// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:21:30 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
JPHG6u/O9B4rgYSC3oilq7F90FSivnp154+oX076nbm2d6VBhM9BOHddaWe4qYc6
9TXlaI+pSrOSv1gqHU7H93vynI11CRDO9617pszxBE7jMO/8gU1v8EOFbvyrSubF
LIWPhjo8WMK1sgKo7ElyYmkLUPyv6H0n8NXS8lXmiPs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3232)
qMgMdyUj8nJA0KGEeCdiPIwyTpCMxLPIpIj+8KcWwy10V8z12s0iF1MVqUaelMlE
dSWaHGdo9Ktmz47tDaow6zXD8D3LGPxoYPMh0mVt0t7MHj4dYULOzUooo5+vqEF1
yTrYAssxwSQd8UUe0oz5g6MoY7bCabpG0jeXWJjmXuvNTc+GP9I8u5P1h//WWFfJ
sr5QOoPAsXTbzMNJoJQPTJi318MXSbaS0KZWYZaG59eYpmd/LEQXuV/VaDdl0ATu
KqTQKGU7W4TZGWbnUdVM+ya5dovQxdOUKfNev6fUNhLmXoMyqK4/MFF/M11OMdVA
CkSwG/23XoHkAFzaKcOBKQ1TGSNg8w5kpSo2qTkvTrzfVgnqXKJW7+eK/l08bRuz
TDt2U9C1E2jlZVyyUnU5MlQU3lkqwwRFsFWIuU40iFnLZfquEZBsyP3r4FTsg9H/
kfgHzE+CF5koCGjHjPoaaQ3oCjjbZmfWHdfW5QBAR4+JNp926TLPfXFdfdlShyCd
GK5bxGtMKs24L0Is0kMsleRZBQ6ZCeNBOq5iVcx05udTkPDdHZc5ketYF4PaXhpZ
7XW+VIH7SzAOLXOZIcS9KgGfhlYAMdKIsEy7Z987smH1YNQ3ROisiFMzktDGpOfg
IKE3P+umxU8WjzEoNBJBvoCtaaufaMkyd+XmdIgTxtWIBptu7xGKu7z1KHwjs3pP
jQp7oKd8AbiwRgQb8jk63ACWVIKXmyUN22C8S+GaME3l2kVIXp/dftjw/41SEG/b
hyOhZELwC6/oB8WOqi650MXEu75OspdvsjOG6G66Ewj/b12QEV+XMhNEn7ejzKQ4
oGdbT9W1LUUxmdDAjf3wBWom34ZAbiGVBOSid/cUW+wLOwJUotp0mX4q7gKERQwh
PKuIQkV9J1iR7gjT76KnLeojI4nltMhMzpPVFsTQ7YNAXmCYGTxBxUjGvIUpvj1D
9vTNMfsc3IuYnD+Tv6If2xnkpWnPJ1v+lo5CtNaNDV6CtBeMX1CNk1Y/tsN9BnxK
Vzy7g4aGd77L0fuoG18c+S/v+Am6DIGWxpC5M1VUuMx5GFqOwb8EvRQNwH99hZNc
8tSudJgST24oPCFjzTgYLYo6B7izz+BO3lplIaRDXwbe4YEQekxVSiZL9BJveEFk
ervXZOp6gTp6C8MEzeMzv4eaHwzsOD8mq8fgG8ErEH3bjLJpcK15LmddyUFz9pPa
Xej0PLCAPpj1rfjRLTUEiLee357wn10RbljgPE09OhEdxjbDQ2PD9YvJ6/K0c4tJ
d93uns7sqWudprDMCxxt26bxOA/Fnnz/00V144rjOXQoWn3Z+lCh88F2PzX4+94k
gBZbGF9lnzgN6zgWJDDmEPbpfI1NgkYinp2VG273WQO2Z/L+dxfNncmKwrXDb06p
FvUaAj6jW5GHY0MLzyafOF3xHigcn5SnY9T+m1QIBki/0MacfYH9dN6sErV/59V8
dp2zIxzyGHe+C/EXcPAoPB1I3H92XE4abhGogUGyUd5TaUxi0gdn6Dj0BCr0LY71
TiBLcArqKDaFiVp8S+d7EwBhUj8FJ2ljwc8SGBDq1U89HtT4304Gcc0PrI50H4sB
sX9x4ZYwEmUXm2/jiswmbHAejFRFT3mBYeltZNEQ7ePXx55CpPytMmUjrlVRpwO8
T/NkU7ar0RYasx/rhs8aNLdujp7aBpT9LmlxA9sqrV9D0J/tirWu/pRo7Y6jCzeJ
8f35IfvDFjpOQAMMrzDw8GN05mSslfl15XwCeqvt2kJyiaf1NHIe0uHvw6hXu7LW
sWQxvZroXeNuSDArMbgwX+/mtm4JdYu6BFcxNtSExsoqy3IgA9v3zOMgEdq20JLj
P+Ex4v16PrHcttWD5+TUsJkNaQZTSwlhfRfS6nPNrLwJe3F9gKS18+QC6KREUzDB
KUyTlVIVhlbUgwQMilFm/RoBsJG+VA+VEPP7PsliQGlyzF0CvzWzdz5Kt0jVLFUl
Cqie6Pg0N43RPlcso06HH3m1AC/euUpf5r85+RC8VxzWkarI6veb35hdHcPpV0Qt
ziEGi2eKd9AW9vcbUJ68EOQLNl0AnWTjzVzPFVZO7zghaTgF+IQp5HdDAmFUjU98
ZqJlj4x0aGnT5CgoF/E0dmmk7pOn+fNZlhcynhXEUGHBM9g2CK7r/U+2ufDkQOkz
elD1/M7anlkh5LVXgZfuEQJWFjc+y3EjTTJ/L61QeuDQ/TQPeyHOYmf/1F1rz92U
Dzzte1U+iXImm26n+6ia9Vn8kJ2VWE9MzA+cU6LAiyVfpyiMZj20rdmj5h76+v5J
COIMoPFAIn6OFz1iujFSKEmkKHd9RkmmXU0RA8p8j+J3J621+Vfob6DfACh25IQo
Vf6LprG3z1++nQ0cpSm026SctaAumlPa1glwTn8a7J4joTrjOsCKS5t/oTjKYLD+
zyP/+diE9+XNwglpIsmH6pniwDek2/ILJ600cOE2QxwXMrmxlDTMq7kXVxmKlAOZ
j5VgIvfFflCctI2wDfg3DONpRGR8CXo2hQq0J1TwI2jb8ea/LrqmAqx+K7l5t07X
yQx4ob0c2N1sKZPPfa4OWv4KjoNEII8h7CrF+0pBlReqhW3lrhAe0BH8ZQJGIX47
iZDRz8Wvc2MCMLHh3zW6vTzV4jy4JrzjBuGuDvy+IOlvtuy7Gn7A7N/p0RmTHUpn
5xjEF6pTZjKqBcFGl2Pv698NjAcDuKtWE/DnDyW6vIZEhNgiMwVdDSsVTZ9u8D7r
JJHZ9HeVtApsoA41+juvtRszM3k2cs3UtukS+YsI1xus0ljbKAVFCRxMOq3vYvMC
zDN5xVGCi4TH4bmsfXFrUQv5OJ6w/dNfoYEBUhpWygf32WKhexz6vKvnjhqbRoFz
TzHYPLiNVnIZZ1ka3QE5pbpHXa9p/FrgqOBzN30baeiSNYGpXBwKpHaWdY5vnNm/
aEmZU2s3pNrCygJaXTd7+ahaCTvlLY3sPHIDa+dQs/bvDPwf3/k7KPDaczuIS8GT
sUhDYVY9gam3EEV1wrx+SZ40c5771/y5huJ1Lqr1QGySwye/EqZTF8IiyolgJrDM
e7Xy4ySjlui9ctvH/+bwSZ2EKez6xqCj+Ux1+ybZMmSbNoHf32ozBz+1+P1tuhfL
zPlj85B+LQh+cvwVbfxX7UjfSwzQREZcgCENgDH9xFlfqsmDmJqR9sciWScEMHGj
Tn3ZePavXxqq5Z/qZ5uKov6rz4R1Lw8HE/oQW8VTCZV9tpjpRsr3tSsqYYeciedi
OGZ/JAIEFGNXDxfgM3J5WRpsWu314RiSpYobg6zlGcUARV/5g8/9Jx+CpOgi4uWX
BNLz99paeCyKuXn6wwvYB/ElRHOAGZccIihiJO7v5q9Gugg5YyAVuAGm082GFVDA
tA45NRjzxqEe4n50hiKe56286wFPGx8q6lZjrhlkYCRT0wVGR50EsEdi+Q5SQN9n
WGXjRQ0c3skJ6wuvPPL0xQraS/ciY+lbtinasVr/izcvp24aoIKHyJgpLua7XtRr
AkDczv4FqfjGSdTYnX+h0WzrRvQYabRviEB3yga8H1a9gxb4S5b0/H584QyjQdzz
dXUtGPAqRnQikPVso175zObWhOQegu1kM49YX7OK7Z0r8bAxwBue6vNpax55i5Ew
hzFDWr5JR4ciWb0UhOmvyyajuYA4LT0WJlQciW9SkUs7gXICUoMLrOhN+Fz82K2N
rsv4e1dzAdxV5Nslgs1395scky9yI291/WxFyLZRl9xLZkMX7jLI8PHMvmvZ6P8t
MXGAseBtQnINg6V2UPKT/JIFdgqYkJKo5nMrzTCeYnN316ymxN2lrCTrI07f5o6A
T5oGjecHqWafrb7wWNgcad9j/tF6iyblCoCCRqZN5zL8FSEYz0AGJE6uZRXvXA5y
1lTOWFMQXRoNzYxo/j3llRurXkP1zBuvCsbs1/RZMS2B8VY71in2hKOq8+nZ/NsB
ayiInaNS8z+plWBaM6uHJp4mLhzz06djqUjPwkiquEQNPRdt2S6blP8Ggrwo9aJK
vyr+wGbuJzESJKf3FXUJQONL3Ue/r5+8FHPsEhqEmkVxtPSfSkGUptToMzGSl5Lm
rZZtWcNwaXo7ghDtVzQMloVhV8nT1K5yIqo3ZV7TxeTb+kApU0UCL9vsSqy2pjDb
7FwUTbsHneAcDlKxKbZ0FRALFEypovY7Ps2l8+zk8k+IOJVqPl69xAFku6At2rN/
yx06mRVNGqQQcHCOjnWlBx90kQMEWewI6cQuovRu1+5G6TiT3t8D/A4xlNVU3c3f
AnHY34/dqKAODii3YjkCyQ==
`pragma protect end_protected
