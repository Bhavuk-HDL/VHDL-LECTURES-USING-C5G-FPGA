// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:38:57 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
exKmWZO/3jCatHMsp55fh/CYSpXk0R2khZwg6MR1BNhKwnnO5IhM/HlwH7J7P2fl
WYqTKfOuDKdzSaXXJupJsHLywKKJdl53zCedVCfzLsghTddP1oUJVuQ1btrtK62V
9fFAjFJAZjVBIpW/KTpD2Q1I/c1kylpzVsa6SjoiHDw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2816)
X6Gkk10iSTytIQhuOEXQoTpQDCwicZrbUmpf9m8qZUby+CgaowJHPJDnWjXwlVA9
EEHnhHLt4PweKHi7uRhVXQPMvQAsaJLoatikFAw7gnoUCDVUFHUWfWeMF/cKD/zR
1erlm8FaY59CU4Dgaxx+/BxyuoyGL1TnpO50pMj6HLzKdxjwv131P43ArBcpAZwd
6EtCBN4KJ9r69uQWdfOLFlImhKQE7FmjEtXNm1AD+iYlMT+LEP8sBFJpwlNAdPzl
sxyjTqNeHBnB+gpNCEqNEFE1A/BTUR3Hj0kquiM8tR4ohnQI760xvHj4IZhOXyzP
SJfDE6zG7OsoYjXDn1Lw80ZAMdmtdcg58lF4lu9ASmnC4nBF39Y6GBr+8twh/2/D
JFHXcY03+oh23C12+GAQokZ2TaLrQZ04ifjKDQtwxkO3jhDrneCuMrlbNp2SAqnI
liaRS2JRu2COAVZiigIi/WZA4FtXUstFWQ2JChUzTKDD49ljAWhfMIuGm6BuKqhq
XWwgiOl7sL5V7NN31OORo/I3WyVCGk77BT1sLJP1cKaBCwdUW4cIUF5zc/G8dEA6
5IFiHE4LInVxLqFnLjaPEiMaWFkyEWxcbPrviYDfuW6MOpO0IfDNYsqg4kZd6+Lq
348U3sEEF4NHXbdhimR72iU/+tI92gYM1QkBeO3NK+wogsvejhakmfeJLUBM//dt
aMjKBcM4eLgR1wvQkYVutY6HeCCemObX+aXlCxJDiiTZa0ghe1PQPVzaxy+WYzf/
2eR3AZUlY51INKb8eZ5KJoGhC7TfYOynumWiueuHqpSdpInG011kN44ND+wIwEJp
pRaWim8P2k5DmrmXkxXqsT1JoGHjpOVPev1Hh4yNhU3cMWbWu1kbsW0t3ND7RbI6
9Whm9RxsTmmYyQ4aanBbsnXKnQpwlQI2d9iuoCnj/F47q/9jrGBY7xiOeKWvlVU5
M+0wqvCyL+VX3QcKxoSkTh+NEYnrqEEU3ehC+MpHAPScveUVmV+YYNXb2mYL4cr5
+j7olUuHOWKEgk91SP9xfsSDnVP/t+dYyJPRVXxH1NtLiugeLbUnqTItWHaXUYUo
cbY2RxYws83Hfi8FfIAthoE/SR42bSvev+283rn7ClqPJURVkNr2GI2iWvTY0VWj
SHT6NvlJdnqLnLory+KnA3w9WYbXJP2jcS2dnd1UNNbyCO/IcaOviwBBj3seamaC
s3Nxi9yzDqzUl3GLwtwZkKI1wxkEDx75QI2uVXkB28iFhAMGeEpV5Tnn4HMdj4Je
IKCGPt4Os1KQg6BVLaAmxuIi/MsucL6DKKIlZXjbzo+z7Z0/PP6/ZBoz17pp+sr2
T/c0y9Wwy+A7xDW1gld1soagsAq7GiZaIWtMx/2jU1+fuBLX4z0emnnTOHK4Hihc
uAMpmmmfxWHrYixCIPzf0DycW+/UhGI8hsi6aq04zWhocTT9F9UXnHMEOPWEBmob
KNVsL9ugDZGZ70mYkyIzVyTaRZSXAWD75jOWlTEH+rinTeGB5Wg0iEkWBodfRCNP
0QRctNQkR/m13aJS9cvZ9s7lkpJ2epKYyuxfz8iVAb4vKNe/YpRWHj7GEdQFt0rv
Jzm3sC1y1BstfOtPyLgY3dM1n+IEjY7cjsEFHZ4Onbm6+kGaizZgA3SbIZb6naPt
6L1jxy3ib5aATNnO6smqmHX0HSqw2b1xvW/P7P0gR7RHtheckE9Y5ahs3TUSs2NY
FYc3dKuM1z8O5neaTYoNj+z3NLzWse0sd+KM9n82yP1Sf8f+6KJenOQZj2pABRN5
7QpL8ciT9JQlofIwJJhqegB1NURL92xr2pMpdlJ61SUmONDmTiNXA2HuVsQiIcfT
5cprKhZ32boyrS4A0pDxBrNlNxutRYGMgaQidZeHeTcStj/O+DorAb7xSm1w8YpT
EkuwYPceCaZCDVIDGTEh+mJ5jgOb9bYYj+yJlKE6jXsimiHLEdJwpmC44n51mfE4
na0e0qw53SC13IROVivd8pTeZVm2djF3m1GSp62mNxomP9yCSTMCJXMVAoRbzMif
DgzOVlxLYoypEjqbeQ+1W5hC3dDt9bewca3ucbKP/HEKu89VtpmoEaOTl0uHrvud
2hog4uEJYpdJ3ijYzsB6dPAKYkre9bMaU0H9sTcxNAOAufsOWBt7tlB2yUIVVdmM
xkdIUUgmbnR3ytBYzpMaAH/6IPc5XWo3/XzHislPJvoX64Tq5+t5J9xzEJclmE8U
m35xexT/877deN1ZyD4ILHhyjvjBgVOlQkPrhD/vmJH7sPFIYBl8Ndn/zMaPJ35V
syMILUhhfVdtB4MWC7v5kPNwChZpgDLyV347TsU/4vt3lCQWJVn2VGs35oumhE0U
9wYv5FIGHpX7js1Q/WYdXDREnTJ9+F+0Tjdqkz+sb2O9TLcBKRSa6yY4IYy5ysva
MZP9BKB+yxe4SuNQ7liA9yTn/QbFyw/xKlJl7UpzM1FmsPFpdK4sN3w/LE47dqow
7lxGMOShRixjyuFV00H/IA1xADLESs/8l1M0metLvheRYYyHb7B1BiYvWQZixYq5
iQV6u9ASBa0fceQ1TD2eOAD1rEdGUJhm3oA1dWuSzSrTcc8peWpJT0tVp+GR3mym
T+NraFgfvMEyrxP4wk3BWUNs7mrxSb7CUULzGPKlj9DlUvS4cz/MOSb31EP7Hl71
MMGkC0ZKz34rQ51yIK61zu9xEJpvTT4pVPWlVk1UovbHk8jVh8RGDZ3IXaZhaiCu
gtH965oRbSHE2XgHXiULSwXDtBShzM0pXFGVJ5z9XQdu5ppFIMokT4bwe8CdTriO
CP5+Fsk+CCIYwmJrzECJHpk/uqo1oejVyg/El7bxJ4aOXORocCbx3wI424ZdT3Oy
zeTQLp83inac44CNLD506UA12UXe4OeQYRutctPZ05jnqy6gwuB3ptIK1aqmWdGg
SL8tu1eNcjpPewLTf/u3LozkGvgly7SeEsc7T3R7yQcVPmlZjNFbWDDOfy7yvYFX
iMlAO7fMgQKMaMGmE9dzEinfQhCINRkVBmmh4uWzWd2aUOjx/md8ttohey2TPE9b
YsXWfV5gs9qu7SqInRTjIvajCc+2ncR4KLimnrrGY0BpB5m59YTTmEoJ+1si0tL3
Ii2nseTeT1YebJizKpve9W7fcwK/Pd7xrAWMKGBYy9psHGHLNNXYIqAcWmrNATjL
BpLF456WWHf3ap1ReB2F6tEkEoWj49dWPmPaKqgPXrwgAkjOmfitK/p1ALgI4UcR
ZVZRQlbSF5FpYj7Zp2IFSOrOPxEW6+tLk+T9gKPG2Kjp/XPFAL2sJ1W1FW5/aTT/
6koIq/7WyCzfcW6IhSUXoAfv6YAo0DcMTYEZpY9U+4xyYxe1BYiKuwpocFJ/Q5au
eP4M31fYbQRZT7m3UbS8cojg9gDvA7XppSZmZ13EIOPfMzyCbmOY/rmTPAFUWblY
9+6mz+eeTVLl7jFh2bpSZfhW6HSPk3fr1in5/Kf2hBfZRt9eJJV6GPftMMhplKaz
SnRi7cBGC5bEEKxWKqstepE5sRMHrEWeDXERFvVKGXZoJHNEsQtkSnlRTbc74jqG
xqXZzpB0jdSdJ67149ePnbKTvqjHsKWMtOYLEl6RjPNhRbUmi2nFSb9hb5RgZPF3
uV/ZRKLgugCWsijl8tTeb2ja9tN0mad6z8Lo9hiL6ogRD8UsKcKD4dTH4+5wsoSW
oGNiuM3s2LWP8ecQA6PnAJ6lqxWJHwHymrTsIRom7Qc=
`pragma protect end_protected
