// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:17:49 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ssyb8IyN+mNqm2hjj2ZFK2gUWeoTMb1bDH97nI+C9hQV7AR8W8PJ0oMKPNF1pE3F
CGpbOVeSfO9JFsfW2AQBBqW35+NPLZR30kDrkHqYwC/6328Xa5CPI/WdKTWeocxy
73yPa8knUpVkkWE59nfshxi2oOqAOBXiqvp5hSjPTWk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62432)
cjXd1mCocmXYO5/C7zwbc9ycO0cuOPrynjonT4/hWy1bYfHGiOXcRiIzwp6r4SW6
EE5vkmk5EdSjco1TpyHP2/6GJNssN9lDPLTOu8ghJAB8pIENIV90CHrow+4GCroD
IEyAqirR8tJakt9mfMlg2HEuu8UPzzcFuBjs9f3I2RPB536iRQqtK/QsB6CmN3eF
OfSTpe5CxDUJfR/H4+4OADj15eX4dZsrdV35Knyjbh4qD19YsmhoZGyxc+d9ft7r
RqitE15TpM4fH8/22ftuaeaLk4WNS5tLBnXmzDGYOWsRMhMWD2ufR6zjl8VhEUTX
suIsLkyXZHWZN4dJBT19JNDOqt6XMtMmGVjBPnK6g3G2zJP2vM4CruKiBIPQZwU0
nHI7JAF2w5w2EABpyCq7A91pC6Bxd+jUHuh6CwhFj9fh+VP1iCRIerHBJrpm0xpQ
dwUYthwWBcPoJcIl1CwfWRKcryzeXN6TdetgO3Az9edmfRRBveslTxEn7Vtpv2IN
KnrHBjxghXao5CqAw5M+GNibWFKl6mewNDt7/Hl9TWJksN5lAnHBXYINtj/y8MNY
gkLeDfsHXSqOejZiRcWys0IoHj9likG0Gt6Bngy+wGzoNWS0E38DP+blFuszzT20
ZS/H9QWS1kou4d+1WAto0Fi1fGbOHiHZALOXgtRtYVbnoOa+bxbDTsaBcZE9P0ZZ
xe+VV6Fej3ltSnV7Gv2xdZwu5Vr5G6VIo3rFBw8B0dd30eDy3G1O45MvZI8NkfFZ
Dqy5UU6uhxTCJNzKmxx+NTp4t3jbELjnCx8LD+6a2rStNfrv54Yf+ICpBE2AC8rW
zXX0q5v0jCyF9rG3Xfjfq5MAM0srZLUU2/XF/fI34IozdgDp7AkroXXLCRgg8Lvn
hTImBu3tQKw2TrmhreuGOuKlRZj794MTfrgTOpUn+OrDAyCn8U2J2qSk8mKEe3QV
IRtPd3zCzoZYXDJQtgQAakd6m10OoYZOHPWMMSKdPy5a+Ys7hCkeX+qqoOJ/8OaO
AsXQA+KszmvOIPGV/Bo13wyqtE7s1+xNIIoaYstovAzTazenq5Q7I4ipjX708ieV
L+7Sr8XjqE9/vssXn91FcuW4zidA/6CZ8LQJjwbNfV9bUj0G1zttsFq4RoFwtajJ
2CJyUGHjqKuigq2iMt8gY+IHsNhI35hOsWt4AfN2i260DXwzWbpWssyVrAsDF30V
i0UONSoIFcVFQcp/K+aJRcA65vt5cc97TgqYFVRQwRUIJhCJt5xULnxrMBw99qVD
+s6HdHv+SNMfuj1IDa8jXH/UMIwarlScSS+G58+4Oo9sPcMopLLem0BJKzaW41PD
XvHpRgJENpYZ2z46fbxT6FrJORckB+2ghM9OjHLP+3ZvtTWjte7jD9XPzIGNbYnm
MSeIB7aOM6PCxV3QVDz4aFpPZRive4qHmsvPRCG7A+gxvtzrDR6Bt3XPxP2uirZO
t4+CN2t+3OlrdwBiSOebbPuJ8YL3KAKAL24UuuwQPPO7lz4KXeEwonJSsGk9G76u
iE769OInYiquWdov9SJmp6t98CHmSI85xwmSu5EKq6L7NzGysqu8gs30FAnsvyqb
JCT0RT/ArAig8la5QcoIWHKolZMlQDPm5Loy9ITtmFm93tGK+eruEX/iyJjv8BMQ
Vv1qowmO5XdwsC720C+GP3s7juwPpdqXJV9/HoFfaX11tTHjIEYMS9M8Vvi/LZUw
F9zfO54aGQ37PjgR3SCYEFOFWugwu6DJ9bQwsgfIBOWNAaQsgcwU6b6S+WvDED5h
iDnyq9sqIrD63GorXa04HJDsCoDX3KNGwdZirBrXPBCh8HbyOC9gzcFmtjvaSNF8
ONwKNWzxYkJyyGD1m0s6ztNukT+lpD7sACLpHnKUrEDmpXinNm1kEVM3qO6be2Bp
fy3yLuvkNJPWQwDTZVY60iv/t9OhUea8B3X04dk7zOQHk+XaTztv48VUpZKvqj7Q
6lXikRm1N5ECxqyjmF3VpMoEZ9ZAURsdawx5jnTXFNXytIypPfiraZROrC1GqEWp
mENvLC0EMv7ZMduVCHZGckFeqoeF6Zq2K6/+VuZTU6ZoOAJRfwzIz5kRSAg0X85Z
I0s+BFgJ7uQiTofZ3oKTOKAF8JQHAnHhFNSLOjb3jMSxFnTLdFDKHAIyh+ABP7iv
zC/hUFrxIzMlF3jDOYWWwFUFSaJtdTd0WoLx0Nutpd87v2r9VSkbsuFR00vpBCwG
O0ftmgU4o7QvEFUzqU1NpS0oZH4WHzGG5+2TFBQ9Ul4hSXGDkecL5p2lEgFRvu0d
JWKjAsHTw8S5cebokyjpJP0dRZZYCN7mfHCuKDXmHcIUfmmv1ItdIaWXPfMGzdK4
IcDu2/VWfvjpuSNJrjWiLIMI4yCOQoDrrjS1GuKiz4uE7Wb32L4oxZWMdwjPHF9o
K9ctjmtejW9N1DERGnKnb8rN7MOsMCa+dGN/8OMvKBUxXG3fMI3MDtbVOLTbp3c4
kR7mZ/WwRMku0B00cMH7Z1HReSRAxigKl+QWOsImniKFWyBYrFrlIGfODlwCdYJ0
Kl7kauV2yl4mzxRBZFJiYLxLshSODv1JkA3Qi7CptAl1B0Fdyri51z/NZm/5iOHH
Mz3JxTPYqb9VYGHJ/7ft5Y7IwNuQRN7e8oUfkqHO2HZQnJO9b4QfvqXJpcZHzVQl
jyozw/a9hZfge1VoSJ79MlWXIZRNvwl0S3vrnJMVwnDdhQfnjj6Ma03C1uB+Lnme
Ljm6Js3tegSgj51MDkAxKifvWYSmnpVUEpMJpuDAnTsakXzpomKofVQCnY+hv5Kz
8bAuJ16G1Z/Z7/gEIX47vd3ocCyWkZeA15D67EN0lCzUhTUcVNC3/gHjQ18Jchbo
zCK+kpXja9di2hAcATrd2dHZsLVLum2BBmOYtS6s5mF3aosDlXpggVEGs2sqOhvQ
meCe9fid73kCQOKw5hccDU+w/kiXF2UCHluDMSNd1Kg+Cnpy1QCG6xsjWI5V0MTl
EHM7gBriKv+iNqPj6yapa9F01EhM/UYGHXq0OWH4QIuVefVxz7udt28Pc68wkULz
j26nsiCaXjUFnj9gpefBoY8RJmDNmnz/vkbZbr5k9YNs+YTaxD/z13AIPpg/B42P
9Y/UcVG12VBC0QHMXFRNHdY6L2AKrijNt7oGpJ3LzHG/+GVftk3or+Aj2vaLfwEV
xkgqoavMCbMKLtnRF2lB3myarUZ3ajhmCmkPPlJpuVIGcNfGGTGR/KRLcEguKksy
SpYsEoT1NYobj2fhsvTx6k78dk+iPmEE8H0JE9MAeRlsMGmFeNAvkGQuYo4SKf5G
h6vwsG1ktYedgBtSGLZ0bLuPjqd/h0o0goxhmnLL7303qnogXBnjTYWPWJppjuFF
LHiJvUzg93Q4/20oYCb8606AX2zbeFdeiDOdbEqTCQGBQNH0zItxG2iuDKdutVCN
4PfNe3M3nfnZsSW69I+0H9twWxlEx3tWANa/B5cwe3dIDdtl6CD5z7YuTJ4NKyv4
FhQt4/DNPfG1BAW+NO6PjrArtdASthuhaoUK+ZyW4USsEng25nYw/sAhT/IwTZ7R
aQNrO1NblxZaaKCIACn4yJIrTgClSrRSJ0WsOBlLxS0raq0BvK8WNwKJfGjAH9eY
6wM8QypL59FnV95bbv061qgOrZmyvdhYJjV6ti4bhqmU6NSlbsAQJJCPntFEXV9Y
fjzg/1VpCERj7z9rpdxX2huPU59qMXr04KImCxPwqUZl48ftWPbkXMTX6dXJkL47
nQh+IJmFxJX2ubnbnwczBK2uxj6a5KWHSmtqMWYsBr+TDUitdTNPQRGx/WMXp0Dj
A11iIS4/WOvMbUUEeawSmRq5zKmCGzUp4Zt7Lfb0pZTOrAVC5TYR6pnNSIbwBnH/
yl3+ujr5iUFhjLOIAnC/+LJL/aBJy53D+w0bKFfjpAmZJ2oXoNJ4eAA5xYeNfMqk
BFP3QmQV4Khupe1MtNLjsOo3eOHLW+0zOEVv6VGrJLyyMxA2UztMgUUEqeQKYOC5
g0qw1BV7nGsWdZYSg3meAOIYlq7Y92VEzuTu2nySnsds7ln5P6FkFHOsr2XOVQsN
F7ycGSJ8bZ09ELDgxD4I/EXWUmNwwxccT7IXZeALjIg1L9r4ovo7TS8HOpPJZhCq
tJLUPZZ4rQq6XhAPViCSLQTatHbzkJvAamzy14Eg3ZkJIQtxGPwQ0aTKDGDYAJ+V
xR0P1FgdiJUCFvWm4nPUXLy+TFe4JVeei8jFWvkpWT1eU6DaaT2rCy97fBhpkYtZ
1h529V4Z+glv06qA2ZAdnhA6SXDWwpIdgIo2sW4tVqMDGORJDb1jSTlr3Gi2gDub
a5qu0l5aBS35UokoOLvOnDIiPyFQQ2+TeHlRXjIIHmw2K++gOQB6/EOy3uQMbigd
tsUFjB47YuaoGsd+31Si93ftVW8QwEIee4xMMVyrqlnc1vZ9F4vNZAS9Jl+VRX+V
VrAcx9VdXexkE1KI9R/PQANFTexNk1kQsxtwVvHPpM/q1ZyyhuZZ4E+gMv1MHqZP
+JaZEXs/RQABYgDRWUiOqAgpIh6yqquRhu5i9vTW1bTy2vW/gDHwikdU1IolDh/7
vbNt3M3Ow8CKeglgey2JNiUGwhfU4nCvPVjsKEjwg1qnNcD88Hfug10RLSzPERuL
CYbwsktLIaUroXfDl69OHZl8BGwfWm6rVJoq671nw0q/qMk1CAfsXi7OdS9KtxAm
CFfyvyy5HqZUhuY6+hUa4TucQKgJHMYbzibCn8JUkHINFK+Yjt5pXS/mGHMU7hJ2
O7LsygJkbBKfXEj/fkVNBQG9P5sYpKXIYmXaOUlEEV2DHY4nIaE3DCLAHGZY5PUD
nB9SL/jYf69Sng/iA+IvaHaioYZSDyLd2f+n/PXGiAYPvEwpKVcaRjQ+M+MKEbws
Qke3XzlKflLEBEP+lJi69ZlqhTHK3KtKJB8K/QkWDA4M/ZcLsvuCnWiytzlPhyJ/
Te/r7RhFM8/g55DEyqH+ds3T0m8/Osv32edQ4rTSuS+LwFh2Cl6JEfl2ZNktQ1Fg
ttVp9lpMDhR9QeSURtO0nca+jiBzULVn9qhDm72lFslTV0RpnIVOZIs98pR0dNxl
fIDVmQPzhV8QwOYbExAzR1dTorUzsl9EppDOZ1Z++RMCUhoTMRzP9h6rn5HyaAG2
VauYiK2/SFtLX4aiNsxKNaCHCnufXETriZNS0SjJAyCrx1yqBdy9YYyTl9M4RAcp
CScGRqdZFK1I3X+ZBXCgXKKRqaOU4a5nYQ5eSDd/F+6vYnNi99dSarShnnfmu9a7
Qcdsceeli42tZTbOrD4c94hno3m50VvB1NR9iJEyaJwKIR/euOAzLujqmxLfeftI
VGVhzFKbLH7V8pZGO8E6ZM8xPliBM3uUDTG11K3sQs2p1wxcsoIJbviWc3339KfL
groP8FiLV8n932/TCGR5yElQ/ONCTHyY7aCyBZcQLNuZFW0jw0jG5J87kXnZSTe9
tqYhPXeM54MXg8dU4wPCaLELFUD8M9iWpxa9u71l5ww/2bO3K7Tr1ZYF9mt8TUid
2eBxI46SZeBd+bXmSXTp9pj26PQQWAQcxdeyiC3yYCvZJLvWmedgGdiC084HRbU5
8jCh6iG0OGIluKwr2bvQ6lSApV1FV4VaeDAeTIP5P7IxXon7XQ87lIKJl4vv/2an
3tWMrufL0XgwJPtT/cGCbNDID0uiYGEXfHAKs1nGc0v5ACEDr00xmF0j3Pr524LB
bfQrXAvsPNCayy/tehe6sJDZyXOmjAFtTmOGF70RfkM498jYzXNCDu+hKdZ4AP+c
U/2m9L+M9dxvDjweXTQyJ41upsKs4C6lH/uYUaNEMvMFNJ9aDcpq8ZZZfyYV1U/s
PhtbbIw7qOz4RLLSkjppQCjQ65K9Blrl6G0aQdcdOBJIzTvA8EEaOPZT5hXQ+9Ht
Yig4ihXjQtGREOntJOww8uhGmFrXsZp+5Hg/4N3kxNT+RvEBMe7MxGgF7wINkAvc
OHvh/+K4cegieXaGvLR3GLwjRPKSP1N9KNBPk/lVyAQXVP1F7lUOOcBdPKgK+eva
7nKEad5/CsjMBAtsCrnKC/eRRp3mDhs+Z3InScmuaTAGfH/3xOb9S1GU6aecU8XU
dx0V6NI7GOa4v1j01o28zPqLY2m1a9ZOu+ZHAM3XrsgA8W6UY9hygoH12NDLWLVf
fNZfills+t1PJF66aKWBJXMf/vMwcnzuyXH0rdRphgz4H4iXDZ4DDmSo/wQIw4/w
aZLi3jjw5bxn56cNOZwGWkIfcWTMkLgyzUVsP/PknDoxXrwhPDPgq3V8vfJ/B8m3
Wfn1E5ig97tvDIseniVdkrKneOQwmwdr3QAAbB9+H23m5OG1gz7vA/Yv4Xs0oNKI
ke4B4b1jAwobD6KDKrNAQDJMAGbC3SQvRBpTlCZwMkYqRyf/EWBj8lJibi98e7FD
4UG5/JddRXr/GEulowQxEh5EEn5H7x/pkVZSjw7f9kHXTJd7Q4gQthnYF6BY5vm8
5pX3n5uoRoQ++IQbyZE8AKvoqwVRGzP7Tkp9B3MyEEPSjGUdWbLHF/XT5twGUsma
VAjGC8JDh2TaMY9K3GLy7WcJKZQdA0JgwxDRfB1v0noLPWwPApIjyW6rdqajJBy/
JWCXZlJrNcfE9QZJsvpvT1/HvQa4fkSvoo62e7SYTRahzCIo6o8jWDe8ZnwxoMqb
yNvaEBZV3h1dfW6WWsFoS/4RMIR7Odnz/qlvJx7rC2+Hp7djPDbGbksV726JsZGO
PZKHE0/xEc2i3zVAd3/3xtjeXpgmdkCOvd1aTULLI7cBrheF1f+UtdxgAJvWJN8K
8BBZtrgoiQDCdZ32giUJo1klHavMOpD53CdfTLQ2sLx0SQDOeP2CE5lzhbRFRMsj
+Lv2QgZ0l/cd40j4oPnPyi6EwuO/n3T/oYScH6/sVmqS7HiVaY2iaBnx2AOb73KA
Ge82PHnoWW5cfQFOLjnizxbxx367gHRyQ6UUFxoWC81GChbD+6AFzQTG43REq+F6
+LnMqt3ROgokKjPke7GgJ4sfMgi5QI6nGReX879qyQJCM7/3G7A8Ix2fFR7UYzje
TrzeR4d8CJ0ejYORIof22p5QLIUS5X0P7R2qjPhvZc2w3c1/7FcHoC1E0ZXEAkMS
G3VAnSxDvX8D70NTlQZll4rbTmfGaVSt67TwoXgHVBwRMFcEEwb0OvOFdbO8s6yA
BBu9nFyq+2CmJ2+o3e6372D1bsktmRKU95m0XXcTaGqDxEm08fdxxflV6uO/sS5I
5fEkyErQOygsKz3RIT3sretfjafw2p/xblVUBsuicrdpbrQgZKC3LXs/Fl7Yc1wy
Ueq7lcOGJv6aGltffRQA4ed9HVWDHZUlYi4AUldfWnDbX/qdZl52KowHcpszLerQ
DGvFBVBCMAVgstRSXTIvkRgwgYIk62+98wzwTbBgN9QfShzRw0q5RbEa5H6d3U0k
b5B/xNcVwo8vtFEv/aHVyLfJeYBQifOWOPJC3l7/Sy7CKbN69bASCVpTJzzGwzRa
wMwmtq0RwWw6yV2PAFn/yaztzih26Si5IXlt4rM9zHLMcxDCZ3bElc19Rc9R23wD
zY667TplJuhZ+SpyLu+jyXRv0alENNgrOSzU5z0QmCgY9FuoMLwAGTOhMG6nXTLt
oQ5Eb1BoSK3NRAk6mUtDrOoQTmawJKMb0njvER3mRVeReEHXgOhu//3u7ImhW7sI
3NF0Lc9KRGDcjvNaJLkucVt2jne9W4DW2RTsTjAF1Rx42qPJrWyg1ImTXN6lsa6y
8CPS65X0JkWGchx61xNIW3SQ8M70dZWF046Tnak9cgYtT/Xq97bXRFjOMFs+nQhs
wAc6sm2rzieBev9riNYweF5GtB3Q2thsCUcmiLXOMdGuJd/2iyxirUrXy04Uqr+L
D4QWjePPHEhITyVzE1ws8H/HQo7Ut707PbjbiMe5mN5w8XrgAUq0BOQoAxrb0ra5
F6JzPbbNbx1Wk0yz2mSklKY26rL6PeVbqW+p29G04xg3KaVWmTH9tAJvNynMzfGg
yKCAHxDh6vEshRx88hVvMm92BXK1WD7WSP+MtPUtnE7xNs1jUT7LbTMVcQDe/9nm
eYR6rBnvRFw7xdX5vWeefNUQ2G3sam/OqdqWLJLmxw21lNh7lIPzI0zrlP+ROOkd
3eLHZKbD8AjLwvCU+XxoOhnEahn8Byf/m4BL8+/u2/y2enTX2xxVqI2R01NbbLSb
uUxVEKXEpGkAfOwwnU8buG34Mru/Ope/CrzfDcR8dDFXY+VQMLWS5gAD+zimMJYW
3F5I95TIsUzSfZD/nQTfBU5iKscZk9oH1qvtfJ4jm/2v7+oTp61f42g18CAa6U5b
3m9j23Eb/e0h6W12gyN5w+c0o5eQd/RyKKHi4b9hdNT0m3wxmnm/URPLrOgAEEXJ
7Cb5+4shE3EMfTHrPrqcx8o6SWOi9VeWiuHDl32UR/hh/ekN60HF/4BGJsFuClYO
xy1L+BzS9hilgL5Ak5sZZZ7mdOXcdGwzlfMrQStYJkfbgvDB4D1IKz5AsCMQy5rR
2GWD17JXLYQjXukbM3QchXqgITek+WvzXua3Jdo+ru+Kkch3ZBb9om7Yyjeg+zdM
DlaM2J+hF5y/pa29rpJjGQXZZpJaVwI9mgCEr5kJk8vaydZC52Fehtv6OwrGxyx4
Al4ccdEc9WOxEjlnoSLFTnVcte5OjMYIRoKqjaCq1fgMZzJcWCEERZdxPsRYcW9+
gWZgcclvvugHvb/9yPslm6/hJtvo+dfbqkGFYjTKc71bzLB2O5bQZvIkMjDCrtdR
LHYv6T0PkRoKsQCBSmwc8CBA62+in8uvq1j/CSQl9+pdnKh/TIicbMsc3HXolCTK
fQ0wdTwdTZQPeLxXnFo2brNZLL/HionVCscxwWQIPcIGHsR+7lfnYTUmpL3T938K
E459sbzulveM2n03lvW4IunFSfNaeYIKZNn9Ysv3qEmgWvnmOcqZ2CEikFPeWPyN
i75W5ej4OrXSGAS043pOFVCLpkt+5CAIxk2REgxBCJQujgKzW2/lRbmp73cF0CeK
S8prDRrzNSAc1zggXHio3QOHZkc/ArQsyqumXT1bmyVDA0LfDgea1M6+/U3CDRNb
N7El0FwpBBhDCAgaqH8xDc6BxGR85+ruoswwoBn5N1dNSNxcDn/jKVZW3SAEHTS3
YWIxdgHHAmzwK/4OcoSJk5aBv0gOQvz47dlPjM60Y5XJKmP09HxQp35W8J8pki47
Ds1nQR2yCBUE9cssVbOeqdsEHsZN8Y3sL0703hQu7u8DpzAu/aIjaiVU9vN4ov5j
HLwjpGKkLTw4G8NZ/tc5KFquaNeKAj5FOPgbBVW5ZUfMxKeG+EnhX27tfCZouWYb
eZogisYd2JIYKiRIQt7jx77B5pGEUEwG9YWN/GTUCOOeiI/8DUkaI4wKxD8ASUUE
837UJw3775SUstE1L8NxDk+rEemeZNOAYc1gGSQeypb57hECZFH6xC/9VRlhshZp
gO/VvUEmTfwR4443qF/QsWoH1Wo0iQ+3X95Vz639xlCwI0HNKDMySfV6FtXWyRCf
ebyxIcrF3u85WEiWrJGfcHw1qH6ljTajIvJ+7csTpI38kPMU0WQHQgr5q7uKY4i2
2t4oHuYrDlAk7r3GOCd8b1R3KaPhQYRE7z5yPJ7U2AdCFohFQjFe/JTpLjJFaFi/
NB6CgYoAiKGCip+eGdaVFu4XTA+KBtTuRSuD/cUmYeMKFOCPryo/QWhiJyOjdlKi
CWCWLcFu8/9j8BvVm9dm4WSrgJrYBZ3tTmFI0xOV6spIlUXKl9KNLt1nm4ZQnbvX
bPmEhT7pnJAEuVEzOt4emU7Jss9reTg2wfBvDlAILAJ54bq0+imPRPIXs91XKVaG
g5g3iAqZH46QPHa6aRMXtbtI8w3xdmpG6PIhBY0/SujmcxPxfjT6OKpa99chRM41
FQfolzT1FSWoHHZ4j4GlZWj3Ex1T1qD82YamIce7aa6yLFjrqeIrXDTeXXyiPl58
OFCKOG+E2SD1MQ92OwsSJtdHr48yZfxgDpKFPOcajEVBOmX1jJkoCcu12yzXLuCd
rjDeqR3KaB+KEEoPR/fm4ZSxnU4n5rtpJ8Bmoxih8DXS1E4QAFcFNBudC61IwPXz
bgXZ7w1tMe+HC+xAQ0Xyd9Gi5xlqkwtcow7/mteYNH2RtrbfcQOU4JWqzX3CIYBa
ETh2jbAcamazVWzfRjWrRjPXV64PL/1N6SVDCOGzPBrPFFxcrDIS6v7cZH7Z86Ju
RVAH7JcXcLY4DFXLRtUHIcS+Ggh0VZQTc0nTjIcpd2Xg2pV3qr3qlibV76mJekhm
IjIXfA88offkvp5J6PXiRGh6OK6/3ZHhxY7BV36MS1qkI2mmRM7UJLqnDO3uBGwH
ync9XtjTJ4D5XUSLNtlBQCSjR05vEYbCwzfNfCI/CGys9TKmEeDNG0v3vGZhaWtL
qyFlczKhhfiPezVPYAI7bJoywnbjI1bSiOgpUhzctgSuqO558UvLxEPsJBIFpAIJ
K6pw6NZsPW3bvagu5z2Cp9dOqcPlXc/cNogXEVe2QjmfS5UMC6kf0KZUPO25Ejqw
WxzU81/66JUeIci6qU8ktUTpYlu36oL7LjU3/IfVFhlCtjAUizf5WF26Jl9xZ8n5
Jmfun2uzK1lbf/IpAhjmw+mVf4WYCRe8PAjgEYrwmTvS9WsKvPJDi4MdSfixVMRz
4z0vTbqh5Wir3YtP9dNe+iof+XcKf/SYBNvwaIc2aa+qAbLVnfOKFIaVSiaklS0+
c2sdoxUXvlVBveWamMFIcuVRYbju99rygWEGEbl481YJRV31l7+dVXspz7wMry2T
BDPLWh1aT5WRu2ZVZlydh3i69FgiUTLxfzdf3vf/Y4oDm8peACjhcqqWmcHwygO9
aVuBymWec6nCOUtsSh67tUkCi3WHbduT/UjcgLgZKgA3rgD3ApwR/fWjf1WEaGrN
GJO5quj4pGK1JQfvkReiT80mdLDsUFAJFwvQTCo/79lpBboIatLdS9DWDM4jeagl
DaokA63qAg67hLt3CFsQG8ExTg/pVuQ3idf6ReOWn1rLq01Hj0cMDRGPvPPfzBIp
joE23wQhaCl66aJz8nxkSaq5Bxk9QkxafdxCAZ2Wb9FObdLzyM7UackRAEanZEdS
6qlFBgyvlpbj0mnc4m5hoIE9lwlZUgf1tcA4Yr95gRedGRsPeb3ZnFJNl3OFfYXx
1/0UkvfGgnMSaaj2QkIJsi3lIkdj4ff2d/7/Avtb+wo2lShNQ8CMgm3VELziqDfq
6EOuy2PxzTmmTVNduWYNZ5GuW56afrdxvBY9MauTl2GGmDcMDGHKqyBs67lFM8yo
QG5aA994aEvZ0AOvt14/7mQ5Jz8V2eyjtHR+GKkhnzuRC6Hyk9/74O6au2L3pkwc
QGnFOF9hp3EX3OZplnPPA3u2Odqxq5glHpi37Gdq4wHrfMpKfHN7m4hR3aGoRDx/
lZLpqNSYxVYVzj3abm9ZsUr2RvH+eOnc1G01nZNrXM16SNrx2eixfOoniMyUcQyE
qe3qSoUOUN6jd+TkrGLYpYHj47DUiX8hOumTPMvaYkr77w/EbQ61nsc2XC6+N90V
8dCFttaY/ZQH5X0dJsAyuL28mR0ZPWqQSTmVnYMr91JdyFgmUOri9ZqMvBF3rTdz
1bFG1gFCjvuV0dhESlDd4vLYVlUGFEXxvDoaCwQ1fbRu15BsqkUetzR83xphw4yW
s21K8BSLz3xCyipikD4dO2Cv9khTfcdE65t0gsPPdVoL82/4/klakHXRNGICbeVa
vcpva+8VcSdydiVkQoUyhuTrSr/+MOOM5tkQlKMu4E5TDnKSDwe6ia0U6RwanT8Y
5OX3pkFIHVkQ5M30DQRbwo4zm0kNXCVh90+25hDjBZyQPq6zFVRMlThlQkfDYsx1
JxzYNVMz7XpNqgmszcWV0/3N1U/NOV8LlgHkoo+/BDZlXhA1kaqDhTEptsxI03zA
n4M+TxnITZbrI6VcZQ7SkM6Svsz7izr82ihWjqeLpRQWbELP9Ul8Mupcye6/4dQA
HhUbp89A1QtEXrZ79k+PTIQP869IMiNaVTuJzCn3stqsLC9+vRdfVTSIkt/tHtny
OCx7SO/TixviC6hd1NJg2ITj3qdFMub/Hhx5Tg83NkPN9iE5fqIxJNjnFRMWx8gZ
ugwV6DBpR9zuv40EgsKBxWTnORSZvtISRnwIs+RnV7RMGPq3fclQy78zpJeZBd3n
sf3EvOWAtJoM6M9N1BDAOMnyilSXZ/j+M/uKQWQ5U6AaD9xHB37bddlZGSD2YI3a
7hUj0nGeXpzNH9e0aSWXl+43KjKE2wQEIPj/1ESxlNH6WLvxlhBAm1MjfQEWVjSo
YnlVVhn0L5V3BJi37o+k6lhGMwfRMf9NAf027LyypmwrAeNoiMtc9EzCIZokptJN
3rhe3o1WQw+J19LpdV65lLGyh6mJyWfBOoLqV1rFiwszlzy+0Kj7q/L+QPpvubkv
7iIXsTqyG2VTzH2PDoGe8iAIOiTYt3w5lwm0ZH1OUwvKtANSqiaebLBoo5ZDtPLw
NNy7p3dtMRXHbhSgi6W6WbT1APYaGLWRPOUdYx/DdRUDRDRqW4jvy+ztnhCvy8+Q
cbAlI2pPXltIV9vnYJHKDfNuUGO0gzzzEQ3ThYVhCpZiCYthhOQjz84vAbAS+hvy
kA7vPcmiebesxXaw34mtlJ3XEfO7oz515GFnvw12+lYIBoj31RgRsh+h8ZH1ZDhf
7VSZBlsxt+y5DT/LrNXT1mkRmDTimgWk0xIfai8Pqmrvo8O/rwWnn7Odx4bbJE4t
Ne5c59vOhNbZ3ly/9sXUmJNy1c+c/1gSq5HGFcbmia1xSFLhqaNckscqUCnF0fK4
qjI64HrtZ3TzlxjSwdh7HVMJ83wlUPtL3tXHRLzMMSlzSNVtAkOlz7y8hmmtHh8X
cSwzxXxDSej+6u2E8AEVWjctjIvlU5xizlo3De7GEdUd48gbfPX4ceokFLmfs5ng
rOESxOePAvwZkQZ978t/YzGmHAZWkGEr8kwGbbemzrQuxi7AMZD83t0bHg8aI3BD
N5pwrDaB1crdRPmf4AZ3Q3k7UELBA9QxBC5JZwvGi53fZpy2pOdlzt5FTFjSa0VD
dom9zK2yWmBnHkl5Ja2Yd+4/yccbx6zn/Or8rlDbi3qmBWiIXVnwLeI2CWwiXQyf
wquGSKyG8lHUXDX2HKFJjtkwtPVSkRZNziMG7A2QIx1No27AL3m3yyYZ5XPXko/7
Q1B5gpJcFSVocVcY+nHz/oNupTVWuzm1WR24J8bFcasqtEsg517Svr0ODA+wxqba
DVhDLVBnXsAaMG9tD17vEKKS62JJKVtz/gJoH9Cfxyc9FBhFc6ZdAnEYJBk/tKYG
PP8O0lfOgZYfsgRCZfzHZ6+YtqPNXZt+vemij+9FIN3JiwzcsKJLxlrwYTE883aZ
ycHWVMpBvzNq+t8e3yKmfbLD2DuhHGtwBEKI8Tf6q4yH02lW2vL805VBmOw+N2YX
r4F5/awPkt20bnen0DdhxXAwLZKj88VZWG/NCQ8PrqIboICLR6nfHK2BNxRpWSfq
ojN8jQBBppPaIZ1J6z3fmeKTIQebF/6ze9eVxvwlomJe37QQcXKbTglcU5IOSFRt
oCJph0aY24UL/+5qPpuCV2hdT5sZMbdjN/uYyzDYftogh86LJDSO65C0T7VLkbYr
qXUAQcf4HNFXaKO++Ey55mwFJ/iwBVs8zTmbyyF7jzqT/qMUZev2kGwnWooFDWbR
dSbjU9hpQu6+tdoBgoIT9Czi1IOkqaxdunZZABEbKcbA9KgSQlMMAxFSlSBNi0cN
Hj4dMo+QV+0tM4TYd1reckpIbDtqNpLw0W5elqnFdqdI5tEbcAoHaMIiB5a4BK3v
9Hyw/0TO/sRwkDXsgTBEbfkaw95lIzI4ikPc8nwlDbkkocSA116dyfrtGUDXrct6
BDqgV3yxZwDtO4XnzFKmiuN2+95pEkWOcAkOXvCnKbsa9NrHlE8wLybNdxd5Sa3a
TY6tv9y1Mh7NcfmGzS9Jltbcs6Swa+OUnzN7ZahwxwqTt2U0VN8GYih67JkZCt7B
lmQsaTJlUUkIMmLDbJ21Q1QlfsWD+EGV1EmUsYyVDU0xNR4km4+NAowKUqnv6dW9
+bjDH7wunZpKQqOUc2/xfoHPUTmsqYmdSoxQnKijLbb12MuPbxiHbj/fwUgoj4qU
fR8ydEAe2LQCjohhlEJmqOwdhamefvHPYBB74OhWZdSbSjekg0nJNyXPNu1rOA0q
ogWqkcoVwdxB3f3QvaV2NV9Px3cmu+9Z3J8fT7sdiguOL/hPtq7zsEmG93THrWRI
EPVaEfbR/chdP4pVRxV9UMMRtcCgo5IrHAHdy287FIZ5JiIa9IDxwtlDK5oeL/sA
j4/VrjAlFux2FtxSTmUrV6TvwVKEoQn9Fe21x/8Y9bcP7+OAOdasfSxCxxeY1w8B
TT+DvyHgBJc8VHrul0ZvGWZAVlDNQKj8A5Z4HbGNtAgYz9Q1gGMV2LtZWpjW8E3d
qH3LLvK2VEFkaEEjsHb2aDK7tvFEpYP154FEyriveGvlPWcQFyTPd5JipEQ0g4GQ
Hw1rzFJ4N4PhxmhzR1TBqIaRnT0AISKITsPjVqolo40OvrbC6Zj1MxvIMUxuvJcY
okOuvwE2d54WEZmQVt9oEqDPdJ+Bvq74y1o1r6zPZ3ehtfASVJ8HAvW/zN1nI/dq
FnzWEVIqc0oyjx39W9bC2lbmMlEKSHZXIJnKzfs+Z2SsBZ7X6kJVYgbvYpQiJ3mZ
6uVky7hwce8gFv0eRBe/3Jj9cuD3r5rmAXSDK3WeMbaKBRGSFeusZ00RN9Z6hFMD
CSwNjq7FJAsgrt3yL+bE8Blf+nQvQNnIUBM6WBEvVOlq8YcWAU1MoKuUY5EtO2Ij
crCgQmNHUXAyjfQxNECy8vjjve9/9MeyNMgGtIMkD/KKEj/n4RVqPu3ePkfQ3lQ0
fAberSAjJwVn3Pjubz4gt9nkpggZ7mEZ+bu61AIZ0QR0dVR5SThtIyETpatCe6Kq
Hb76YcwCm+ay9D+ADSfv2ZM5R7RLDPp8F7iXiNNuNprAMaReeHAwQzPleVs87D6o
x3BkSAmMi43VnEL92GNi2OIM5mSjB3hZuTL0tIruPnKdY6lSVTusQ6/sIl5RQj+s
LH3RRwgEhKevlFkFX3vCp//8y6kj/NI1eArCHjcbzL0Zp4HRRwRAHXxY5F7JUZGs
dl9d9Mfh0bEpHc2wkxpTdn4EIFa7YNTTrDqwAyxbbjB03sms0P4AEpmlOc7nqoaF
LTIzgtP5osaKx+ttuBIfDdAIsGHBGKqmKqSTZ3LZg3eRTDOKXNqwb3FruO5QRjb6
070VAlM/2tkvDbt+at9ZJWNt+4bary7L3IB78wxyStWSK9d1TmnRIougDRifw5lq
FtMnmoeeXmjG038L9wSQX8BIfRN4wnbNMnqBDvIYYkYtOHwE4NHKIRrbzlwJlZYc
qCevIf2uwgWwld64U93xfKIm7+jilBsBlRUebIQ6ipY87rpwFXT7rIEuyl9YnfsT
Xv2B6jgdhjx9teDw1TosMwyY/RwhBMqSt+pMpGSelDgXnvEL2ofNGS5uTzOZd9mv
maS2THeRuKLhh7khv/zridVEr45c2YvNQFL7OH/79SV6MnE3LsB6amp2OGnU709c
1WRDvG3D30ujIgPlbUUKmesG8q7VEx/xWMMBG9YJBVVp5dw+EBODb/g6pEKnsQI6
4S6EZeZRq1lLjaVrPIPtX3m5YskMCo+Wux3dvyLHIhUzAiFvjYIJXlkyCQYmN5Z6
jK5NJyVKNjFcLMpi0uSDDuBtbKU2042BttWpwqft8TOgV0zoQOBcx5xQ+fzwd0fI
Nt30XbYgtJfBk10tfr7RmA2mKYx+dCxm1l0RtAKu4GwZORgvkr9e2/+Ib2N/cvco
kNncnlZe+jS7MVNJtp4vXpsNEh/moApXKolk86LimbmT02X+HmSf78vl/lXVaGLc
kbj93op/GMN32rpwMuDbfy0oyGvUrEGG9snfEEje9poYf+ktt19yuVFjfQA2ILX1
taFhxtCkU7HW55P7apbxpCsSjyc7oCxZ/LkC/5LVDzTXEJAWgzjNXu11A03NF4Li
YVayVhd1mr39QTrKkAOS+2E5+JPiChWFMvbeXvG/okiQoBRtc7uHcVZMLoMVHtNe
sEGQSy2zdJTs2yycFPo6WLy27m54vroN5O7mYw0gahU3DQjB251dhfq6gcdP7o2y
In82JuYfWIC3+WRV5nBy/3hayvsLQ+76EFMXMILIMqcsYdHjf/H/hxknOWkHnW//
uz5TkoxmcK4XX6+iSNrZlNcGnKh9j3hJJCw+h3ty9pKObJKQn4ALrAeeSk7jkZ9q
Zfw8n1iCFqxtviyjKtnQLkfrBKuu0+NAKw1FhJ7wYpZHMdmDCr9dVqtCrH7c0mc4
EgHeE+R54Gk87WKFV30SQCrCRFJBF+kLvC6/WXhnwCKRGWi7qFXRS2PEpx6N4+fJ
kX1Pfpoa+wwIjHNDVtM6e1j+CzqSaxtIQepd3Vj1DprDCHSr2QJGYT2G0yMmlPTO
6npq/1kT1m6dztfibL71Uq3DjAUoRiyGtV1b3qv1JQsTdBWSDLnb+hNeoM/oJxfn
GmE5D6QruQfhoC7LjwA1w2bDeuCTb7YFrWo6vxiiC399QNUVBhbu9A5XnsPjXDYS
FKW9aQvaL9HmrAgDStucf87G7+keRrNmZYfM8j9Nk5mqFlOcsqs5EXzKfu3crsFl
9U2udN+25gFk0A2NlAuMwVHxPeWqIhflK55+1yHiAn8LeDyG7ikDsLlW8bwjhwTd
82sM7X6JJBWCfb5bHOKl3CKqNQXnI2qCysxdruAOr8y9aZE2JxFjPdkAVEAvK3sy
YyYEogZUsEjhgy5BjqPT1kw0rfAnQueU/CApefruYJAaSWNVrJjiUTClrCbEab/y
cD6J6AQWojP0qo2pYmpgVbtPdLWBQH4vDdHD0jiWwB116Z2UnVGD7SWIu8KnlWaT
aeMHAXhd2g65/ObjkhQIu1LV0dYrInvMAJsS5xCFFLUHleSQqh7LfoUrAJsGJLJp
ZgFRnkKqAyjzWIJYGZhD+Fl4BVg9B929zy7hvELxC3wPslOpFs+he8or22QULOjd
T/XbW71rFgC3tBEC0MnYtx8yRi9m6UHiHEg0Bz9Tgd3ooWC/gge8Cpu4u0xX5MhP
uegIZn9zApN/pU0khgPKEGo2jjx/UpB5ib9WcOBTCBGf6pOlxvc/SMcjdHJfwzXN
GM9boF3Yx+quUVVW9D1tCL1wqZ+cIriF07BQXOcWIsfdJL40fO4MzfVjZVpjpLj1
RREprjxT0pINYyAu+HYr0IMi3wbv2Cb2ZQBLRsbvRKE1GbxLNOEsC4NT6REC6H0O
51OYuNn6UKU2GUBaKmoUKrja3sJazczvrkaICmt+Agg+iZy7eXLQyDqB+WB11XzQ
MOjoLENSetO/uO33UiXvDL+jw2mNVPMw38LzRD1cMOf7E6C4Uac/2SHG7U+iWp1x
wt2VJQv/fCfvtKs+aNRB9SbXt7XVvFKy9g12p8TbYoMVdWNjX1szjuumvUB9U6Wa
sRXLk1kKh4TPH6vCGgqCvYT1GH5qlz7Q4/kpwmG2KkjE1cC0ZR0Kwib+X72q3fKf
BT0WmGYOajK/haGX7sU63XAKI0hozlEh4bO6gOVbgU5LU86ZAcaatmLiRREPVrym
tKNQIyL59av+rrfpPqRKwK96MuYXs0U14SzNltATGr6YcoU88bX1QXom9re539vd
D3xRWcFh0jF0TV5YVAUpKxi8tVUpOdXBtEPiqIe/3TnpKk38fDXpVBPPf3E8/y5Y
MCsMEIai149M5F3wE9iVlO69zBwpHYv2Af52lxb4xchUJqxI2nqP1fvuCoPKOPy6
whOF0RYXQLSf4JkchMkZN/MVHG2sjmrfHyO2A8AZDrDY54H4DWyIAtYhi+piAIeZ
u01vulxKYOdZxkk1UagqNbcVIUFAOsAUMx5dxJreRQXBU2/7i0vHmAGAAAFrAexn
VUp5G2+6K8bmj0IuPiwK7cl2HE07kkLfhDDOtJe0xlXxbR+Mc7G+Eq/K90ExtNIN
b3RFhk53zPPqedr81r5m6G1LV5pbOI+C5Ge6b4iIGzMpY3NrVjLXOVuxikNH5reP
bLer6Z8+0evg2dHkxCFFwgDO9t3FbIm2d4C5YF+3uVGhA8cqfWnn7b6dOehKao5E
RE+BLAdoSHVaxYZhLEVegVz0d34+8Mrohbu4vcPuXhjHgKTgK40sTRKHHUqtu9Rw
zVrujBmG1tk3CjGZvDAyjCCwBpUJZbMqIoHD/ugmgRNK4tgti4TKFzvL5ns3sE3X
fxjH0jjOG6+isOqYjJRNglVDfZCLET0EeyRYaYtIU2Z06f4DVKL4pp2awCrCvR/O
1dNA267ScC15y2ZJsoAkhmVnPvvg1uaagfBltE/8jtvewlbw05RYIq+zacQ9K0A+
++Vv9ns1KOOAdqLIYepMVrJkhWa6cc1wAuqC6s6Jg9cgRpT7Zw8omwttF8klN/oC
hDLgjfDFwMUIzfYrBC6Zs5mJObMjMJtS1Zj3MRb95Z2OKF9P/HB0L5/Imb2JYJ/M
PQR7lyHSDpxUAI7Vyk4yDl7+8zz09HOBby1is1oqiOS25HQKZBpN9GT+WlpGS8i1
KUXRBkr5GXCkFLm224CPLgX+Z4DOGQzVgvDBGGI0feiQC3vnR9cuAGBTdZsEDdrh
PwDymDiZup9hee0QhafJNL3nAqzFbSY71M8XGDz6Wo7TBqlSZo89JWnY8jA7EK9h
y5p+hOZ4imTjcDc48aVJajzHys7s0cgVyprMQYScqQwu8h63wbMMNx9WgFSetA/t
duyw+zIx9I/j80goQn+hWOppY8pu5GnZarT9jgpCLw5pNW+gIUltBcdM5bV3d1uB
G2GwIFf5T9uheNj3Sr7/Shjd0iZ6Bq7QNm6VvIwR2jEjahoR+UPRb8gISGj+rDw5
WoY82ZiVIl9oDx+DRzES5aeODt7CHz8NyzMdkn1xvckor2xw7feaU9mDwsKwGpqq
de3H2GRp9sJn8bhWuKWTFSXtwO1ZbeSEcOs0+NG6RuvgeIoOa1xW6ISkKSTg8FMe
jUUJe0E10z/G+3tT5RDyGrnSwFXsFWK3UmJGmF05t2u66HseLolPSr22LezFFAle
xI3Nv4x86G/k+DPN8ebgspb0ety4/FUv+NtV9zJeUuyWqEsrcDH7mawfbscsYAQE
vbdC20XGC3plrcMSXSdJjs79MNugRFP39cD+GkDp/ZSJzqPdLBSHEWqhI+MX/EMs
LiVBC0ixU1zHJtDdYnpDI9vXXGpRowLRA5AZjkK7nhPpzWvgpjkv49Bapd99lLL9
BnfUPB8GT1wno3nWolniVQIOrzvgKuEiVQF/zM5VyPNQrUMsXTBU2bhFICbUgIf5
Cw/13/sgs/DHx4QlHvqZD5kczbr/TtrRCiOCpoOVM/dikP1QQ3OZdrSfG2L6Y9yK
863JrlIh67aIWQeI0rEggSqeUqLcjgScA4ZPJt6rGzgu9voe1AuMxpTR17xW4Xfz
r+ZZvt7Bdw6NASOeXkr8GBr9IAz15w/RU1+bAzPtn+w6GHCKf+qhyB8DpTKIUufz
JnlH0/CMAJ9r8irsVzVzcyU7FAkAB5HfbrfMHn0S4dVcJf5wJDkGBbcbma1088GN
VmTRuwXS/wOqfACR//9THvvpLdBNHNYbygFdybC/McgJRQbnNUr6AuCmllSDryEk
GpbbtKhwcN6kNXE+oBGl/N7YmgQXnq8R5iuE9lca8CcGiyryQtIRkA2yEdP6c5pi
B4O4WouWOxzYLPEMYQ8f1cFlts96oWon4PMuQwC0357lO+HoC/GLp2kH8jmdOpcT
zbt3Qi+MPGWxZ2ORG1KLM7Id9g9V7+rxa8A0mGW4LE99Mo1TNJcSP7n0CDJd+Mgc
ofWs++BB/4gFBkiXVBeuD7+J88AOw71jth6pTFLfRB33YndmUH/8Gi64YikQcvn5
Yd7cY9cGVwfxBZnkXxlv8QVaDLoWFU4kVlZ3PcfCEYUeV43j2xxRrX3Egjwj1m1J
mzgX5rclMVgfzn2DFN0B0CM5Uvj4DTyye1o9Hht+MZuWtP/6NbR2+0VjD5G70VkF
v/FmlWYMBJE1FgLJDMBVM6VyD0hmezdEIhJuBd1sVR3XSPhy/vzPCDGwcvY7XBoA
p6dzcRRfxIFxomEC6eRfWP29KD/9OxsPlaBeudNr5CtFuEaKj56tdtTXrguQKTKG
TUNMzm1pBvIBoxUPEGg51Fvhlr02S6lDL+TBHPM5+YffJ5KshWo/W8N/1RnMub1s
Nj3tZmE+ZJWo0LETr5JcMXkBBja8FrA36ev6hB6GC1dwJbi+5llasDIfVF+wosWB
qlyNjpkQzjLfZ02zu8q+6cZJdVMy5fl+emZM2C3Lx6fzPikYZRddJaWjUMA4wef3
lEWazGLv4XYI7Wjq5/wFV4lQrNNpCgzy2XRq44S3Eod9LdwODMQyE1gctPQrJf/0
ji8nbxFbGuIezw7mNNGh1w4VWSdLNYu9wz/+xiiddcat8ujGxpwNz2UnJ+YXDh67
Naz7tfWsDP6dT92nvIFAxhpFTl0kwkvn3pJqzfdRN9ywH4zgyQ34AWr7SYKAX/B6
S24tMdy38e0JNZZ4IXh9GK9+KbTBrhCs6R1R6MmYwoHh0QYqbuRyYMR/p8uzbkq/
6BaqCFRi1C/J8B7XqFl1fPA3pmYI0DhCz9cCCK4/OO6v3fGmec6vMIVDC0MLfvRt
2azk91pOG+p9ETLGa/T7aXjgeHYka2s7asqC2q3CkLXh3FIpdHlBUq39S+9Q/pe0
0luFjIYifhrcT4ZK2U3MRCi0O3fgpD8b2qjhGN6mhg1IFC3hUf6n6YE6B50VgsY0
TKQfmWR8hg4qn/ThvaKcMhJ2SfeNkxIVUQW+dndl17yKD8zMwf8kKYAD7hNHtK26
hUjf1aAwF3FB/Hen7h4TP6rcQFXDdzxeOiA12x9sH3dREyUUHpJ+6zdv/nDCldGG
TVF/IXzkU8NhYjJlDvsILf3xczcsocRA76oxxlI5n6RmqAr49Ih4OZgrX0BouxCU
P6e1A/b0zyTTh9yjyuSpB27b5oOs14VdgeHMCh8xNC87nro1p1QPB69NrRfVijTZ
2tN9j7szjGDw9TGl/m2F+f3nr8PC3aH7gMFKe/qQ5aPlom2MTNAA7V0xyERXZJDi
+vHauKsY8FA+EqMuoGHuk2yuSNlWInd3dfJwUxDeTiYv0hxOaHZ+fppeNHUARoTW
gsC1EifvBM6Qw7V/F1NHDvTl9rZXN6WfM15MibscdLsOgAQOt8YA7Fv/QpGYe08i
lXi1ZA8n8GDv2oZHqhU5v70cARoREvIgHmjU0/XFpJZey7/87wvdlEKKD8VVFfok
7kKhhnFrpgVbiBWY6VCLzuM4faWDpT64vsQXOJejfAZNgQ0F8qq10Qd1p4KTLdLI
xyeXx4Ovn8hMdxGJRix+fBkWx5qGxbSaFxWNLEfzNuuUl0CKqJPNHWaRjSCD4sgF
4iBDpZBRC6t62/WHkFeycDcZpq3Q/P0eUfRhB7p57q36mH7podUTeRigI7SKSR6w
HuaM+pyE6FBEEJmfhs7atY4/zqus0rFQq4Tw4v1bLnyvALE6ji9GET+ochgolKka
OyDfrsKAThJd4kc3ZVdKF22xi9IaT+lAnQdUqhEkLIS6zHcmwALlqlq2JMKM5I/J
wX3LdZs9e8tMhmSycIzVL5I7YCfGGZBuf9dk24XyJ4A6USJ9X52aI9EqbmgR1/fG
OT89Df/CckW58xw0SZPZeKc+Hvoo8qNyGhwMFDVncm3+1bpmxZaCELRH0gGQ2+yB
B14sZPItCzA9B7PLx7ze0nlxDTxHdtZSwb9PjzP7/2qKguAsMcqYaIEqMBUjKoZb
9HS+/YeSX2gbTg1yUvL4pI2HATW5NFn3pOuAkQuQ6bnJz3KsR+4F33dLyTULf9Mg
RaZH5qb+15q94Uy67psMmLplQbxApEsW4NMSaTI8VBE/s24/3h/N1q/nlTY6y9Zq
XpEyAmIYHAeXfuRsw7AJUg+mScgLhbtf0Z69nB/OqzNrrkVqe6aGAHvPUgrkg/pq
XOoyCl9Ppcc2rc0mdQ2CGSK7vNjmOuc8iJUWerGGX3UGQL9I9OsfxfwHVu3ugAAK
0HRc2zTSxUCjvBFyq1T/8VtBF58nDh/oxB82gmnNu50QLg5/6c7NgQvfz07Ba/8s
Eelz0fSdabiU4msMBLigi/esApS88XP2BGopaZJKw3EfWcXj4QMgm3GNwgnEG7JZ
E9p8n9b0FGKxZDQyOxZEAF1rHRlAX96RICOfdeK72FAgHwXQQnkm7rZL/MkRKCkR
JRVow8ui8q0sJp5OZO0R4jNRTPplH2SOYwKQ+CqysIKtMfgVWjdjCNRT2Yz9Vqd7
n+DS4SY0Q9QS4lDTuScw1LR+sKBL6nzIAxUnatMuKYkdXK85oIRMY1uYkjaJnv/W
JL8dh7CuxRFYZhOTdJ7oObrcxJFO9tlJL/KjQkYVnpEFqsUDzjel3vpj7emQBkOW
izxAYx+ZqcoQjf5YAZ3h5NQWgc1GQyOcOmfaqcqLkIGow7LmtugIvrZ96zhhMDZi
G+eyqOWTXYyWcGMn5lf66yGYjTFe+mIH/MSQ5hxkwGRyoSAuRoLM2gCLZyXtOQ/q
b0ixVT0YGLlWfe6avdDC7dhkRlGV7Ek9BW1FytNYiXBWmRSledklom2yzOENL8SD
idXnw9RrUZCntuWQ5KXuts/U3ZCLvt+6yjqaXK70yklE20XMpGAOiNMhlzHSDLiZ
5F29RM4RQ/USg/t69i7ntv2lvjUIobRtDoSIl1pFIbXhyMJtLEOYQPwGgm3G0El/
Pe/25gkSuUhgyDY+jRTU1+WKSsTTTCUwdDiV/Wymai8XegcI4Baouab8J8O7Dtjb
r46nuSUYWEiQqqwzR4gyMevkDEhvqkKOX/vkHhPexWP+sUDMmnzKKo3D3buK7z+R
IjSq+4lNq8yl1wJguSD+2RP2D4dtTzNKtxgmoqqjupcepp87Fl3101RKJuXNNvNM
tCrFZ14/xyZH7bvWONLY/+Ew6HaPCvzSjZDgBI6YygP7YnUOmvrgkQaqDGtgdWT0
bFgBmfpUtpK+kwS8FSiWaiasOFT4MJoWu2CublVaxNsee7cde5HE33lk3UGHCy6Z
ZIZX7eLYAUcHKgdft+5zeG6keCGowh/W4rYwZTkVbks/E9rCnWju7SaHDkWT7KJE
LQ1MAmOsOn1Haj67pb0IrTIhruGHUMasQeATSjfAEzZfNgqXW7eYxdOAQoBZZtKN
sl7tVuv39WEFuURY8O1+nb8c/jmis6pJZVL9zIkPbu7NeW6FQHB5ASOdopwft+CD
WB2y6/mJICd0M8iugjrYZlYGnlC4x10mpO2ZhPQ6gTEeKyb0QsrgrWXjcPaRXLrx
5WjsHmc0mI8AFOI3MOohfp4XX/g1H8CpcSV0YJMpvScxKPyTz19LHIYPZTFYlq9r
RU4ij5jCuJ1AqhQjkBgX2G5Zo0/K49ZPH3cr+im5OBop4vODsvWj0lc2BiOYz3su
+n1kZmhgkIyvlF0fihPgtF/ueShXgMjhK2Ercx1tw9f/fcv9GwFjwqziv2v3DaSm
Bp+OpkG+W6BDOegBi3SI0oBRCiuXOcuwsLVp9CZukR9T2oINXSOlEKGRXVREbaf0
Z8qTtvMa4tiiIfi04VuXzM6aRAPU1cAXSlDqM+tGBxBePj8LykcmPoKR4YbnXqMd
h72y0tEjM2iZSnS6xyEmi/SzI6LUxlt1lI0Uzo292NynDlCS693+spGJJ+jkfXf2
pKXW8dVKb8fO3oPgg0Q5IoOF02LwTRBsU0MBkcRq9OjGszATRwhYPU4vINC53nms
8loXOjFE/Cq7W+jL0KrMtjQdzKFAOujnLD4nq+YxB+cFHKghBPfTs9pAEQJJVbpu
7B9BOm2Qlt2xQvmDKTVjYwqHdaGED1PR5uSCZ4A8kffyPHXGQO7yfPh9ASy4W44q
jdCJLK20RwMAukDnHbAl3fYI/aVuc7ssoPQOK3aYbxZGeTXGRpTxjDLE2AZXpG/B
pHaXZIKAd9fPANVih5E96btqRsvSRCMnmO7FsH3ryhQzJGRavMD/sTvPTA1m98O+
gDhzS510tNtu5/7ATNfsxTrJN67DOcWkSGd9+K1dZLl3Wu2CneMeoLiSYc9gTedk
Ur9GivBNfeKgzvr1v8Co7wMavoG4YhH6XUaeXPzjW7grB1LfZzmwMjG5/c2G78j/
mGAh5/rhVA7hGmtsTxJyTOjAY9yweS/PbBYaKM4poR4zrmX0YdKYdLaLGpq6NwBz
Dwt2TBX9kfrqO9rieVMA16oSTrWTXqJVdYaL6rwxvbiD+sef9R13pNzzrotnG+Ty
z83+WbAXJCS/36jXKV5/QBnP8L17dmOITbi/V4c4v95e9V/lTtaWBeidEzUn85AX
7EbwMtygJq+U4tyHrBfU0Jzm0tD5wXrTYqlJ2Fcn+TSZ9OnwyzuF3K5CBD6wR9yk
IYcKpJxO0FPRZuSfDHuFjzY1iRitsm7JFwP/69JlUOJ340Ku5a4YirG8V7sHbgPt
OHhBtwx/YTk4W1aPK8lr4cgy0RM/1ameV2PIeQyNFlykzM9Ux+Fjul3c1FI9huIe
bfSj0LWVTUBzXcKkpgbnSyxMNjuu1Yy36Lxaq+WuyrohRDCq80s9+lTTsF/u42h3
W9LoL+PSUiHmUGAad80cXnmgyZ3wZi/UDpzoDBkCsB4rlNV3If1dfNZlbGBO68+v
9xVnlUWzQLzZjW7P4XcJ2MYAJJN2w+2YH0SxchKaN3dum880eLzrouuIvgtYZFn6
hWbhazhkn3BcFR9/eWKubPUlDIFMHu8s/1HM+W6EKTNX9iekLR/xEsAE4PKn7wY9
p06oMPEyLWidkffz6cf1yetuDyRhaIs7ct2/F5U9Y6tDN5OsHIXPRTyOLfdPFxl8
Tqd2FPD3JVZLjN/3Y+31bPu4GWTsU/uHHOMTlF4h+GFmtlmk8iADWNgtWsN04Kjq
fUgL9m705y2vLV916BT1V/ChNF+CCTg6D2mXRmwHKiNf5G5+y6m9wNuQaNMcK8UH
z5UAfxgU12YBC/11t74U0g4m+T2Tq0O1mH4e4hCh/NbdnNhmdtennsGQJ09cBSpW
+GqklbKrwQwe7dzzKNsovqUlnyfH5cKNEcfb7W617Z/gOMEeHKn0cwjEdzdUmUMK
3XxCikcZfDu5dhzsCumzzx864IZ/ve0bXU3PNde9zNmH9IbBZpkJ8wv99DAiMgZd
bgvsSZWQE8afz9pivzGNr5MYOITnE18eRTfZq4GjX7FHxse/GyoSS2cxGQofLx8b
8in6F1SaCaK9sG4nnBRQ6KUOKnGFRJZ2+2Scimdulm/eUn6gqCpbtoR00ZpXDRJo
Nk20mIb6rpizBRHEs93gmI82LiPlaXuvOZhQz6e43Rioi6w/yJwHgSz2nmN0suBg
xSlUeKm/BrP6sbvoVTpmV338tRH3NqRiMOuvoKDdoLBMfyOfGg5LriWZjEEBuuBz
BwZ5HqrB9SEIEY48ibTx5SgJoYut6raSNxl+ozM05HPbBMw53EwFZqNYEkNXJawc
iseSzWmAg2rPGRXryGSJbcG8TaZmKoqQr38PJ99vKZQrNV05HQzY5S5C/GooV4AZ
Veqa9a16pc8PqJwkcQ0oZXLE2D7N2DO/8mqqeE+p+lqWVshcdUzOl+dMa18aOo3B
Rr8BYpTDsiRjOnw+mT0CRVo4ZwL7Ca6+jNpvYOXknHT6qpWj8gbQaWg2v6ByyNIo
/zCjOFTMEz4pSv3umcLfb9XhACEruCtw8Wzft/afb1y0mz+JlxtE6pBBEhynQ1Ew
x6xSiTw+Lll+9hTE/4S8VCIP2g6u9FiweWGmoZw9za0N1vFrF/jUpK2TWDj6g1Un
QgcSeeKdOQCSqWdR9AK2RQ8V2+KtF3WttFIJJ8vc2GtoS5LNoColUMMlxqwgN+lT
wJrCkW48YljWPHXD+Uqi5kRYm5VF6Z2lvgHRA/4J3pvrvgxCs2gHJBHOC389ATaD
hBoiJ7WIrdOKDSeSHomrD1jqVniwtHpYglZsdcvyndkcl0jIMbVP5XMPde3Kokin
FcDdtS3sVQkG9jaZmU+KUcP04pVs47AJJ1Agk0cxv4zwA7Xpt8tPASrUlhsX3VBX
PIvkXB1TWiVqsXQ4V2a7ry6o79fSS54/cZGH/hHlPgTGpaac9ZhsAl3rOXXO5Sd2
oyCI29P5pXUW9cncP69gj6zVVj8NATHLLYsO0HZIrTi+z8Hd7XsaYiCjHUghGsPf
fNBrXB+j+ra0ZHoWoPOmk6R0bolCkwESniCD6o0t6+x0r3V8HNFTzcJ/s0j8A8RN
SNss/SioUXflQ8G1Ej4zYFxgFya5zDOrusD1IbWUtroK2Xt2x14mwGZFaz+VRAHG
DKbCEmmqR+5UgydfL4MbkttDB9eH5TPKLBJOLXajldlATOzTRSjVuY7PXrt0Bq8H
IYVz3MZWPCq3MYqZv8vPUv3Ad2HnzZS/czjc0yB2uQxNik5Un26tjKoeyHnJSSjR
2uWLrTbyXkl1ugT1B2hCd9TFPEBIDIaupYxfGB/eD5+sOcaTALmolweFn6Tn3hCp
Y7Bin0YxHjM7OlsD5amrApBOamnc1OEkGHCdPnFut2omLZG1rZr/aUGfYthZ3su4
z/yj86d5PS98DOt78PVm0wab4JvzreEJrTjOwT/XJBe+sCLgvVNl5gNGf+J6q/ZH
HiS50wR4QTo7t5s4vcHPdSLx3+pYyT8Y4ZdA1rxTbFoq7wHOon0u4REUKZRLSYjF
3wzvoMeCWK9BjS58ADu/PTvyBGBvsIpvry6qJjIsePdHLqvXDkue7MsfHjzfukHT
sE+zmC2ksNd6v25VEBwxbW9rCv2RWW6++fsAcMX9JusppS6cLzG9NwV6fSPT4yjU
0MhDy4nwDfCFKYEezmnlgE8+CtEiC6LuX0ORX2fI1459rBZySOcHmr6fWuAPvXc5
rysd18sao/BcUVcR1HxuepLatVFoqEdBM0a9CX3wfUdIelj+w539PGJw0afCIR2k
/cTMtIlsfecDH99fy48Z3K2UKW6MJV0yej4I5ZXfwlDhFiDsuNYlCUn6i4z7B5Ke
+/VIt21TE0EnY+IuZ7F7321dJmCx4zJ9V2/8djrkk2htslDiV54pV0MBKH93zT8+
WCigcTPyW/xd2EQNwR73oFSPPXsffuxJcg8Se7yyg538g2NvxeqvOYWYPkPbSdbs
bvz8nUSpwXIpHRIJT5HC1ixkLa9s/IkvXDTupgRY0NqrK62FwEYnzw5f151bVS/Q
HZIAq2vfRH35S5AG8/szViP454S4ZfCIbaNXQylfr1qHrhxKyAYH9aOFREMuZnuA
PGMuH8TJANDhjGVPIUhtSaUF56XvTpOWXNMw5lGxWaMxSLOMPgK2/3QjXOAWe7wb
lbdZxsNAZOCZ9JRd7eZQ1whl+AJsmBtP4Oo0eswdr7lC13dzLdb2B/BODHVU2kiO
QzkRxOr5QPv6canUx5TPE+Wfitdg+mKYoc7gLnvW93pXXJewEOGNIm2h090KSmXU
/67L+HJbkHv9uFmv21lMzYVx8z3+WhDMFzII7q/OhAvJlNiGCPrqMOSXYldcpjJ6
uMmHZ8+wY1er+WOyrKvjAzOUAkoA2fWo6Y3Iqo+lEbpgdDxmeoKk/ibq+M/+s4Ug
oYDQjV9mjwuAI+84g65HDcZRv9nqHnmfTuQmNp0mA+KJYfVHCV2Gom64JtQNx4qR
p6MF1wTG+5r0jGcWjtPrZbTtuRGBlFxyf1NsR4H6KS5uhUhTCW9cb3q7me9W2ueh
xOOWZYzcYSG0i7YSXRxrdqpk4o3a7AUMtVHwrCWyF3qMRD3qycO9A86Eu2n6fzZa
ht4x/VFSJaXKmLDtjbS9MMtyTJLWW9njtWtJRrSaUSUs+T1PwNDxkvP3r7889mEM
PfosZKedswUrK2wn8cKehlpw4reBY6uchTDBGPWPShatmKd1mUWxboQHNtCw81kJ
lywgD9T3b56cOqMIcjW+19YYUU1/Rbigl+6wrmvkgBwBrbS8Qts3qMY5vlLwdqrU
KuVmv8QaQHgoAAjzcegZKaRufeyFWqUhfevm5r8r8wRKtRrfwRBf0zPWNkuAw/9o
Xhm4iHTVN76SlterEzeTMUCRsWtcjgZW1wFeqzgG6OtUtMUP7geFa8S3XCdcZMR7
4crnof5SgMbCZH3/oorf/OgXqRcUROTGYRo171PJJ9sLoFEyEYX8snZwhQQbfOfZ
GhnUvnJ3m3npLaw/s25Z1u9eQKFKkz52qi8O6+EiAZOZZ6nrJ8IRXtqH/qnWnjKw
tzivekHp2TUOqdLohCfxC1X1yUcTW7y4Fhfp35qhgVAH6w37eXemt4o9Qe7O7/zB
2Ss7YqFGKcYFH24vtFXrg1OfrbBC6+A7Ck7dAtfRZ/HyQCOMo4Ftxm2rZg7MB5x+
mVpW0Q+XGxI0q+Hspxew5o+ahv9oWi4eLmNtL2vfg14ez2WfYElW88QhXzNpxOYC
L2J5jZHhNK2ZBw9U5z9P3pEJHdJzC0mDXLluzK6d0Q5cVj8mhOynI0uvF6ayAu9y
JNpuEmvEpo0P1ZZ81ZVZkrDwUrIqhCzCxsadk9jwBiMPK3DK5eT8Wf1UOM9f4vce
4oG3JS6KpcgvOuutd9qbY6mHwOR7U/YDZEXvM4mXduwhqpGl+XLPMyefdVvl55B+
9/C0EIGV334PEib/gg1yF43m3i4ZLUN5tvf5hY28Z9ceMHC+th60kAqrHjTA6Inc
ake6WdD7GuRJkUJtkTF/F2zSL3MQa/ikSRqZv3cJDAOYHrmw5UJ1E7oUKt5iooSI
Lzwu/o+M2Tih17EBiPuTM9EjSa1OUvnunTLH2efR4JXGAv4HxchJNlboAAIIgg3C
8+ZNZbIucUxE+N9A7YFHyg0ppvNXW5hJoO0mCTUYZQy8xqc3NhAOzqXlLX+gKQx+
djQwE3rlabdkewZbAnhzRpjaY1OpmkQOlzanMc9/M06iKqIaH1TE0qQHD2WHc6sq
/Inp9r0LRMM0a723SY48+sO9/E9BKx2g8UJZAVjUw3egQNlcqr2LD//gXOWFglwc
2AA5s5Dwo2GuEJ+nXWyFOp2R/gNUvEgu7ojaisvK+LOg5HUNEZFD+pGCc3auMaZt
LJk2BMAjR/IEIXm5Dxiv0LX1FzCVM0rIeBO28Q4Nbvs55sJfndGRif+tUZu4pIcV
vxvQTMJACzFxxi2b+hI9N7zhwwSJ2oCs8UcNG1OWttDB2xtNvfyU0UvNdd4NGN8i
fzCQHazS62UOP4LIG1c3UXPRKnmqYQ8/E8JygziapsuPQdVTPgDjkFEFWvcmHbUC
EPFDzugI1uA8vRvZzz3c47Q0pQ29WLh2PcrUAmyNGYzPvOwj/W7Ik2HUenuMp/WP
EhG1/EIe4QQIRZFrqlTD5Y/qYkWWGD6+HrG7goIsAnLdycfTi5+UlM0hdnu2X6yg
Ur+J8hqj+y1U3vNQ43ugd5SR0ncoMTPUtAR2uFpddBpMPEbucPdMoCH4iGydK5DM
rlq05tLaS4gWQRoD5VSyVFz4xrDCDvLaqI62BRLWyneDmDkfhx0C9XOPRBsPX+vx
PlJboPD4PXv6V29JcWF5EDaLoTGfh9KP9jnv8N0cXZvVkgRsO+LC/OvpXd1VyAjo
XUDiASvVMad2IRWeRfL3XzXgDmoP3tp/LKUHbxv41huzkVhj07Qs/v94vApGpxJx
DBk9nmI1giqPVu1A5HZgEbOScuH4AWv2I/oWmDwOnTeARMcvl3fq/NRr5XBfytnS
MVtnZDSqpZPtendDSfkh+G0B86cOy4luF9o2o/snsdiH1v+tHFEWjimFsGJ5QOug
7R81opTZ/F7HMRtftMDZjrOFzONH4AAFaL3IJluGM1tY4TnTbLKObQhhMwSd//Y/
PB/qO3n6GXSjaVdoYKiozI/8ha+aCiEYOqYJmJhQFBzMXu1dWB/3TicuCxG8nq5K
xL/FyHXK2UJaJRu6v4Spi2JEspZSWruAKjrlkrUwRuXumJ44XkKJ91QkB6QePhnd
1z+8xZPLWE8+vj8wXE1CrbvTyUKQbNKB/Fomq5hl7CIErd1htiA/0py0f2l6m42M
TaVxDcr4Ec05NJVMEwx5g1YakXbqKCuk74y5pOG5kurRtZICJZ2yvpaCAVGv2HRN
aIOX056uQn6OR0ZLXIO5DlbImuXV11Xq2Z7haNSz5uT5GPlBf+cxbUynRWNTikDg
vKqSS1hoQeDKuBMh8CsnIUQGNAm5p9Mb+isnC9QIjNx3c0H2NFBAQt3So0S+EMit
zl62cancEZCEVApSV2Fb890llVGH6TfnI7N2RjJe/8+v9Q085PYLh+RK0F0tDUW+
jQCVqCzz5wHsYaoPyYHK8RdYEGPyb97SKQlq9KzYd9wSVusIwnxBIa+KiByXEnH6
+iKTF5yr3SFnDKlZlewZTHrVw8u4/WbjDn6djCKnq7MVwjFqxqBdYJD036kNcrw3
MpZMD6AAxg7WUO7eC2MatPlAxpQHEpScg76oCEt3DpngCSddqIsCvF6JtnR8GTs6
9/wluOdWKa6YKFLlK1EOLmcAY3PnpbjxEmmP69879wgngvZtjMc9VK1JgOqxxm2+
zAKH2ESXfjsqztLU3l7zrxOS+V+xqlvgGA0KK8FvCvEvMjDuEb90XhXn4SjN/loy
3Z6QCXtrkP7C4X5nVVBH8GPyFl0FW3S4LidREAWl9eQjP2HPcF1ZOozFgRZ4iNjF
Rcr5jZ659onSBOWAxh8LQBNjz5OaRnhM0PB7MwZ3szq6yZKGaa0hTRzZ8Cf5Fut0
uoN/TBDsA9pHMbylQ+dWxqGAoqAnCGFVPHuz1AChn2bsVJzQ8xu1zDUFFnuE7AHH
a/CM/9bUhYHVvUC7KVN7zMQOAkfW0CE2ZnglsFtL7LDWZwuGLDwA88KOBMCn2Cfr
lnri0+GJ6XkTtTKjCcjuRxc+JfkI3aSARe6O5ZOotk1PWEi/EWBAfrO6l1dYWDft
MlEZVHRjUq6T25O7F/Q6/c0sTgBDy2Tp/JhyH6tcmbfh2cm1XrY714iffAdJA9MB
f6zcjHn+AiDFILSIdUkiZaqmCmFWSEjZRqe2nwj2fjZgN8aVv1rQ2kj8EwwXpdfL
4SJzCbSDtIONU9qS81JtHyKSQOIhOL/Tll9uI6cM70ak84DXp8oPppzU6+2OgRSC
sbtlSGwaz8OFZ+4SlCAVZe4IlFBCrU7hPRcSYgGJfnl1u9tMNj5YLMl6C/5JOn1R
4g+lcfv4cxDWwv5ZF0PtAs+M679BtRd506BaZMQFLjtiZZ0nGVaR44NQpovdBnFH
syNu8UOCS9fKD7pqsTj7PTMvekYu6W0lhAYz3N0st/gu06xVW0r5T4lufFcIIaSL
davxBo5scpqlgMlIT5VQxLe0cSMFr/qJAtIWgsD68MZuwl5B26uTGIcUAeJC27HR
QwEnsAPUdvqcpSOFH6puKIBYikOCWRbG8MjJip0ytZEcJc3qANMzixOxHdAbwWQX
HtIzSYru3bfDP7lc14CU4PylCgJpIlT0FMvgKfHd2mZpsqrGzOkxeFzvsrG22Mro
vNKzwB9XhM5l5+m7+nAVWXMqv1+zuywgWVEEg+8Q9TFqX/c3qNnW0ZgKLTDiiZgq
mB5ZzU5t2On1g6JHGI73g7URhMEEUfeTVWA1bsu7wPQdWtQW6do9+aM/vPaeDwMj
AHL6erijlA9KpG/IaFg2Gk+X4qOegzJgObR4PbCOj+4dO8t0toYxywpmgN17bSoT
V3B459rN7pEPZlKUToGWvRReVUrpfqFYyeNzh1K/zgKQDVQaiGHEqG3B9M06rXUg
FbNZj7f5JVDw9O+bREwJH6SKqDUSwoau8CcOA3GKLHHpRHo/yVdstKFluqiHrkA9
HMsGelEEA8yrr+adgX3U27f7Yh4o3Iy37NKq9MPcpXOGCUPguh3ZAQLGoF660TqN
u8qQWsrwFOUEWyndQFQf72GhzkUPLaINjubAAhzMHqqeeOcPtkJuL/TwB0p5qKD/
EdQLPLw715dDqF8b4kVtUCsuKgn0u4D1HwCHYO5Xo8q+h7CKJDOwCfrYwUtqbanz
gV5hEiceJtHDlgpbdD9uzhSbm6QQ9DK539LUsym/w4ZlsPMozfkaYyBNZILLZWXb
LMU9lCU64VeOc9sVKrBocdgl8gtJOSRF0tgfD+/pXuMRL6W52KMrGHZoB+WEx0wl
OCwNDDfWAjWffWKb37J4iBpvP0SW6u/tQim4MWpALdZLKGOOyg2/DegOopO+iWU0
FRFacCi86lJk9F572rETylRhoYs5/mHksuINVCpAltPpOT8nVAWbVdZGTj40Mf5b
ViL+fhPEhJznHHQ7Bgxu4vtpw0n/Mj24gQzUTFW5P9Ym58Kcl/DdalAGHMktoVHB
c/SaO7UwXwFJqCsTOlOQO861aAy0uRNGHI+P86N6xVq473I02mwuLxawLhG8y4rj
vwSpLZ8590oekDhfbZxYmx8bJcOnTJsKr+DCwQCSJyS+x5m3YLTgpb02XaMf+ydi
Pd7ew/TKWzAOxVHUr63eYHZGhbpwMDoUebX21zWxnQmSy0LKlIQ+BhINCAQcporX
1Ptqw82GSsAUdXNt4FpPt89IAQMOVMSGqoTmbCXdqwhuE8ubO9lb+b6ZH2vwXGQA
doN9dGOcNvxGLGLEGGrxQro2CHxm+Esi2k2n5KKNNOuDw+y5s5ZOlQ6qGaw3P6sh
XrKC+ieh66NbUaZ1fLj5DNDNsIaN/MG1mz0ZNeb5vZVJ9gRA7zYKcNHpt6oWRxrY
1QdfI2ST1ov/QEwexY6og9ejkt5NHlkVRGPGmvhGYySp4nKep7oGIx+R8ar6WtDc
vQkQcRutdK6bBi9g/tOws3eR1Dqr7BqnR3d5BKUUY6qqBie4aXTvVw9DEYW05Iwi
oaL1Ov6lu1sgQU7vbxG8lT5i7oQfp9K6QZP8u5nt1a+GTmDI9aGYx1Yb2I3Jv4vU
mSoH7N8WX1a4jYfimL0PTE8tUYZAe38Xh8RmLlfSSyAwjBUh+a9+B14663oYYmWj
HCNptQZAGWmNJrQtJa0MhrUuH9NaC1dfyo/tLuivKl+rt6oEbC0lFyI24dYeDNTZ
18iuRLZQSmRS3opHA5yJp6SXmTQzgyNAFIKUdRHiCHUBd5M68fSs+ZaWEAQvPvXk
Rl+5OukQX2WTMavD6LwOJ6JSDS8NVQtK50TezoloojaH+cBWuKW5IdHVdj3MkU6b
MsqDJBMPY0jWeb5swSAspSU6GTDVClF2bzL4H7Sm7fN8QkO2sDePPyQqCKCepHHt
XkkXZexbgK9hDTxnKrTZI2WEoOCCEzKz/G50+NRrohCaWLhZY1sTMSYSfIP+MDPu
9rDuaEBjASbVayqaYRp0uXGNsEz9Oa5Cbg1cxRJZ4vrDDHQge3bS7ln+w/ZkNHad
nZD7uLYczb/7QCqlWHwsvOL+WlwBDoyochLsKOaNY+kUSwwL+9NvvN/5NIDWMLnW
2LRlLecgfdhu5TZ7Dft5Em2GkFUncphtH/+aE+5cHg4KhWQI55/ULe1V8HhmpFsg
IrsNDAlJ45lUjouVv4j9Ln+Nc65MeQl1ll6iLzVCKCaNL1ScX7qTBy+xdJx8iw/5
qRva7qMCdXAfoVw2pZG8F7x0MxLs7S8bh8iJe1vIo1hESxKw92UXPQSky8kw1Mhf
tpFOBnJcWO6Tyy+8zS5Tu66wro5dsKYo/CGJjexbKpbciYgrsqj9wNwA/zSsIfyl
Ahc3UujXnxqxZSZ7PpLwTRbtiiCLS8PbglwKk4GPuoiUlDOgAEQH+hsuAArKCgJE
oyNx0XQ7HnXl/V+tamMHcVde5jON3XJfXyznFqJIkEinymgVOTED47JKreAahu3W
tVhCKhrvzRoMdJPRfF7a+ZUM5SV0PB7aVxWBvUI28nCHnKJpUV7yjwwvcoce7DMT
wDlxbWHQTdd7Zmv2d66bpCLge+UVIhfjzM98+dig2uzOhrp6tQ/hvA1kU9nI5L+E
3aEc11MGn+IVByJ8VqWbHzWG66Xx9FV/s9cYG8xh3ZffCEVMZGkaPupjhAzpScm2
xvEa/p1csIhAPNL6XG8U4b/bbsqQNugWLBpU5Q8O/lG6Ttk9bIt/OWoAWvCEFX6m
Ys1wX/KXKpyhahi90KIXy2VwVVA3gRQf6Vt0mOnkHm3boBh2gESXX/O+LbjOdwd3
eUimn/hEDRhhG406MVb82qd3S9uNUrrSArFY54e5mYvIvNo97ziwmBIkZ55GRzsh
p56mXTu/FPGJAMwE+79cJGKyVsp3jW0p8qtOAm8dn0VzAvyNX/9Lztwyscgj0zFV
4rM0WiXulroV40XvebSpAdI8QDrhgidAZv+/MNrQpPVQeDFd6CCjgcayjVL2cwFi
vhGtMSnFS3ZbyIJLMuLyXUEKtI10JdRbUvtQkGUooTaQVCR4emSPT+HLRnXjCEEo
Np9qi65/dmM2FvUoG5g9l1Jjd4k2lIgPiGkkX4HIam8sYpivPY3dk0LCU7Ud14Dw
8h4ud1C+c1kUs5llfq3/B1sS/Jwwx0StQluiD/s5B/mMDvzDWqTH5BbHtTsoYDLu
I6ZrLwubjzV/IK2czQoQCL2mEB3NfklT4nPR2VT3EYvlgjRI29VWjXuUKd82d13T
WZLUoyNHGOZJAPye8+/YfztxGscm3gYWS9xgpyiVx0vHmwe9tqpKcV2q8oxQqbSN
EIiu2Ix0rjV3/4rMOGcQYDdBW8pBZm1vIqO+afADJ+hUMVDhjcb54N5iSS2sGtQp
zkijo7h1dnYejUzRue9n8JDwXgcJlovhBYcXVmkzBwzpOn48nBI10c5WapmgkWcq
OWL4irx9QY7MBhDmzHeNSl9DI86G1TeLZ+KiWBeqf/AAMl9EgG0G7qE4dSdv0nSr
LSiC33EcbCaYBh0S6r+jr4VgZKjZ22wkoowUJ71XUg7K/+Fg+wSJcrEadQ+5YylC
8AJGi4IzBojGxnos4E+w+9eq1gvKOcTJcWeRgFxMpNxm74WBS6Sk/q4nvkOUm3UI
TpCZAZqhJuKCIIgF1oDkH622ivi20GMq2FTRhjNHeW9yZkLJevCPenTjXJo4NwbV
t2eLo0ryemOHiVbBAxvv8RK/p6RPH2F6PbwSMcGHCO4OM2EIn5/Sx2KtrPjt75Ou
1JazAMGtIcRFUbg9oBTLlwH2v+pI95X3/opFMn+BSEAm+rvyP/Vin55+HdPCezP9
MMnY8anjBNLkIuqZRm6P/VygoGH2JGVr1DFytbyflYJ9NI/+C9V3rDeOTNNlb7M4
FvpTpAXO2r5SWMdMBIAmuLsI4GE+xeD78+YAQzdNCK6ZocXSdwmpthnBkFaLwjPb
Eky1i2q9srBXhLopnL+nXq/pBJJlIyki2r0NKYwdEDqiz4FJdGnI0WqlU5VcWX1q
gYuz+fugk/Gcc6e03ehb61O919+JtHi6GkmyD8+o4AH4nzyvGUNOVSbggC5nu2Cb
LVBMVSoohX2GlNmTF/kvMjvTdLn16KZGMZBMMGNl2AL1gjlv2NLGKOSueUVcB1H0
JvAOAVGgbErUTDmX1C08V/evRFTW+IS+FQT1JqZKE37lxoY/tff7vhYfnIEu2gqp
Xg84k3zRoWirCpsMM3nJHpM1dR62FzC5Cp9z1LwYMbb9QhSkJgPCv4b0YhtSptUJ
K3LT6qrmgfkif4md4P+102/BTej6VNuvZSwJRXo6IsriFxVFzoOZznBMA1qY2+e0
4ZdnGlkaXegi7tNX3CYER0GOW35rv5cRWfV1QHBLZl4ZvlMTMb4nyTpv9HLRqXOZ
ugMcOhqPPtJvdGJaj6MaJtx77X1MpHza4gMr6indyf1cuSKszPAdqqdpW5+1uHlr
B+1lNY5SRwpfRU0ADCzcsMUK5UeFzaJzDrva7RiSEkgbIy/FokUsZc99mswouVIP
oBKWzXK1JwxkRa8vVFhwZ6MQgULsEwyTFjxAd7q+CnKBLs3QnT+fI4A2cBpqYslM
3n6jEMQFtAj1BPu4stS8hhvGkkigbnOa08Lc2luioa8TunEJ3qKRkZnzM3KYR8OF
sycK7UsizNNoeBSjA48aR9OQ24+TjGD7NZZN7XK8Ev+C5xEZyAFe8AJ1vgoSpSoo
t4Me42Zw09RkS+GDJhbSana5Sdf+u9ofvSAGKEb8eeB8UwgZX/aHaYNRFK5EYJ07
yNd9qziCc4oqeWVSD2x0dHO37jHPE0qk+dtrCz78g56z0ecocNxYoU1ZsORfmPKZ
GWGKwblJhAd8UMah0kRsjDJ+z/RSxr9nzHMKuXyTh//MAaTwuCjJce4BIz4BeTNk
Z6RQ74Y6JWcV0ZZXk+baTRbQcrWH8i9i1Ry9ZBFYuLciH2iaPhUx4IJFFQkyFf+z
3Z8OnWopSzJ+HO2HYQpPBVdQMZy0WpOpOgZBtsCuWM+BVJjckhSiht92edDsGLIV
GcHueRPcHuPtgxEGVdMWLK4WsxziNLtAfeyofVJzi2bXh90TciFlXkzE8zSJUCPV
i5S+XYM2VUffl7lqzRmqIVwc09y1citBZCzOtB+MI7Rp7GO7HzcPFAaekZzuegTa
whQI3/qB5yH2GCe4zZt4OtwnTJ8EMyhmZMtQi/6bZddRiSUYbyvjhTgtW3B9Bj0i
8W21YZEosrtpPKxkTbYx2plfU5FuCNjR3X5mlNZKNYYrU8wP9R0q3povFxNrx4nO
r6PwK+Q6XjXURQ6u0rCq0+nVhJQYXm3WqSDRrDol5f1bSyEWPwKyKXGbzFoZwr0m
Q59ZxGtPFvDz3urFZbJwWdiwzTmzFGZfwXlcDJ+ti7PZ08ipuyAQ2XO7sTm0ZiGX
66mwqZgHKaEczAZcAzU+0pdD7lUU65CRFRAA7QJws5C8DtnTudrd8We3/9ey3KLE
RngH1tfPjC6nsw7ySIHu7S+YXmYKmN7RucAwfwIJ7Hou9KypRY7bCeZfeE4JwSFV
DaRs4Qbse0Zr9cx+pb3IoNcWx75aL+Up7G/osmicciuqHWoWK9r+aaEr/joebSfH
B+JNRxE9nGdY0OzzOfUe6aK9G2ENKW1qOvsIY/j2eatr44/pI+FmcqpR9h/KVQjo
umiu6s6rjwj/khpydYq7ZjTmzGkSFQEENhJWkt6b0qqnP4ZVDp+u1rquQyY9ooLN
QwcLALU4xlp4hLWafh/HTgx+dveIky/y7YFsLvk+fEELVFAi4FEt1smAvjWcAgHQ
z2/fXIkhOSn/yA6nkrdEnjxcsCvQwmod9Fb3aFnrh9A3tTgUB6yNdo4ezshL3ONu
8IxzEvYk3s5pdiVK3g3Nn3LV18uIqW06PSC1OBX2qSs6K34iof9L63Vq+so+JQ8F
LS8VVj2f6/OYR2Fy0ZGFqUagT8sJ7bq0aj6x6ATn1/1Psaq/UbsptpgnfmgLRR3u
Y5V4NKs1IFbndCKqTJlaZgwHUO1nXik8bjdRe5ufhh0tpwPsHTireaWliIGOJ48G
wpo5hpklsZnrX79LVQznES2jgIbD+4vfvkR4OQgilVYP8LkX5XIDWpJyprZJoqEM
dU9pali5cJ+lpPbaM2PZ2c0RtqwK8/TmlZh7wwzaipxPHdgLgeJaD/7EEIfoueHT
NiTMgo56FkU9DVytRB6dtJchu898uJT0x1OlLS95VYYVdxvLCCGAtX3DHRE8OiqT
BCFf+56yUCZhHUS7pDwwDvhKBbsUvFzpcnSmMRxL3uNsGALHpZlPIzwm9iXqTXQT
7Y6s+g/569/qdYoaM+C4uWUeutrFMeU0ejs21zDiOGW2C4hfUTT+wlnWlZ4BPfD0
YhIJawNjn+axmbztsRJwV+YJBS4ga6KOCxkDNnhJo9WMjSoEhPdciZYuV5TLbaHs
E5QGzcg8KtG6cdKNESwkMRrv2WBS/4k3hkpp3S8XWQW1dR7Tt9CFUoSCEulxCLY/
mKvEYiRDkg+CPQMYAyV/S3kejQTH87n0vZSjSaOTOmBdmHEraMZGtm9Pz4NbogYS
kBjXoINTTNyvaVhTw+bXd3F4GPbWByLU3gGIy95/lu+mWt6JVq1WsqvivbsRgcHZ
cuaLEaCOA89MkjwNmSH6STbHt3+GfbQEpcuC8X6xCaE8eNYqbJ+fmdGrYyXiNGoA
OBKmBfKx0Y+/u3IlT7MrZH6/bPhlnTYxHRNdzV/MuA64PnxNlCrUSdKd6DOednx6
eZ9yFEQnd/jEaefa8SBR66zM0XNHAncP3VyYA28EvmCWTeDNsVQsas+Vhxz+KgUX
OJNEvWjD4fVWtzdp1s7pazddGybBrgCsPMHZpmKUYq/6LQnVDCoPsgrzKHuNoqwC
JANnnjvBhNjQSmbhOA2UuOwzRjIxqB4LS7o3NADvzykjxH7fpdooIuO+R8xkqOom
bPdGM6GeU6FdHgZNGtbjqCL/wPmoY6+1v0a9beC8Rre+46XpUQ4r/z5wzOEmbuOe
bD5vXSAoVs+90qa2QZY4P3uim64T9rSflDFfQsfwMqHwyw1HJDyB1Ev3l8WTcF+/
L7A5P91oSyl23hJA0Wx9UpmSXCoKsYHCMWVJd6S7HWMVYU7oKG7/kSyczHbaWhaD
nXg3jfXVy+oOY0k8dI3nfLPML4jVJwNX3gFD/GEDkNK1fChpdo3RQK1Gk9C7ZZcX
I+DLpS+hs711GdCZigChPSJCYpLP32NQ8qgOB2EPi2WRPNQmgXsR9jT0EwH0xpfs
3h8rztdA3o4SfDsanLHx1J6VSemXZKglbjvGnInWoNikO3qglRrxDyRV/ex+DcXx
VGLJ4h7DaLXRyIGSmjrbvLknhsa/TmCUY8yM9q9xaTPAyuz/KNo5h0DcXrzrrU/p
MmwLsj265x00nfvY0glT4nJJYH+XOjLMSIzcOFnR617UXkCKSQOa+RDi1RixbpNq
M/4C3qWuJt/eWfE2jlrQqjC9+NRZf51HR9+VrxYBUn2elSbLaLJDrn6Oey5ZZS6w
CdcSbzoyak45AFVkldzYis07viy4AQrgbBrmS/a2NAdcnHrRzgdBhJVm8jSkuQh8
w8mMtIu4/UMKHWDf7IEMoeULsi3qUi7tePABkezXnvq4RhBOpsP+Y/c51i/WvrpD
L476Tk3Nxj2Cbeh0GFqSdbTKuXEvXgqXy2VA6ELfCUdcBYH2T1k2vA0fAOyALcaj
9KANWyw8jyMX+Rxya2dy7zgQj+0JQsWx3embKqrRC5U36GcnxT/WdTuI+0wRuk6O
/T238v2P9NhXI6Cq3x9+aB7beWdnPbmiy5ofr2AV13i3aWT8/CQrqXbezY4zvsB9
G6rokbvKiDz5WX/tB1kdQcZlV9xKwAwoM5OVDCoBeygk1fulpY399NJGkYV/60kO
TAp6k7+2M4XdnUj4aM1G/9AdcHSm3e0jBvPN9XcN+qAXWZLXcLkF4rQx4NAZ37mu
2Wt3Q8txvcejfYFFFjVTC9g68iI+U3r1vFajiqnD+xcoqit1BIIn9G9mS1RFSGEl
4/TB7dn/C/4qtujLvbEuIKUEJILAQ9WFVEXBlc/31Blhz2ozrUn6cvgKDXWyZl7G
ZatYYiNYZQl0jRhAQWIWFmEJIDVMtKWes4L+my021e250vTwuMUCklshbUPOSO0B
cyscRX0njBJLXoq8mWcOhD4zrKRnEtapLOq067sKJblOdfEYhIGT4GyamlWxVLz+
+4zR8VtE9RZjG0GfGBSMQNbai3ExxMg/igBoOBRyLIsbyiRrbb4pi4+QlFRxL8TE
YdWBtrE7AtcIVA7jIsimEx5J8W97dVJURZWIF9BK7ngDSxeeOp4PAYoaeP8L0waU
W62d5Q0CTSgKHVQaDZAZ5ACsQXxkXL4UB6QyLhxqE22/I4+XFZjvIkVBZOGpRKdb
9+hpjA+iSkJ2giRuw6owfzWaw2Y+VScUhPPawXUY+e31IWsl4sYEHkzdtYrdcR6P
BndaEsPraYc/g3hrIJwYCy6iEMauRB99NF5KLB+FpPqbXgaMHbiiGK5VfTA2KyII
p8E4C9oYmgL9cGB8eoURE7KLMFyhApohfjtuO0LgRnHiX8FFnodfInD5y0UTGAUJ
yXyPW0jK0XfIxxGwO17hKVT7lYFrReOMbGyxbgsJCWC9Js0tzb8Rwewe2xFu5RD+
dg4B9HCp3+VOe3O+nLKwhBxp6EuQ6duwjFT17g1qjedCOxw5EqrDQonlI5HJmTNb
uGSz9zZHND6rxjeMflE6tbFIx1f3QCNaJRedFZmHhQkg9uan8XmyKNaTgiDMLrp8
bAQwqh1A/Cd95+RSPjrgdGfvFij2nN4hhRa77Tw9frEL7EjFM2lF9llyNq8QvRCa
YqfQxjyquAVfr33StTL+SZfTI3d9E9/QUYAGYMo8fus9ckQ8iNP+MiasSSCe7zjm
FFkioPbGpMtn1IbpqRibWgQ4ukrlPUSIYLTpfl7atIZPg/2WYRc1U6/VZI2jhvYC
3qhHVtPAcDCYXUJ3PtdLbxykO0u62SVdxz+PSHZCDmlX0eIAYXkbaBuIPewi3A1E
s6bYj22nkWt/xRIxS7FkbrhX5EynBDCgsLJLT2SiBn0m3itSh9EOpDq/faa+hfDV
B4qORwB2132cQFNS55ZXIj0G0D4AvAjPFAfuKN2ZFhKDpPo/ihN6h5buMkLRMbqw
DCYH5Fcz8Z6CDhiE+Bnu7f1lmV1Y1hvcAquw4WTXRJ3Xr2vFbH6qSXW2gdbF4iSV
m9clD7U1sesymiYvJQIpz7w/GhooPSjcDcPI2Lics614GsxskCD3xXDAFvAYPMAk
S0KdviHdSPQRs/RL46Nm3GKKX6sYrgKhXJjprgUvLKWSjC2/7b8bnhFMGoP5O0c/
bJovRAOErIofY/HZhaedaSb6DWkea+eEWudbOIMPU4cvZ4cPul3TctUvjm4rrKhS
ycYKPYOrz394Jw1DrhMvJJkITi7h209rqwcC8VblNXCP5+I9TdfU5k7DttarPLsQ
kZqehQEfVFQm19Zw2IBmLKTa7kYJVkOVMk2ch5ctKsmXL3wIBbfCYYLAq5wqMoNF
Gj0SImns2ubAPlCZ7MUJAV2vadfLu9RFJIccTml2/daNJOlXuMq20ZDHYtpSRRjP
3x/JaBo5eLvVgvHD10piiX7N0zgiLenhPYSZInYP1QMk9uOuGzwCBXEjiRG9F2mE
VuDXwRbllZx06XOkThUwFbNVD448vzND6JRaRM6okBBVpL6RMMT7yBMZKq+edgGT
kP40f60JJxMZo05IANHntsVabwiYD3OBvKGR0lgeGM2Y0mdVJtwqGeqMTYr8b1O0
3bw7K2TcMQj425MrfMJ+tvCf38BzxihHCIGLKRDwhPygDQgUhfhX9Ozf83XgYSV9
NaOxfNTAK6SF9H+AkYKsICWg2It4qGLH1LSbJiNFg488E5N6yBAyp5RHBAj4FETY
Cvjy9I7CunLHcnsVzZqDETlbyfSstJ9UnHooadZo726LyJznuHvxDZOpTtqZ3fjJ
Wgaj/vAHdUy3XrMxXKhSPxrAwFXN9zSoW6E804v5DKnPbU68eay7SAOMzo0SuyG7
i7J0mOVLWX1fJC0oiHrCC5yC+xgvSO+SrufFFVUlXNv9CIoePB+K/O1iY1GOh2eC
dokSiaW6awCDNsDz7B0bPKW8YEtN37TYeP6g5W8IQjIkeyS9G/vsIWFSrtmV9tz5
/vDzLCbVCUVy8i9rYSeVpB1KP0fEbHt4Y1oEVU+3ZpgJogvWy9koHUdE+cKFxkdO
EgxBaZBfgVSMvPKnVFWhCBiJMQazJKFIC+7vFxP0DE5Ud9Mkn1Kin/vP5q4HV4jV
VyQDO6fU21r1ffUAe/EquyVica0kApNixcPOlrOkj6Y9BLwYNkASeG/V913QVDvW
cFZN1atASt5PFpNNBeVoICzUoPrykbxfbS/epHGgTrOTSQJ8fyvCt1HDO8yevbfz
l46g1AUBjTwcjbMatkPgS6o5Uwbolm1oCksUKkp5I/9jvSWb/nulzlbFlN8xwOzN
jInsuop/Ho43f8IPv3spYf+Rf9W4MVS7fhzbUsS6QH/pB9XRE8lZcEpXU4kfz2Yl
u2M9HS/AzMiehxVNr8ThOsBlH4YhvbnToNW9unwiIu1G4cHlJJrP9BjtANJf41HY
QR9eUT54I0RniQLYQeYAT4HZ+hOigEe+6WQxbPFLxKbDTuCG3cvIhM/ZRDeheh5V
LJ4lD5lQ9ewetz81n09BbaLPIZtlQXVbeh9KnKqSsurSmFIiRlHXK/InpIkY6iZg
U27xnQr7B74ImySXnUcBTMwK+dqAZ2FRslDunz6gk979MMbqsJnqaJtpSfCW6xHd
cs2VettKqZv0R73i0ZUI6BqAwj7BgtDj4pYx23wtHqzEryqMINW2gKGdV4vl+Ohr
u2BhfqvyQ2xSgwTs1Ih4MWf9DktmSfoQ3U1+leSmu4R7HFg93pWS6EHn3F+uYaRH
jDX2N4wrsTat1nApY1V2J+BEK7vRW9u2UtE6I59/Fpq5Jyp+vv+BYJVuyxMnLX+C
VuJEAbYGN+hW1B6Bc4lVZUQY8dqTo+1HQYB4/w2z03+4bSI9UxgxuJf2a7/Bw86Q
KkyAOcLzmTsQCnNEk2H3vJ93BoISgMsHjXXuCgaGW/GX0NGJ5JowIZfal5FicAxp
5G8XQfZvJwbDNoLvOOnPykdMcdHSzGQ9IRPerzRFL6IkF6ww72olUnQmv6foHH6b
qIGeKg4HEsJ5qq8ciMkzsVi6XtgBpvLlQMJ+MbRVIVrB0wC/o87xGr3hjrjeRHzs
wyqGh46nwCjba5eY2m8hAxHaCutvNi+Uoly3lP+zcJd1B2sPw+MiSWcdnK7BTgwp
afmWcBnPJzL1Mbrb4iw9kID4aHsT+su+Qthy1LTftAEemcfIjqYnuQXJxsDPV2Po
SL+MoF8mCEn9s7DIUZ8CBAB80rN2ywIB69lKIw2edLJuebnn1gFi8M2I43qoGy7K
txSu2W3cEyhxxBhBbsBNlxYxtyY4aNGNQv11rcrhkKnFTqxBYbvRzK3wuRCHOFd7
ogfS6bLqo7nrPvCn1U54HQH+9SlSEgYWZJI9diZzh+jJbcbvQou+8FwdSRqzzF1g
SIvZxYrQC9lQhVLQECoKSCyrc3PmpTDEPzreioweFsFzN/PDoTe8luaE/x/+6/7I
IUp8DNO7efLM4jWfjqjsbYr0wQBZnZ7OhW3K+uFQhogFEUFafqLiOgWbZ3JmdRIG
Rl//p96ppeo62tqxSIh9wEf/Wzq3UuXCjQCeIbOkhU9OuIvV12gjcu8GO7CRfQHv
q9YRUJ8uvP+EVrTXqlyBrbia62U71TniT7meFy3uAkE0lJ+gIL1xCzpNxQq/Rsiq
C3j/XxEDiNsgCqBIH+8E5Q1fk62NjDFd2MqTC2pwWyiWdCPi5+3VqoDQBZmkQ93T
eZ/akgS6xEjLirQy7lVMPpzEUJTuqzJ9fIaOnCqocQyk+fMC6Gns4UbMcVTah8DD
O1JkrDMNRfERYaqdStiqZ0wMtNhoFdCfWH2C58gdNBgN6+DLrHESRaajxCj5wltr
JCju1uiXzRpct35UJ3X5ffIOALn/5duHjgfbTIOHUFKfRo4X9ph0wKCLTO/wJy7C
P1tg/FtfC32EW6vq3sAv901OAUyEaa7IGZR5mYnWaMJd5wXyOy1Xa8uXNnMTkoF2
U2xrvhU/zd9CPswAXlcJeYga5PC95YdZwqBbuckbp+j6DWZ+tQPK3UQ6crp/M4w8
y4xijU49cOx0FGqyWAEJ0CPLiTJOuUia0rw7pTZRX1/RQqfWanMskymtdmQ3eO2M
gh1ujiAdvIsfOYIachpz8uYWBPnuB/fsj//uwO3mA94InZ2whklpjFwfufrIYsVj
8nR6RFQRQhpBpoKG4F2iQSAB1iKd29VBFmTFN4VSESpbIorx82JBgCv6JyJqzRuW
+RbvkLT1FdkfmfCGXyFxweQhfa5oNjKnDDF/pADHAMlBsqA4YgwGB/ttSQsJ0FLW
CZj26yeUrECkdnGZBfCX1dxu6zIBplH+nNvKIUdq5F0XeiJ2Jql5XwR2Ghbn0iS4
qhXKEPXW4gMIwBzs8BMwskkK+RLy2tCMAh/f4s/SEEXcqNzKYia4ktsp191IS+bU
dqYopQbeT8dI/ybVn26hNk54xXF2Rt6Ads8l6a/9xitr324QUsw6L26I63YI5bRt
hIgWgmQeKvkOvxotx/O6QiZRu1+i0B1gRPqeyNwoWvfnOf3Rl/fnPIFBAHNy6L6W
fIvcOU7gF0rfM7SNmRRKdpJJqsxErb6zXeULtBn9gn6dzhIfw23XJy28WRYjq3NA
ZX6BJPDcNhg/GX2GXMyqwcpPYZNMAOkHjUSSRdFdnKjl2NMwMfaK8rxj9L2aGDY4
noc9G7H2xkRVKEY33Owq13+aly94IaLCRLySqKBIs6V10XDVx7ajPCm9578HS0/W
ksPp3EEzZBOdGJXzWHGpUoSqjwWi7bhiI762IY0Wo8GXj6lwa6x++e3wDj+PkB9p
Vs0LjG+xcGQNm9T6p+EOW72oyOQ99tiOmxEncgmqGABTzBJoRN/zXznbdsaUd03d
zaToaBD+TjEpc42XFNHag+TCM9mlPWDCJ4tN91OILFwTaMX6v8E3mclPaOm3s2/Y
SxlnZFlu/oTZlH6XZkUYTBExK2cRZ47C20V6tAiNtxn4p++veoURR4+bl7fkHIr0
sGA5ZDG06IQIDr3HamizVNYk3PrpzUGydxxY/m0C8TmFZ6K4mE3gQswwy5ch7Ngq
sTfpU0mLykpLFqHmZTug36roF49ZUnaWazt+Jb1fETNm+oU5IKsyJKY7veYNpX8s
hVY4Djl8uUgHypmLr6/27c7o7m476jfYmfTwxWLf+K0XwtW5pWhIvEb+ALLH6cXu
ugg2M6vLWcYOOgxKC1bRsyJwi+TkhTFaVMOjV/O0MZSVqPeKbUmjCbuLqGMmuOKn
N91YQ+4Jwyy7nyhVuCjGKgRDU0Hbw084Pdc/pYkx4O1Kk0Xn4neZVv6Ke1fhX/25
pCU8BsH+xnCGMiTcavAnZsH4J/1N/a4zjiFnBxEwdP1BhGQbeQTyESgtrllXbTT9
M5DU+Gg/elDm5UyCBQOCLCNehVjs237Z5Xn2Ls8AU5a1qDvDxz6xoP0iCfwOhLqm
A1MPA3CAz1UuvKY5BzKFsKvldGgBJe6onFCZuRVwQF6Bhu7FqYxRi3G4SJLwZjif
wPZ5Y4BlC1CpBvQZn2GPFPSbDW7h2YZAkF/k1yq0hOOcrKserf8rvDEHSJ9y4nqp
O/kAIffquKCL5NKSRMdSEMIaFZC99kLpsLXO2GHpTy9zOIm7OLrx0hWIESktZ1NF
1pfRWw0fJWk/ivoGY8WqXLQUlBbGlVk7u5lyhCy3g6KYVIYjaYSdULi12bkZ6+Ib
rrj7PHbD7LK2enJjVA9m8NYKLrIVOuv+aEhEsNf3f7/q+4w+bjSfGMv90e9RM7l6
H3wpRrlMoitLFLhwudM+Z73T1Dft896Zwh22LJ8Qrb3G46sbPQw0p2GfprEzvF+t
WomAVJYLSv1OZ1R3h+C0v93PHWu0M+C7ux+3bVXfewVpVCitSg6VoA4VYqVgzLC2
3pnAk8eJAIl8WTPYm5AJN8NMhDWMQI+VaiEi8liph68KcFs3903jfcDxnV/r1jxt
+zPk4QJV4HRJaNxUiX7eefS23QXHo5ZwaI0cIhleDuPPxm0dR64A6SXBiiKZsAI2
ckMZ/drYSSx+ZupR5FjdQknvqTJA/pJdpm4q0AaFKbDyAGXObhXsCqwYKh/uDRIH
uYYtUpxusD+7ooaOVXvIJEWiQH8auHRQcAMDzg6JsCgMhXtIzt+9KU+/l7rm37x+
UJ74tvBdRIJ9Qu3HPsDM7ItpCVRtaEmYhPotoRaMjEZfjcSYC+Ohw2kjAQiOhZX7
TCcXeuuDIO3+93xc5bplgZsJZh1vSaY1g1eWL2wvubocRxxkZQlpTTh/cdbbgI/x
dZuBS355uXWZWUQjEdFTRk/67jHS2hTRR+SphLmXey3xyGVZuKagQxZm9Z0eJPfx
t/eTrH1f8yYCEWkjPS4rvoU8X4a0cCLJHpMh9UR7jG+Sr4t1IQ2ARdbixhk+WEGt
wQRWR8sGntq4Rp+VOSrFgTY3To0QflTl4P3D/TMnnrejZIpsGO0HXh2QwOgdKq3v
bEipS6cWsfTWdqiDhXR7PxrHOQZ6B9jeN8toQnNPNleDXrMaCyczPEZXeXrHIy1m
aQjOR8SoIm+DJw4vefZQJ0mkcO7dyY5JGPnzJ51pjQ/IsxJZNeuagLd5IK7ChKBv
Nli86d2LfHj1jxhA00gBQ7G3ldPTpXGZ9bYNjOXHXbPYDiXp5czLN6xxuXdjJXas
KQ4dmIPGZL1tkIxgLMko3/QpeZgnxzTjxi4P8P5AmZj2vffnSnbaFPGpY2DrXN8M
On1SURBVbaD9J9rKhKsvubSng5Xtthvob9xKn0a7ehhuxxqAx/GRk5MeLrlD7/fK
aNdWnJUVQRMovP6qR+NrXLKmsdDVKgdygmREFqqThi7DoFz2rtC5bNoCnVk8gQCo
Uo2TxXdLHxMvZfENihbzGo8ePTURdrAH2ym2K9VOs4KLQmFs4nR2sNVePo91xprB
JKuOeT63bP05bkwj17JSxW0LpHoYI1Peg1PVf73A6dEUhRcSQimf9qBU19B8Zbgp
xYS4CTQELAUlRM54AosCcOy6uRaj8kNpn34okwt+ThjZkTcxvbKq0veFAmWMMLi5
YS8h8WdBRKDzPflYdqlv5zNAoJKz6RIho+1LHFQRJTMDOlir+cRPW74pcOdICols
sFJlkH3sNxNABqj1CwOAqDzR3SBze3GMOUf8pSLmpyfpZQksn20s8ib3TJfDcWpn
6teKCgzemcPnUAGcDGP8Pq2+hne3Y/qlETyfrUFK0ARGtjP6PlwQzTC1DIHRibqC
N51lZ01Jgqx+ZydTvlVhJL3XYVrmDX/M0qQn4HE9FAkVrqFmO86SzFdD9S764ef1
oxsh6xVxM64WA1RS3WWp20h2YPkDSki59pHRfyOB2ujDiMOvfrAPJowBt1vTIVFk
dpLimotnzSOgYOBPwD7+imavpug5METrVxvwGm2gAoawpr35D5f8e/Zl0RNuup9i
8RZsK5sl74H2R86a6W0L7wcc0PDYh9D4sBOxnxauV3l4WOa3l9txL8hcXBSBXxCX
6ltnJ2hSlhBjkusKET9cIXa4d4O6r70Q7SA8OeFQt8EsoFA52cL0h5JbbElstssQ
TbqwqCRtGCYnDT1Jm2ibPwgItHLSxOo3EgRtfSkFVbODwgcjRwrAPkjGk96QdOxW
O3zBGXf6Po88sILuWyg7xLyUuVMwwhYE318P4ia2kMz/R//Dl7aLHBxSpVQdl+Gl
HMVf3Nfk9WBj5Ztmo9OKculBkugJ7/jfvWxOoTXSPEupmhJnszzxOHNv4nVsxufk
kpHv1LjlaSF7pWUIOzNB1ktyvlx/Qy+cykRI4PslCyL3BQ0LOVeDKr+APRhzUreU
dw2dxR3uVpTXuXsIdL2rlU3Wc7C1lu52sl4VznciXjzwlcbJb2qxM4XMM7pQN159
KyrU+9Ak8JVuUrojBrolR3YREl5jQRks1XI56BSAk0ZVvGDAnhhPV2C1TwP36Vdq
LVGZqGY0FEJULBF39dW2cyoDWJHAhYELi2gaOjsywQVW+u1UoBlWhnDhDz2D8rq8
mxiTOLYWkpce+OGWdfgsiNJ925CTGTwByLw2KfBcu9NowwFiojBEz1j89tfixlz/
1iCviItqdH2pI+x9wMjjWG/Zag86d8Bt0fMW3Am3A7XqvD6pemKoI5DgNAAW3Fys
vxYf6INIwlNOviSglAAQTMlcmlBtqqm/aZDsGLnO9Fktx9MM7I4++1EQ8+ecIQXJ
XN8X7F7lSgw5t9MdkPG/Qxq6REYxhJzpbWHFUyKc1Coh9oy0N2pVZg2tOgdbiOJ/
83614a/AQvAhWfGbm77gr37CeGPlSYtt1Kk6GumMQih1q44mvzaE5MBN1YMWjs/1
5ejIYyGe/jV7usqRE1oQ2ZqO9S70bH4dX6bGO+PoHPM+0K/rR5gGJUIhpN39BXRL
BSvs1RgQWXRJ+jzn4y9IWN84GCUZNfgyJ45jFuL6pqqgSdJz9FoKXC4LCFb99IeG
h6dh3Si4RCx0l+ZDeNzOtwqbXPUdF8Y5tB1nKtPUuCQ0NxawCZYvaPcGBer7H9QU
DEpYkzQvhKUrGrIh4ppE0meLgJixus8F2wpYGtK7bflpt3cxffD5HdsnKjZg84xe
eavpoPaCsnAIVnk4As4hpKKH2DHsi6FgDl1z6T07CQ3YP5gPDoOjZGJGa7K0yJZe
FuzBEXbyDiwbUoVlsOSwMw1QgiPLnx/9iXiRtNQOEhJCzDGY3zCsZZsZ7R7NNWm5
gavIPP05ahbbeqabbpK1ty6nKaixJLa2Q+bV6yX+0sVXHcqiaVpTmBKye7A8318l
Ar3arHctclE1lx5vb3cPqcMxrpr+APWk0icj6dtdjEqnxGQ6+3FcKovo3mebzEWu
dhkJyyd9BNiw1/9vtTDK4/r8AwP19IK+v9NU0O5Q1rXo99v7v7VOMnMudDeANdhc
gcLapHL+FnBpXaoGN988tYQ3LAMxiD/hijDzSlH92LMJ75n52zHcOyZiUe+BNcse
NR2qK+90l6PXEwoR8osB44alH8dpEnhfdgm7EIYDY7znyF53GhevtH3b11cAT0gO
k2y1J8WWdoS2sYnWaNihsVsl2MtX64O1wVVvgKVDxqMKcfRbJtoVZvaJiADdm1rC
Z9QQ7FGJdXgraOE2epKbvm9w+a4IF8VW82HtQyVDdaBpKcZR3LLW83VdlAIZRAV2
tNN+o1hVzpIFuPxoaNcAJhzhU+zf8tK5AHAt76ObwXm6WOuwRbhidskUUoxLkQ1p
QXq3802h6iDn9yJ8toIrPJo3duOF09KO6gGJi+rgtR+KI06GRU4jxW19OQvXfwBa
TWIBn1tqISzZaHfZn2XOjSs0JbpE7K+XS95iOndT/Q99GCbZvLTjOX8hh4sUOGVT
WQ4/TzapICLJZbCd/OlO1jwiFdE+6DpymzU49bx1n4zW8AfOBCJJhAmDnUv/uuAX
kuRVCP+cnTvAsqRYERb4K9QU/ObIrQyWtG12I1bKxKj8AR4s3Z0hstLWAuH2iCya
q8SKYrcy0pyRPInLQSmEIvO5JZwpBTW6Cr0pX2rwP/uI2UW8lhB0+gyESC1Jl414
Q4d+98P+NGhR4szBvaZDOalYFIdaLXnmq+HEh1UQKW7VRa2G7Pv79Tamj8pGzC4U
1WLtxipShJeM89IeJLhjiaZ0EijwGkTSajuyBbigJ8TnZ9w1kW0rSvr6l08y+cHX
0vQVeKpZY4oDH0nIHe6NfR2gH/KnMOKoCemoianRfN23get7PK9I2yUI7EmFa/I3
2X8wUyaSLYrCfhZjZyy6pskU1nRTT72HxlI48JlxU1U51lo6QKrc3zUgtetA3qtg
7Jw+K+whfsKKg9T3cPjjBawoKvKUhG/F7U26xd42+pRsvjdSVgmGEpL2vOl3XZIC
MpCD+qDITd180DVS+u9JpoJ28Cv2daWYoPbBKs0jQepGXGDKIlYjWh5+b+QKWppA
F6s/Vn8IUWl6y0KtSfkWS/pisV3mExjvW6EbgkMBuD744vQ9ztSi3UC1g0uVeWn9
DTWPoJPTkIcbkaUOfksaOTFiPCPvZO6qZuvfXIhlpQ3IicACYI9jPOSUQbF0imgS
sbeC9md1ML6dVZ/T30JcV+98U7AzJabL9+60rcVj66qN9lh1xp55YeGsr19Fq/Qh
x9ZGq5dFYygegGIG7ERTKScVJKfd76hMRuu2XUllwG/iXMbrKUi3dHDpq7asZNh/
kTMI0HewWYn6e3Ygg6p7rSXXaMwhiFXJP2bDGcmYByviF60O3enhN4EuUDRDbYUf
syK1bIxJ12J7RI5RuM7jgLGnelouWBgFQ9MG4mzCsZ30MnilEp71alvl8318w+kz
LZ33hmS0pOyMpT0pehTk72bQ3z8fLfQCFlWH+6gsdw43hB14mspNc9Nv9VF1fD+f
nziRZEYbJ3R239LvTrucqyXcyTqwODEU+BIJPdpGpye1PDas20CZXIN+QpwXLIp6
hZJcpxwU8qa0uKy4eUSIKbjXmC3muqnhfBRE44kp22cKTo5MQiwpQ+gGTSqI2AZF
WrxynGdrorWid8R6rTVyRtDkva3GLK0qT5AJLCkQ9pD1NB5AIWfC0xMcNQzSTRk8
FongvNKwO2n+oj4J1Bx/WVSMff4I6bpQayC4heVtgjMOjcgaEkIaC9uinkbbsL3s
QtSkxgGSLXDE+sHO3Red1P0rth00bBs6OYBZuxlSQL/vN6IElFWIqQIQet9gXXJZ
N3m9qstSkWZ2U0SuqebBq0lr3Y1kEOqYzZ/tZj0ycLnpWgU3Y//wdVJ2vY/bSy72
BXDS9FtNMLT5Hu511n3Lvahw90Myoajbz9ETUIzj5R6XtyKW4+TiMBRZmH8bC9gD
UE9G82K79Canyasb3Y//VZOiPDFsnsa0ZFLMJRvzjzNuJQUiibNaNYwVf8tEGF04
3KZd3Or3kdMroSnA6uEHC/WfcYamj3+43yxaUwTzhCW2wpxOPIqpIvyzteXXSNI2
vNBT7rvw7/K6sMS2LFgUrmTOQeCRTjwhBLjfsS88qSqOM08Q8K7a2/mDljazKkck
3w3f1ikMoGEpFIDU9Kt7h4dFMukztHZoLupTFk0zU1w37I89w2zADIhOJbmfpoRy
si2bk6Cke5aWUI7AX1CW6A4nzx+QsZu4fqLIv/QcxwR+dvmF27ZpvAlXyP+hEyep
VgtdIqW57vwkHqzPTU8SrZBeF5tc/SKd/AxpIDD/FQ68jPcrTQKEq/TCo84xkyxu
Nfdv/wAqw8N9NT21CC9EuRfT6EZ4Fi+O2j+giOBBiMSa0ZZ0Q8zftu5pjoZEtTvd
1H9W1OnLuy1ln1+MJyZEbiWqHSkKkwOmp5iqMcpVmM7RC5HJUxApQ3nMuPjdAyb/
oKwQH1eOvHwVAkAMRm7fAhr5Rdd//G+nOQs4t8Z6MCGmWt0Tg2g2AMkuAbVu/6Ps
uL6c/CIeHo6A7XWK3WH1qKCKbwKZeJMKuiuv20n5e11pHJDlMgp8pinQRD6qaRj+
ki9obJIeUGCX5PIDMFjKWcAm+IlWfgNuKhvE48o462Xm1JRmA9CVdgUHaOWpEJ3Y
cmY2IZwyiMVL8+3iIhMWetLvgP3tgHrqv3o6arjeGHot8dhNcvIULFRjkrg7UT9e
OBEY/Ml4yHsSY2F5AAo6Dw2agOfnMWSusjbfamy5BB7v2gryTk5c2Vg9z+X9uXwp
l4cMA6txmga2wwDOVT7IBJgE5yPQ7SYddPJIV+vIosWnuJ8pF9zjCx7kH/zuB+NM
a2oAvDYHdcN7M3CLbcQaL8DksDcLie4HoddNnUd1U0eTIf1+7nVM/1QlniMBAO9P
5FzXt9gkeDiHlO/x//sAGW1J6l+OKwgPpYk97uPMcje5f8h3OhDMC2uqg9FFfx2W
Sjz91TIyUmtFmkQG2hzLf8lkvg08SvLN7BBskde5t9wly9GLxoZlVcvxEBzVy/u7
NyaKrmJH1PLBsthjE6Z9ANJFHTQfXwF/6uMAQXyXTCX8I+J3uZKHiOnHi6nFYMTv
6kQdZycmulyTWTNahO0H6Nnd1Mj0oYZAOkkXvrorp8RJOXA9P6nf9UeyvYXJDJG7
QiNj3w/nPW63bLa+3RASx+E14Huy0Bq+epwNp5yJuJ++S3clv8BOkNKaFAYLYX+j
AehP0qtqsxYDey1ltVjvkuh4xLIudXO2ky011fwfPOxla3k/rQEuycZBgg2IfJQ1
O53udGzzYig/j0iLLpfJAxXlFT0Y9rxF83kihASJwiOMJ4LlZtDvm8tEcEbCyAVf
JAo43mO+UG/kf3eFDeAvT9I94KJ86aVeKm/EtMximfL/NeUnXy0GV3eLt0n7yrII
wnPA2OYm90mSzEZ0eFN9BFTEPlaXFI0FPon4gJFfsQHvvt7YccPF5jFurrCRUz4p
kHoHWOgTfnCscc22T0kI92B+QiLlHzvz4dgMe9LAiy1BwqNQoD6NniVG83MW+u5/
7tRNqVAF2fA8i3pzWGC5XWuHHNmJVMh5875w2gikrl/JVajq68iIf3CV+lE3GaVg
B6VhFud6QitNYCSzB/D1wCI8vfs0cGfZNXgSeUmvSsuU1Bl0wbFnV8PL3ZD+/FNO
84DTS7B4uLXdLqz4IHNg4phxztGfhhX4wkUx/VLEFFrFvwmh4Tk8VQ38ekkn3mN/
wHv5Z5euq7554q4axPAQPlr4xXOuua8uIh/vT49k0XFut2aihA71sbbRIeH7YgN0
rcgEQQzcMzXYNUvWvNceW8uWUxHF23PmtE28kx86wqGQYp8afCz5yHoPgWBkcSlW
JChh7rfNzWwvWa0j24WYd86koWen7SkUEo1G995woNzmjUyzcK+ZHh9Ak1jX0NPY
QlImKDJkSIvivIviE2PHcFSFYmuv64q0E/MnwTyFrO4FaXYRkHxhkg1COEh7v84J
Jcm08ziqx+qYwMbRznpI9J71onVLJdZlZKGxJK8F1OjMmuz0V1V6lrdozXf/VnAh
iwcXJjsSYoHt7QvcKofEBMXzgSB62kWtWiyzBKt0p4jbA5X4unWRkbuxSj3oeU5R
FdCzmPdiNSs2GikU7jXKYGiQLr3cJ9f6fkp2yo6AaFUQK7BCdWve/8xISvvkMLk7
GSWskGnCdn2pKzTLO+qJ6jrMYfxIZNpr++GcYhEELMQPQDNc3IBKAmZYZHLBo4Ug
zYwKUJCpYUBRuFw9f84/Gwh+eNEn1MLEBLadYv5V907i7UWFqncgc4a2tMPxxS4h
hrxsKsJiLZdV4TFOaFfd/D0bT89GopyQn4jsJyFDB95SOOG1kQfVsQJXkGcAmkU6
9Do/l/T4wmKOEUmKDUAC/mDFNWwQk1nsyC81sjrzfbLKuBdGxsXqHK7TU2x+m3Ya
2JpqkQsr2xLlXbe9aaeNe6c7xr9W25NgWNEjtUaS3qO2V7pVAg9kBG2IrbrYdP7B
EmqYtTflX+WM200pZiaZdfTlW6k2eNSPDhQawvj/VXvJOTWkK59/lvfmNXGGyEj9
UDSzXjo5GKVQqxTxvOHdurPv5/fsk+BZm6hy4JRD0ff3OFO+4Yz6YdZ85WyipD6Y
/li8HLkdMHjsCI9v5afcI0fbKuhN1fF1l/Xcs+oT9kFeTENKJFmnhoLwON7b+rl6
D6Tc8mDDJBqIYCUk2Ivfp5EuKYHaoQWHfh1KMfAmvrkc+5ANxzWIsUMHhcUz7aQZ
abIRvMLjT4vnNRLZmUcQyTka5ZXCa+KvRu8118QE21ZYpiw6v/ubTE/u4/pwY8R1
yuGTq/DLPKKjMRAt1efYocnP6yfEyv0dJG0HCmc8sjELP0rri4APPUZwPlkHalZ9
ZUIBFno2fbKpSGtE7xGH/IT6MtjrbATdqdsCNV4HIEJC21nHB1M/PEmLUodZYw5y
WI0V4ikYiOXCpHsy0asIM0bg0VIQLHcEAsdhmP4NjPI+Jkkep7Rmy0vFj29lPRxD
4cek8ONFKGMII01UuuVbhF6iErZYZ3UwQLQ+rF3skMEWXWd08xYWdgqXd1utEVf2
PhVNWWjLcKi6xZ5NUto+wp5kWmMQDq78nezy02TPWME4JX9bOjSKrVuD6RVBmKGr
v9ic8YUKg5qc+OnORjwt+QoE1bnVA9ZpFFkOzqEoiLErwX7uR5yTKdPhAiFLfUVZ
4mulD775iBqg4MWNJ09njAbzTnjVfPm32+XY6VYyApWnYDglsCFmukVsRn83NkPG
SLLYFLQK7SzTB8LActseWtUCD24XaLCdby8861GVMfFJr3ngp3fLH4Fsk2IEnL7P
Bw///p6KOrps2OL2pHHm2/3Rm5pCTA1UDqeXALQ1XKCMqDUsHcAqBXth+AM8yu82
9Il8jFwNRWuP42mbb/deGLTuMdUwTg/up/hylG5tnZp1RyDgqMPIw8PcCVz318ok
YZTb+0Aw3HjgUD4B2ZX5ty0h8atAXEgTo6HAVD/hnecOCWxDffnSykLuYC2K22IO
RXKjg7aJ6C4uenZfJ3013xGIP8tZ6ZqNSoDkw9jF6fOGnOQvIybqJ2qNHDkrRLq6
8b+1NVditWKz+k0ljMwx8Y/Wm+TPUb4chs5g1zMK6d3Oi+FqUDpTBc/kgw7Ginl5
bGCzYY+wjHwBnYOWKBnOaTqfM1wLdvNNwuDUCLxSM5Jl/p68qEBEB5di2piSJP7w
phfNY2Q/44GpP0xXiTU2+d2BKeN+4tb0wSYH1P8xkY0ciCq2DfPjJi+l7jO/ahb9
HFptOv+9NggUGtGfhf3VW/nMlQjnrA85IMpIOQkvloG2Yih6/ceDCCCH0w/1zcoS
H6mM6ny/bOrNhl8BC3+2wxTUE3akAJwk80Laj+HQsjXZYp43hXgZeb2UxONNfwK8
YS3Y32Pf/XcWyAfWkbqAmWvC07+Qi1pbS5UURvfLJsytNU1+ByZ0I1p/rGgqzoPj
a/ARIxDDsK4ANJx+kGeVI62K0FoAdV6Ssz/Bj0PkVJ9xGTKOyomiO+kgusDZe3DY
mnteFcolSprnhsBbFef5RI/dSE8VMcDcDNBdTb7Q3QwJABhg9BgW/avXMfl9P1ny
2P6HhvXiKU39ZHlKwHn2kfZYqGN63HDCwFRi/SObfXVbMtiCopEXBvSOY6bs4DNZ
nG3VCq48eDLTXcoGsMz9m97NvGAUuvPFq/jnMKuDfxObA9ytwrw7CMtuhhy6B47C
yzG4xLTs4eXuAoUapwtlmHtE4U/TLa9jiburOHKuHn7Jgnyo/FdZd5E54NVlYp3G
KUP8J+oKOnM2GU7i5tGaKhsqxjrBNPSvbLV3jBAhYwGhb7dch9P0daabHO2X0lvw
C0EFezn41MHvSfq1/6juQKa7fzzrO2hrTksTOoOl+FxhP64jmAhepef28K3LBJND
R/CYxMKA3FcTwZBxSrEVmTheqHUHGla4vmfWvQYly6rtlH1jwQPQe5uQFT9Glnji
TI3xuCo8evhgYecOHZhCZRo+6Gqj9XBVvhgF7NdoieBF89FC62j7fdMomaBdpeV0
xjGc5uM2aJKbLDVvWG77xCLxiniYfnhj2akWui3NeyUZtUgCUcWCfHIgN7ljKdRW
aMJX5RYvfE6sAQ38z3x+Ue8yzThsIWabZy3cBik3zHKqIMepH2LC9TZy2JqUxZzR
TQ6mbniZYw3555jBiBxG6/f7DdYgZAgqe+cRLovt7CQtGfwVbvHI+HCwDfZvfoxb
QNjvlGpmi6uMmGAhPQfTQiq+NMm3E1cpcGU6yfPjYA5IA8kqeqZtM1OpNRv1hLvs
14MobCmNmMVe/ekVhdtOVIqU06y7LXGoupNjgKNXXmQdi2T7PqS1v7lwahRSUVBb
xOF1vkbZoMjyefPhtG+5Av9sqqiYwm2KRuVU5bDovwg+EiztM0JmCDgYMxi48g92
09xZ5xmVLtfBCp8J1PpTsxuRXAwZvKpEqjvXg2LXQsopMI9z8i2kJL98Mq7/OEy+
jd4bp59ztuAVFMEaR/NKNhJ82UaOFU2OTUQkNUX0dkcsoXryGN6jUf7X6gmd6oJX
2M4ECLVJu9CWOZ5cmmMg5ttfnnd2anIlOhD9t1wL1AARcvwD9aM8I8EZFeLcGqQ3
wf0lIQj114GvLD3JAPmbEozGn3RRBQ9bm4LGf0xIsIpVfckIyrNDoptHF1lm6DLV
e3YomowF7YgcsvAlR5GouLYGg79XeX8dw47zmMuLy7PuDZ8wzOHuWVOMtPUOIf+C
ch148lo8EYjofmL/0lOd+yN0xJPkv+BOEkmVKD+otN8zslQ2yW5k/eQeYSesFcLR
hY4/Yi7Pc9m1/BmJx4KdnZ+lhqPCqTZK9VbOYdu85lVgyrI/BuxnLjHiUifSXtXH
KYv6ZwbpS2WsIdrH58iL4qZOqxwJ0MlO4rIydGEXxukoFAsp1AQmFVB+ihrciyov
Kb0zNqVdwD2pad7T2JrgN/SUclBZJgx2AOB8Aao00td/7D2yPHzGW1Pqo6WRbCBm
iQd4n2yQerP2XHhmJprABrL1dWElxNXWeepUnsJd/8ocZTbfWxR7TAvfPWdZfVJl
XIGW+J+liEP4xoJA0PuNFk9aYqQzBms4X9kMAhvDi9uEIbAfNQHWe+3ixe/Jtb4s
1SLSicOPCqXH2xK4uEyDDG1aGYo/+mn+5EGG0W/kkAqWQd7XTGb0B3HPNZLBWLPA
2N39e5LXiKZn9ALDqTOBxviyITc+SAmJ6lskaRztiiCqxR6dtZVEPO0kCHmk7/bt
uWou8LgsYPNquVZw4Fs/RasfdWlcNuuWxBRyo1DB8UuKWs34pwuL69Bzoh9dMwYA
oE8GiMdA6JNdaQRiWAlBG9re/9DQTD/ErnxWNUaLQcmNlKvCz+UQPCZgUvWbFxDS
N1mKLpLLiPKU+en+0x2OTq4r3i2RxTP1Ko5HHAVFTBbaBbnXsb2xJYQbru0vaSeb
PI+rcWXd6LMT72nl447TUne0uttUfGbvz2I1ki5lQyTZ8jnbFUuEkvoYIoC2O5RF
AEB/KzMrGOecyptYEl8DEpwz9GwfwTCVVvwjJg4AsrHPyCcBbhHkmjIwgsYa6wKu
psyRlw/4zhMpR+NxNUO6ZymPYSs3Eitft3wnG+XzX3A8AX5xiWM6aPTiM3FxkU7O
OGjse9k6hBkX8x4A2OBvMuduYd2Ad26CNQW0BtLjIAVcEWQHs14AiHt+dNHpJ85H
oSF31ERL5LBBWzLlaVVwO4Q+m/0+O6qCqbZbRGnMJQGUOZhWzO1eRkrUBvGDBNgu
nycvjfxTs5VbPF2OX/bHNT3b+w20Ml1d3gdkwSq0WF1n4NPICDKRm4SRzQ4LEyi1
83lTgUi9kZMSXBCKgHCEP2vD7Uejecq5t0hzDNBlolYVN/VusufdPjNHah/EjXXC
YaiAn6RBxyYxLbX8Z/5nf/sjCHJ0oWw4VvpORoesFHGvDhJQvcDet1XnqFTXtwYy
SdEKGMniqGqTLwuy3ViXxBIdOS38pB0R4wfodLl8Nw5ye20vHkoSvkp33qjxcY+T
LfQooR+6c9HBDKrO7SACPc7VvXg9XQhLUyMMW5ZoMHm2ixxfI3LKsZ0tYCtZKrVK
OuMQtUf4+9g9vih4lxrcBggmUemogQ+D6oSUjPQW2HOa8qJpHZeoEOfapByuGO7i
Wkn/SeCeB/oDAHpO1r+HWMMCU3WS+BHwVuKoyE0PvWXA1MZmbmM6BdiNlUgBepCl
t0xCUJRo4+YX1r8kx3fu31qd9ogghK2Bpte/SlIf3WFUcYnlIS36HCzej0sYVEkh
rQ/SAwOm/DX6031FghTR1+uSHaVOe0qyYt59o5MGsSeCzXdIuJu6b12Zmc9YCCNb
MN19IyJlcwhmsQV9da+PsY0ZMrgjwS+0cW4/eAPtFMEzocixAIu9olQ7e2c7xK3g
82dW59Zyrvdtgvb3FUVdiYB7uGXlrPfznlr0eMFEyHSStJ48yBMuNaHupfet1zA/
1R9D63CWho7YwNnHex520ORNGAWRtRu+oM/EaGwAPO005/dxcYmib62uNJL/i3Wi
iFVPCEP6HerWC3/u5MgD54RJ7xqIbyq7WCu3L/EVm3oql5jtNDKSskirh4r5riCf
kJ5w5nV26RWm4WGLzhYIYKJWG4l30+9UV3yPnwB1zTBwZywjGs8CFsox39iRAYGM
APnCWmc8Sj0p9qnBPWX3/DzCLxMxQQtUZpXgzS0J8EcQI1Bo+g6lQzOyWBfbEO6P
DsQlZQvb3qcs6JNfC34XyPOXEBlCGwU1AwEIXzIuX8EeHV79YA9PoRTlAl9Au+lg
kne2ySZVMVNxWOiStu2v1qSbkBj6mGwbt3fc/8b776kYRTREfW8rvg4grbYms8fT
Cdio29h+avyQP22MzgDrhPJZF20isQx+PcEBPkXIHGklwIlpNXHUeXJs+GfJlNtQ
sErZbLr6aGyi+78kfD9nou54E4Flt6uPoNLpB81gbouCAucS96F12tGerp/K9bie
0Z3K1CX9pVx4KZMYSaYRQaxRTTkikpp1++oqSdBbQDzuavYaRHXXDjhpZXewRu01
trJGiaVS9fu+emnPyIyDGFZZXYl1tE9xde9S//+1TiDHW0/MYDvcAlt6Sww3Wd1l
6H3gDeZYz2wp33+jS3BI4Vbf3iJWhD6wYgIxJpZ8L2ZuWWe1+L41co6ogKiv3hEh
0axJ7e04IrFgwOmCAANbNg8BpQ6mY+V7l4UH+HCdCl2cTOprumoGyXPf2JGXGGZ6
2OEtIdGNQtD7JNk2xiFlmsBJOs3rBW/V1HrBn/cPYWSumh9EEqVFFMkgYowcNSVX
ZSPzZA7yM+sBejf2Bk+FO2shNXZv/Mec2VcI4AyDwxuOOtL6nAfHlc8oLQf/V2ZI
chPnqs+LylR9B77ADrmsuocloZjqjAyaoOGP9rKgWQO9oIu1nAcpeGLyG4vrus8B
8VpzUNs8FRQlOpvYusurUM0YOzsvKYOI1GCi4PaG65m3uYOJbyyIfdcWmBSRp6qD
rXmwKSfdJSuukasBM9sXZ86FXSVMAN8rTu2pYDDjrQWBb0TCK1n8oIJ1gFFNIP7k
ySm6Gjadc/S2xfdXJiq1GTKRvi/5+GJK6uwFiv8RAFiJCwI0zCujAhFYERfiPZv3
gHQ5sc0CZVW50+g7Hj/xGyMFp8a+v5Sv5DZJzWLqW+s59p2etQuJu03nBj4se/Lg
L4anA6Z0uJ+Xcqfut3dTjkBRi3D3V/hki1l82ZkTrBI+TGQggzBKsVQTCTaJXzNB
xPASJ+OohqG0JVv1j7FkwdKOh6IGuvWJrjNDNfAQSKhAq9nSMBXU10QA2LFlNTyW
toT8faRhS8EtBOV5w2Gqt/RQ9vC2COKvqikrH3eA67kaeFJmrw0YdsXHzpBOOlMr
odRMTYn6l+nm6DTYZVDXg5MV3IIAOKyqDs/Et4VS2uO3X1PVP21nPB871uvlwO93
R3OzGVZTJKykKGvZtcprc9d1Ytf2RnmN2mVjmfBnqnxprN6QseMa0o0PBCWQgvp0
8D0rRCSwKF8b0wApdt3BIyAmlxsvXB7hF9MYH3bImwCISXIIUQk3Q5cppBG65NWk
rjyuDrMbXA+wrejaX4m4xJDaVniEUBl4Mac/3iQabPQxOk2Su1nhhigchd09Jimi
X+n5IG5KYQQeP1yLxUaC35McdpBK3ULmInN7jxNC31Xooh0hxtK6hyx+pw+b1cUY
wcgZtevBn+6UrbNmI9+zYFa17b5OA+ByEDwXlhEC/TLRqFBzGOtHte+GzrpJnmLw
JRs34TSFADmTrbTHV+lVUVUHgWd9kLjs1XT0MSdixWoFF2mgKb2pCtlIjI2SfV0e
dphlMdx0+BkwyVgf+Kq8K98lEAJgbO2HShZOCQBy0AINxaTCQ5JuzF1GGksjIdvj
+N4frByZJV56bJs+C/ACWMyuyhQ65lmbDeHs6Zv2r0sd5H/x1hA2A2z+bxcl1xHR
PpMBiclKQhj1PZOVUi3I+bjbkphfjXGMyYkkHojQSyLmm9+w68LywShXNQxBdgD3
XjuAQHM+hbniI5ZyxNW/O6QRtsz5fwLDcJZt0LsVsYMVYemfkly7053KhS6+KdYD
9U2fS1rBHNABhaB4lBKd0Pjj+3ZccFalpvSTy1g5aLo6fLiOzuvWgTOYcur9BeSq
J7AiQ3ekHJhNA22eQHbH6VDsHFEQpk6Y0rzoI9pPxuXNVWdzx+JN51k2jwgy7Mbt
Nu4Teu4UJKTZvAvFDCybV1t/CP32WcVy6Ppe8UhHd/Pvvsm2/7PIuDdgJP+Ly409
GoQCJLxsq4vxPD9yMH2MR7srPl030b/R4suuXRY+kf58hF5zKHM+MXm0+ZA1bMr5
rMvFvVzb0op3VuyPhNMvnoOWGJ2VI725m4qL7lEzlOgiQmPtaPNvdr9JRJTWHyFt
YAAZr0nQJfHbQCSYCxmfDs3ssC7TQo5W67RQAZGAc3raq5IegBnapfdit2HVrnkJ
6TtvoAd3cnhK7DIiquIC+r/yA62XlxGjyA0YWQOLghr9e3P2sAY6hEcY8KScqXUY
gIGwjifAfsov+Gjh2IA+P3b9wFpfZtoJMpG3baSuzpmMaaZV/A/BneptuKjmYn6n
DLqAnh7BajUjOP1w7PUDU4ThgqXHEQ9NMXk4tiZOcdJj8Y3VeCToa5HMcadWXQKk
Dou1vt1hgHIbooDjDVKddpe4D7HgRzNPZiHw/DYnsAmbhuE0EjattMPeg8twNmC/
7NL8Lc2J6gNRSLNi4JTHbcJ0eAgfVvvspld0K5sriy+VMDVS4c6JkWnJKkEANHAj
yKOLaLgkOz9VLkqMsGyYnEZsvdlT+CpKGf1KOJPQ6xMm3nkc9xdOrsRx4JCeqbfg
10iE9U325moKcD0aXp7XnPybjnwFxLs/ibwc80rCMzQGlIINHn0Rdi8j9TDXT3Px
ix5VVzy/AGDo1tOWiOQpkNRdHqTewIiRhFnvWfQq3vZOyPnZTzOfyDpY3waLbS66
S0n5YAee7+2yJ+cT4xBIRxLLvg9pOr0ZsHbT8h87ZOXO1hgEsRkO0loPQ+zmYkVV
CYeSLnlENjsTs4GwPGhdYQDcnVR5PIFu8gJnjNGljNCvss08ywsRO0O60U3C7u+I
N2s+1r/nLzwwxxCxpc5Zg+7wqkrH5x119292H92cB81pgPVBErzXd9h0iDAhgOhK
G3jbD3NsbkCpOcqB7QdZ6uZErnDC2iODgCyiJry+lxvX3oUAeFAvlEpw4BpDQRfW
Df6v9VoFPfrXFLx8DpdVJhcfrbRBXLUfZFsn2rz+T89wexP3XmXeQ8MwfpFPke5T
zVl4zXLLOopYP/fT9Bsk8NbiYsvIcXnhEAZUSGMzfxML9Hg3g0mCi73xi8jL9S/P
+0EQ4vGUHg/I4ienrB+5pks3VibXxpDYLYT1nj7APGDNeZHVcASvg0xXpSsq7Xqj
u4hP7ZkbKs5JQFIfPWqhUsxmjQr3uVR/WDlu2uEImhpTYq1rRNnzjAwWKhVadDmd
NIAqA+z4O1BYH0hCzHEvUaUg7eeudAX9CQVFe4adOZY0CRG32CtvGLIStW3BgqqK
KP5/Wb5QaslyLWDQgiZfR4pRT2mQfHOpS5DHZOilsM8NJS9yJZ9lEKRoueBO8euC
S9lupwlJ9wZ6RHnG0pSsF0/xmUixLX0DxQNzfBPfjaxJBXhQhNeJzNU93S5wvVoZ
wGAhwBB+b4YgbKE0t7dH6yYn82MOm5NzOVoTSU6IedMRC29SipyKr9nzRGYzf4Xw
8hcc8+cDAJXj0cl97stf0G9seyMzSYg1U9nIrvNRYJE/GfrzR1iwHkNIJbUlegiT
YT6nDPu1LXmEudbsTsgKqEJq7FLhkY1DOwwFOHiRqAUNYLiMJaB+biCYVPqLNpQa
6uGo5Y8AtnC48qIP9Zg4hXQvXmtm40EtPt1HfJTjmbXEyQFOULJIO84/WaVz7wfJ
+wJvI6Q0d0WqSi46pTTKOKekvFZpqp1VluJ/qe6012m8w43anMkBn+fq1ut5OVut
FQoeMVSWEW/pCE40bc+ut5DDHR9G9bjHgI/hb/5m0nxryjOd1zZkqFs/oeVZKcgD
7d/glV0G84M0aVA2eE3HjzgurTtsrVYjCiInaF2OiUDdgUEvjdHNfTD4YfIaRtql
CQ6vJukyuvU/LERIl6jX/OGnwgI6/qAeweAE+6pgSfOeKdXqhKgc3Ibd4pgW/1se
ZB5HvctlVyFfX7rXn8PP+OSrBNYPgqgU0Are/hN2244/0ekDEZ7cdN3hopHKWg+u
w43xpt75G4MzR9KRGGJOB5vAN8llmJU+FxMqS9DgyHwy8HZkjcoXAn9lbzwP808W
0ShzXBy20VLRmP3/la4Gn0t1KCSxlnbNttkombkCr8pAGOsN6vvCF6R14QWg1QTz
Xf2jgUejw0X6oC3Z8vQWrMXFtPRBzZa8JWhrssQ8Ircd9l/9J252qLUJDttawLkE
vSMZ+CJ9MvTK9FuQg7zGQdl7Bcilue/aYkNDJKQJOJ/pZHAGwXq1ZAYNYpwOd0YT
FfQsT/VNKtnd6GqzgmlcfSgFXcgw1a05GMFm2VjYn4HFull6lRI2h4arQEiNNojg
uPyq3GDChc2uoyASO1ZO+I/ihK7LqzwQAs97mv/dnhp4f30tGk6Bff062/Yi9+jD
EWQkDBNx5DhEYyiFcHSPwU4iH0bXiuysjvU2WFxfLfM389POluHnJqSJZsoATKxw
Vv0ijKNuUjuaW9Je1lTQMyuDFe4v26DIg3fbk5Sgi2RWYlPJXc1d4I0XLyAmNi1Y
3HLY30AnUnaYXVsWt6oq6aoohh7EiuSkSBKEVaw8QmIGVxLzalUYf0x86Q7EQGjl
GJOX+0dC/PrmmfR+Ld5S+BhH9XRtJP5f2xC3QxqRc43oBdvCmEaJXXDO6GVAeJRX
ZAfG7xWLUIf5rVL3KMyJEIz1bK53a7s7B3WHdS2FVeKGyVHVjIURi0aZW7w8gFIA
T/50wApUDX6Zx9CIizr8SNCVCgCc2tHzxO+lWpLXnmKzwGQMxoBw589hWnF7udjb
oAKIlf4r3Bdi4mwDWzdaMMgJVp6f2v4fx1EcN8FhJF4jiN2FDNTzGL432GWvCcED
VWvU5oYNAhQv9i8tJimbNFLpe8S1uziUjwC3neN0vvHbfeVPIxc5hmXivVBQj1td
zJGA7Dtk01ZHUeEPCVEOu3F+uKZL7cmhAX5bOX4Zp+vp5JOV4S+WL9GfvE2ZPR6I
hEO7gseSu9Si7R/ij4aJmLRQ+EoL6jMJXkGU4s7CXz+tUzZOrjAJ8m9sElDnaTnz
rtH9dtlL2kI922I5yoB/70XDazEQDeuDl0tHNdVfLEeVr5AAaZVs2XOzDN4HSTNN
7A/LK1Bu6qRSU7xSminz4k8sDfYUTJJvuv5bmLEuHMfG5Lap/FVrVPl1P3yvp9vf
DOAohChZ9ZiWqbTtLy73sxw59QhpdXyuKn+PBYS5m18qbipZttaP6/ZqTBlmZLJn
Y3H4G/Wg7L+ofgzts/GXD44gikpeohc+4W7CB3v8GgoFXocSwIdSmOmgZbH0XkdF
gvdGWARQNT4oVHgdL7db+N3pVkd2jmI0TW1Wr2pqQIp15Cj0+rCVBd+YeXJQaljY
nr3qhA9uMAM4QeKjA5Y2A7q8Bi5QqG7xHqJXRZ4wYmdtfw6tNxUrB33XnYJ1XTk3
JVfUq/AHjYgcOoN1rUaYX3/6I/jvJoiZ4w+oloquelVZI+5VrfjRDnygUkq4c4n8
HvNg+rlMbra8sZ6mxyuy57j7Lv8gWXIiAmKQ8Onolz6YB/H7BlmeLQl/vqFfXrCL
7X0ZaiiC7s3qpoulGRI49z1JUSew0V6kYHB/OPPr6Fpt9cNsnag5Bh8CqIi0UB2w
hHm2SdNeJikOXMJLlsyFYoBfCiyX6DhXXoh/1DbfcBFKnqAgakP3qw1dwcIrCgHU
ob8Rq8bzk0qCxuSjbJJI6OBL9BhD0TC8uuZf3xrjTFu9AskeW85EJPbSUOpAFQ9P
8ZGim62wKQpWJI1+XRTChSJgJtGtyz7yHeaPWfQ1H7530jJY+nFU3Zo3njYacgc9
4agXagM/ZiiH0DFV57T+2dfZkoW03q8VYAf6ng0WyUQ+GJhEhBZ3SilBn4rHKwp1
qoas8RwgtDmtl0m4nsuYjXKMxheqIw8nioX/u9aR3NV9efGKGhOlKrlKtGGF5PG1
g/1isNrAyi5NShxqLr7ffbWEfqqz4uDfLkrLDii75iQS7rWlXkhwpPj6mAeHgtyC
8I+HER10bmag9Rfa5kw3CMNmMcP2R2xWvE1tmI/ZbzwHmAhXWRxrHEW7N63r2uAX
kLfiukrbEC1xqxc7MVk9BsY1F3VQxjHJElW3g0oazO4VSzCmpJDmMoZe420UtHpQ
FSHEEGUMp6b8FkrN8884N8nJW2FxxrmVEQOrfZTW3ZCPF6x8rFYfUM6JMQ+zJ6En
wKqLWX7EmIdZuOeJDwww8TPA3qF297TL6Nkde5ROx6ITdtBp/kwgXUzumcgiiL2k
QQVmxR03x7c+t9Ncz7LfPQflF3CHGuGKNObXBSdlsJMjVBWmPkdrtCwrs3E8i6zF
Xcsx6fC1RCGJRJgWGJDlcZvRB9HuXDuuhQcmqqT/ecTRkOMCJpLrTB9VAYxCwfM0
5wVqs1Cd7mr8m03ePThK//ddCWKVrY6HaCn6R4HPD0bfb6NzZDCtd0GOMNbgHQTr
3Uh41Bnjl9njrx1FnohLsQGTNfZrdmRjXmnFPjG64zSRRGddOZMnm6zxIW89LYYr
pIsqUdr8wg1vwoi2Eter9otp1XZsL6CSeXP6OwXVTBzMr3V0ENa65YnlRLDe9pIB
S42V5U2nR0H6fVN2RGPPaVU9TXOY9+Cu0qTT0WFgQpnfCXJ/aGyIJhuD/wpqIGZI
gzc7asFbRLfG9mB5jEW/IafYhX0b+oDcb67bC5k7knIbXb/43s95QT/OiWGQKztV
gdhisVwJWHtfXBkUfhMk/qGw0YFwAOwCNSO5h6Zf0oap0F0bgk87PNQW7gNFOwKQ
5P82LWYSJcWXO5GI4vGzdEf769gnKUXG+nzqLTtbHIXUH8eFqbZ7Uw+Lg3MxmiDC
VzwZcY4Gwd2sBzB94mqDt2TCpN2kytJSA0meK0aWSmTlz4aK+KVyG1Li59wb+eGH
iazemuJn7vvWwsr4dMVSp3TTb/c32BM4awml4mCzg+jJ97q7uxifKFwnmb5yk+bu
v6Yl3OJADzkZi9Lkddl06uGAnXUkg4ZQD/fS+cL6B7xXqGd63fv/zsJ2DoFD6WsV
Ia6i5bunVxiyvtmehtBcMc1aAfE8P9Hacst39mEWiKNnRuA0WRHLL67qucxXWOsX
e1D533Ii2fLwAat1QfoUQ2pX+7W2dOgMGPJIdLdTR0t3BWsdAD650nMHqdUCgfi9
L2s6JcW+l/9ouAUj96ZSftKW8Nmo/3TdM536hOZtnfxI7d+AyytalJVgAqSNdqJd
pqrSPar3Zy8+a8jurOUtT0hYYEd10rmuHsUVXPmODCFr7+0lw8BnEJNLnBtoLxAm
685uQZBhguiRMiRkwyzVgVi5VS+iszdv1QpeY88m8y9SQNhwUhggXW+QbwSe3LfF
RdoKpwiJ4Tn3ogWtKBUtE12LNjZ/B4vLMpqpqyj+OxOdQEBUt3wPH3rGnAcQHdnr
bNaE69BY+JIoRNEdKZOQVXWl+WnPYyZcb3dUFhK0Voq5W/CAO0WBWxc4JYqwgWyk
QawiqsQao523SQZW2rT6cYclBcqdHTKjhouU0FF1b8LwWsbVHERXbYWbP7EEvdob
FVYVMp/uTl/pByjuELjn9Tq8Ud0XXYIFv3x/50lpPKh+lZy4PKv8TdqbNALZVbWK
oCBqyccU+B++jhDFco7Xq0iqV9/58bcgDtmbvsvwerPRU6nRRwe97Mi8/iqO8Zvn
m8AO1H6bjcVI1+SKmd2XmB7n2Ocnv+IGd/eXhj9j6yWUNjO/A3a9aOSEEAUU3wbx
BkowRIWz9RMIlNpbLdwDLLjSsH6AeoT8/K9k4kQYomhR75de+X/+Qazk21wa8Z6+
A7JQFH30v3G2Fos1GZiD3zmHJKs7bIkqbLHMy1c7rDTzvYRbNXcP8VN+CfQxRgzl
C0PiTNeyvU05LLgKLNv0KQHgwTvScDuM6vdYs/RmPIn//vxEwH0qh36WDD6sBjLk
VKwYflcOywacQxE8ViswCDrIGDobNqSoBVUJJ0jqP32CL8OZ0PPrfTiF1p2NRgOm
vI2ifFBrvl3zOuupE5cfAP+jPS/gRMgHh0OsfNvJt+fzkH3FmfMw7UmqAEGY/7SK
9v04DLpIuJjKz/aPSYb3mpua1nC84/F9hmmUYUA4lz7eGCdRkX6lE638tZOJ0bIZ
eUz7sngPNrwwzC0KFCjGKPm4zr21SKWrwT4vn7+LhEFOhceTVA0rXwbAYCE0Tn7P
dVMNN4uDeVyqiY98V1NIYTlCK63MDT+aNwNJescRNVDDv9CP/AR+S8akwO/iLikA
SxYDiC3iWCc3n1ZjYGL9ggN57WCtj6viFXe8PAnwjVAFfGCsRH33ramkHdj4yTBt
QwEcQ8qVHhuXn/WP5IEsyQhLlpYwImlKslivRhl70ax1U3QnKH/1ZG8VtAthPwSN
bZ1HX0aRmxSpHk2i5FySNi4HOQvODv1aGo6NR8bgcgjDgr+TB3GLrPJh69O984CG
C3ddF10heiCYgTWWwSEk/5ptNo6T/HJKwSs7cG2thePMX4Sq1XST391fMqIKa06M
oVo9rw+OlHlCFl9kx7xj4La9IFJmd2RxVAzN3l9mXdG/g0V1NcQ0WE5C3NlIHXfd
ZR4GTkxQ40luJyPtagl4AcX2KqIu4VnBNL94ciUpTJKKrp9zLzWU3XlIE7ZlUi/W
ZSTPEE1rnyDcDABEG6OqBhrrsk1j5m9rOuNhDoZwqQw3/8vNMeiKsw41/qhF1eLZ
olQj3LAOVdTeSaAqCQuQBSNEg/rGWbzL/kdgqxbZkkWC4+bAMCQbTXJlDkOabPH5
pJh6qUrjRYfA/+kh65Xi1seYUc2CqZw3+wn3wkrSzSzvwJqfHnNZze7x295TIdg3
nmCzMVGIZYhbztQUCEKPXkrKnn97oZJQYw5Z1OKxCVeLnbu1UGT0MXdqkxC5SdF3
V01hVNBf31dxEUvtCxx1Kt3Aus1irpuGwWP81stBleWfla+vFLG4TkKksZCq1s4d
xGxbAG1KRIohlJok3Qj0WbwOSSIGdLS/A1oriVEE1wq033AEdXE63kKPTL6hIXQ9
+yhLteF1L1TPbfGdRzhvMK3W6kwutgvfexsoDOB3q37o5av6RYZHEI8M/b7W80y1
lPEqrUBHqdGOZQ2AgftKZ7/ifVciqhtf2EPQLkBLwGQFJl2LDSwAmpwGav+vpVVx
s2CIRlC5bvkmSxmaaq/Gvfd+xzd4sQnziU/X0UN5SLPLcixQJHWDbifsnRdqmIoV
aRSZOnAB1OymOrXJJRQGkQOUBNkrShp+Y1c1ZMljJCtxQNMam7ILM12UNluty7Uf
4Odv1cCbgZ7UXpjYH5pkRBExzH6zlxhyVuNd7+2PbHHymAwq40OLvp+wdkDNxTL0
1x5gxOmg8CA4MHeV5D19BEkEBUzUXO6xBLOLfHBN+9jv/4MDw3c+chtRgPhj1zfH
8F6SvpGH3QsLbzSQeQ27MeBMmKXKJ1tTHfUmUmrmnyFk76Cs+GhW9AoiZx9mcjZH
/Yp4uc9Bfy2kxOJgKJ8b1lcA5jIAyg5mq/coByO3xpXxr1XvWBxtLr1S9T1sbbFE
tsrmJELJo6V7Y6LqVXG8nlSQv8qtMdGsDBwRmGoQOv9BwDHjDYFNDJ8V1OOrtTGf
oZyb4gwqKEnvrwKFC02zaGysQHYxt2MmmR+ZfF7r/OSio/2EpXS+p34RDLiXi65T
mHrs9/XCeY6aZw4OFupZEhuPCI7G3yM0+GjEPvGS2RKGrKD4p3wOutg9e2TAcpy5
rWv1f/xjdAnVucs4wpnbYONz0H3w7cdTKUti/sdHQrMxKSTTeRHpjQElcr0mIJPo
ZED+CQcxWe3mztJPYuKbXCw7cT/Om58cKJgInI10DqeKlYk3yVg/zapx9rikrztG
mMbRYgQjAuMmywBaARzRjyYQo2xskeL9wHZCahDIWaUFX190qgxpLybbFlsNfJW0
8BvO3/39xdFOJDjgjiDNjzgMzgJJ9n5uw1FJpgKWTTaF7XWQOtfSZUVepdU+Fkx3
ElUh8+Ye3MWIoKeiHeVOKHoXgmXB4eNxfh8FWI7TXSknpd+mA/VQzVoOnRViJau6
kKoTMNPcOXEb+GjEP8eKsvjjqI+q5hTK0dFO6Y47wxFpSMdcS39ujSAli441e19T
3cMFSMZCZQ0RgIH9laY6+C4yNVyjrMNJxGAuIsdZrPnFDp8WXcRlhvzwVURtul8i
fje082wCWvN/3GydAL0GKHaFPBmsxcTxAiIC0V6oMKnnjyWSC15tfge5q9CDKcRe
XHauJwJxims7tAcdmImJMtIyGzij3vDc6XtsQ/YSyeUkjrAsDn4G0Ru+J9yu6QtB
DJgVstlk5Msei28njOsVuPPFUZ4h6HeP3tZb8E7f4+fvSL8vGgOeyy6ARMzHjhTn
WN1bcUMLjrfjrsiwXSHn/2jjeRNSh40OMwqB/5APryCeYgK+1yMPWwbgX1BoDR9V
RIni7wnuiEOcnQaGgLA1/wa4WQ43B3q9LanNRTA2/M3z+ktMrcys7AjvWPgFqzbT
eF186OO8L521eyw0jPiqRYiOSO5wo6OkLXEO3P8NhhopD3431mDYXeZL20e2r5Nc
fYHCFE6mBZpcipuu5zniS7zRBjnqFfTk1CrIpjRS4PxOsVopS/GUNNqnXV1nCEGX
2obmwXkfCG2QnUZcNvffgMwl30oy32aSnCg56SlAvyL42IEyb6C0absZ1GGfpheS
TAQ3wfZkxHuQvQaEsh65QH6h+IgOt77s4w+6YkXjT8qeXlX0KWM6jod5kUvcuSPc
rvbSgiBFzBODGHTHWF8BDzmMXQ1YFCLtKyt/s//H1h88qVKDwjff7lJNdmE5WSWY
ri1hPyU7bCDzxBMGLi3Bezvg95GoQc/cwR9SS/blVTv4txlSMfBYzL+LxmmmlNjK
kogr06Otji8kv02yIinbyCA07wPzOUu1m/Ss7LA1xYhxaEafRRugjwFjC7f50OrN
ZuDbe8h0Q18sJ8TOVcqB0zjouNkk4ILomlTA0EFZed0EFArodB96MmjRaUSM01Vw
Y9QdcPI+JIPzJlCgjtVL+u4E3+bvw6FPScvHduoTKaY8j+pE0bDwpNQT/yrLD8Rm
hgfBy3KPajHmUJ8vTFNfuun9EVbjvVa+bujnNEjhzGFliSZ/a1Ka2+xpbVgDfm88
+YnRvF26K9fsNOswTzW+PWUjGLvx2hTp+Kw/bGtULxbS79cG+aD9UNEBPCiuGrzM
RNcUazOdGERAxWeQ/VTtAcXWGZO8aIqwkWn5ydsbLTWrRk9uhv0TlSRxy9oeeBUm
IvxLnquo8AVXS8yU/6hpXPpxGy6502TAxO/wwIX3lYdw6V/M7rs+aqPhAbo6BbMT
4ueqzKmnTP9La6UAArrmNPjX/0B/eOSXAXoXvFb2cZ8UoeESXe4GmgLo5mXL1vGP
hz5dB6tQe6Ipxsn2KPrtVSt8hE8rxo2w7B+iTAq06nomszqyTMiToUhl2F4swldV
WyZ79uQHu+myppVQKwIVgFGSHSC4TFDqC7vQ3/nkryHcxZ3o4PRKgzcW5cb+TZ4B
+N8IK4djggl/fvv63yVQz1t7wdCzNYT4VcUWO3EVN9X5uInNRYzrRbl937cC+/EI
8i05tM+aoiYxIr598O7wXEdJM6udVp5yl203EBhgeN75lVKz08tJQM5V29StxTMM
ZxfunJ9nmpmRSaaII4W1B6p2sO5hsNATqDfvTFskc5b/8/qLVMGuNxPwUgaaBLFY
/jkbNuizam1I3TFyAgled+VLPCQ2a0hvl+HtS8Gc2N5r5OARzvVBcyFEmJLjiulB
mq3O0aQWNKjYcmjw49InYK9OBmoziqNjsk0gQxNdLgnFiZI60QGs/oti91v/Qg7F
S+8ok0tlcLk3zO9BBfKFP0qYqCPPzz3P9j6doFOgrOGGtebKcV1QFzfsBsstZTQg
/dPvP+cbS5kBRCkBHGoISoyHRFZKkNKSLSgYxnVpdU3L7UGz+9zP3tIGE6RBCnQr
KlXAks5BixUuC5N+M9YJNW2I2ktrwuZVRZ073raAb53JfxE51ex1GaIF/t8iIwhD
8dP6Or3v8eiDVsLboMXQSpogKZkoF1bbHIKVPHwCMMWntYGzt9e/lkHkztL8Ruvk
mtcXRkfuVl/j68jIeiuxyjD4VXHhTvkT6oK7hTDY3QBX/p/cqT5g5jzXgKhKz/jt
AK1hwdhYl3C7+Vf8Y/fPZfKUscXZNk/mXPGhknjBrGruUno+cbwcxAmWZfgkxh6M
sSaupiYOVEvriZGvynvUb09YK1fHXSN8dc8kPzP9RwpsB+oOrFSgX6KlbEpWuDI5
szfEqN0nc1ZmlLeeqnV37bH59lHplQ29VbTjlWtEH54PRnLGg48UlQh6e1owfLFi
qF9BzChqSsFRKAFJrOZozeXjuqssDhpaaaFLmYHa9GIomTnMSt+FwPMHpu4zFxeh
RvnY0lSWYZxnzrXQciGLGp43TAZjdk+/78oIsH9NuIufCbhD2WBjJ1ZfA5PW9eGz
HqbB4BHHuW3SKnom3IDjri8Y4JPEiks6iD6xbCpLEu7OuV4Pd7zwtdwjdXNysRTu
n/QIZpR+RsgHx7pOlDLe/UkQYqWRReutGegs1oUTeouQQ8fcpi2qQbOTMduXNfKX
adJ6TIEt+SiC3MMDTZOeWAhRe0Cffqf78THYl0aIYaRYNSmr+CYM0ENiHXaPn8YF
vytFq21Ro08/RpYHmj9xbG98u9GzayZ27FgTcgkV9NeVnG+/rknIVXEpnNJ2oTBS
5yYiZezSBXg7Qo9QzKnHlNOWmZI66TOkLPAz6Gf/wA8dX1oD710lZKJzCsU1nNfg
8gQoeHiwrQfWoz3XwkLcNT8r/iOj04605YDMwZckP0VvKqPMtmGpBN+3TzzNIP0O
7X8771njH69+QNz4BcFq9l05bYA66Zjw8Uy17feXfjcoidLe0DFRAK7TOedvugYC
Qz17dBEyGZjgW+4+rRfiVIT9VKQIYsE1YDeUjxsx5Q+232+uASiS6vxjj7Vf0+NA
ohi1oP6fygi/CPQdB6v508xGxQE1y1TIlcoKwxAHrtujp+QmUrqQlc8SgGpqzfiO
w6UkvIc7CVCRUwszFsJ8nBa77x7L6ssigm7PfOytokJjVQwSJB+xUMTUmFcRfQvF
xzaUh++nAUszA3wdCcho14bZrbcFD0GAZvTvWf1py4z5mzTh39oBhGAOLMlAqZbn
1gYX4Sd7dHpUeZijuN2yOFAaMsqVJ0KuIiIE5vBBBxYpaHNwl15dcSqmnk3ll86i
bS1H+bBnDJfEhR5tXqgmRs3//xJVOfeBbALboTID8ObIkxo9UyCfSzaYMqxw5G2q
zO+tKHqLjV6r1kUkgpHC3Mbn37nABKahykeas5OEeplmND2IpBf0/QqlQSUXEQ8F
RS70XxfGA4hBszFdcctRb8r+XPiKaie5+K2MZ/5oJCulG1rK37Sn4Qftrk3+ufAE
JQo8Lgpsno9S2vEU/fEoR9FTu+8SGKGIVuepx/r8WSbNFTLGX6PJJ5V6aXMoPcoZ
ZlijPbjLypUKNFSsSie1KoJ+kYEbgb4t8BqojGyBqIVcCsr5usVmZJ+LD7RKXAjF
hv+mIqCm+Aij2SOMgNYKfeRzh0Cn85pgMHpBG0Q3yUns8ZalkAxQ6TEn7wDBoef3
EgIsPDnPIWOn3sXidZA6AuCnHyY5q+f9VPcjBC0Qyio3wFNyU99xU68y07B2um5e
QjrS5AHIR5+/64vydUGodbUPyOPyfZTn8eo3aOceLEjBqjZplzNAG6LL8GG0XeZ+
369BpbFCrzvaWUg36vrWEdw7FhP87aIm8ySFLthEAtZMdGBE8Bx92M0D91gfLWhw
MS3OiuirBg1MYSb0rpq0tq3FIraYeBbzMui9n1FjTr1aCQEDJAD1qWEfO1h8p43E
L3v+QrXdvEUEO2g1U/CuerdRObNDDOEWcnou2pvfLndhDrXwenAlDgOZxhf7dV2i
FpwZSDe5KRjDINv9/SCfoIIlHwcksYVqcjVaKHye8GizE6YmAkCl+5Nm26G7lYpi
Ydcl4QXk7BQE51GNSUcxZ3HaURldSP6E/GqXooudTMJqyrlHULEnfPe9dptiZFCb
qgN8Pfo5vlJvEoHcwdN1/yqkZRAeSPO5aHLgkUJho8ZUSE0YjCBEDapN3IiJdGTb
hsvce0peKUbXTZaZvbbfYG/JVNgZe7a9IcKg0wC1N+msZI+mOJJVsv1qp8pRuI6f
s2xDPS5Sh0OFEYul3VlgrVdxOEkXluMY96sCn6+Tv6phhfmcu7DFjOOdR2o/RiBR
2GD67iuxwCHxoUeg2NTOPzjJ7nxYGPQY6fcfG5JpKKOpOAovjBk4oyX0zQIV9mFy
fXnnS43ZjydeYGdFCUyN9atAx2+Q+ZjkZDvu6NIUSynHmHNYWY2mu98EpUgWWvtk
lM50jlhLIYyYXJ4fSll2LYTH5Ms+TsBYqVtMf4kcoFdb+XSyYoInajU1mpaNwhgJ
FXrr/1oj9BJAhZY1snTeCrhaC+7E9kGMU67r0M5meXMGJvDMRmXji/ROA43zVmqc
lT0y/AjuDZRHDL1oaE6SEIsB8eaBDfqVLGNXq3aDNA/IU+6Ujzp0kUrtAnqLGi++
FyLGMOEo6wW+BvG9ml/EE4LJI6yBmGuDBpP4/3nr/sulfetigbDxDlb7X9NskvH0
uMjfISzUHZi3nHy+8v7seW4JYaq7+6+f2e/BWB146f2jc3igbv4bBtbnZfamE4eu
+vUhsduXAvmcwpNZ7jDuwI5NzB1sIjeo048Cg/Igb90tGWEBK8/PsLAwAeAzLqOc
bzDZnaz3V/A3sWukYJGOi+7D/ZBRkiJGbjP0b8nPhTul86/zMYrQwh4u21Q6N2lM
7TyL9XdnZ1i6CwFNXRwuHfmX/99VV7g+GhiqE/a0jWu8SKUXZmIFAbsFD5yCno6c
38nkHisUc7J2gyGUzv2s+qJYZn261GaS2v5yiC8Ui0tZ8DmlyhXJiSNGQhnkf5GM
blNpj29Lk9lCiYZBz5Qhl1nHqLUr59O5xL6vHYCLuzAjU5fKJTNcFif6StmTk2bv
WTKGm5sou7DQzjVeZXbMTFvglmN77sP7bpyzUxrtn42/Vz3jt7hg5oN/bqQPlBxq
ziHkOxR9ExgKAXs3FdsKaSLc1+Dr2Em1zH9FU2Ohdxa7ttxn6+8xvNjwCflhwFGI
5I4/1D8yrkvrnvxbYDSdixiCe37k5pcbMQHcD6QwGHnxaL3L0x1u8TJ2mKG5WfcX
yFvMgS7NmytyQN4E0kBN0Wn8Pm4swM2AzAeW5KcZR13on1qMOOVyQy2TdXBiLPTF
cDe6JAU0dJOBtwxbegRs6gF2gTPFY2X8p/LhI1xl+FdFTl18nQuTSci+LE0dIR8c
T2BbJSu+OXKm3pINq+DgmkSrCgNVBobK4wTjnxnFztU2vTo+tEU3mJuoCqCyiNU6
mzBmlKT7n+fQDxGv7YrcuDcG4kQdD8Q+Q9BHF0gRF4lSo8vp284Vl2giFZ6rS0ow
4hhnR2jMdCzOCUhhjZ+Ofz/4C7T0YtpwdCqcnspud4UizQLpyWwKnsdAj0B4ls4a
QRTDbSU3AHQfGr1nizj2ePEtdWUfQ2TLd6LIVZ/ihQj28IfVrPny/TdKZY4Ll2k/
vNklCirrE64MCSE0dYctNx2YuVUZIkua0rTdCRRb7uai1S9mTb5Q9wMXK+EdmehI
OZYGkkl79VKNG9hBlPUrFxd/TTrWP7AhFb3RMKU1Zbr3414kNxdb2ALE6gL2VRhJ
er5ndBNBQUowlVfZywX9wLiDyVk1Xk+Kt1pi4tYpc49wZOyGezfpCloKhWO7mH6B
dAznerQ1a3BB3RU9NJdOzYkoxHsetzcr4nSR2/A7gx+HnUOhLsjMRIfcX33/A97B
djjZmlA8a6cnHBLOTYoYbJeFn4ctZLSWa06vGp6/mL10zyMiddZhKKLpRUPfVwPr
f24iMm7JSlkjeopAh4y5xVl2HvZs9DSSXXgQYhY/wLitXYkRA8XLxqUescdXSLeA
8u4kE4J/t46gFU+CIEBr/gPiIv+WsDEaBQf5DMcqDf85tRG7qbtxWjDOmkvYDeYi
1xBt/tzN2brew4yp7yeMCE/YjxqnfiVJqfydRJyFcxv3fpLAbtO7X/Xl97xwikam
L3ZmaTGVzRVRL0n44SzQIUtHN/1eaFtb7hEVZLt4WnbA03wpt+9a7lGn8GzgTLm0
nzda1BnkC2oGnxOc2ud8zRjJzDATOODNzqPbcxj1pvJDnPcDTBbhVROjgI1QUtYr
U3K388wvoJKb9rQ3vka5HmVjgE2wOVJWiEO6lvJjnuUn+CIkBTjENaDSLMosj9R4
np9EQJoGiyC6uJgJuD2iU31grRPsOan6qJmmi/JHe2iEZFHzpuiVP25UPQSdTFI4
zCeQjJnY3CSBoefNsb9qk67txuqqSJMG9XknLTz2dGk9L4FMjUb+WKNp0IXCAmVx
tljr7BQ9YkCQXtAFwnWeX7kNYjiTSn/Vo5aukrowByJ32y8i+NFIiXuApJMm0ILv
9xKJqSKyVhLKC5gSxHLOhF/Zck7dtl9CTK6WqD6P6+P44BN4Q22njRbfICRhYLMm
yL49dTbbJBWu4DTGv6Xbk8La4kbczifiEqQg1It8rVhLVaLyPn8+2F7NzqxBd2YO
51BU1AK+Fo+gxOWZNb1vaUIYJ7/DbbocuGLBmltoi4J9lwOoUk8pkGpyKI+wyaY/
nkm1O6I6RtJ1UEiei6+gjf7WAN7i9R0+hbOO/Q190RWP8tgvVIvUvflIEHigQtey
Qtw+ObSuky+yxjLo5EgS981Oc8/3E/F/sYl7ExhrbvLJZHJIfduKpaf6O9+iRguY
WSoN9buLkRFfm/k1mpgVI3U6xdZGs8Tzq2WldSvaDB23/7cSZClEaTo/0NQu6JDk
/yB/WlDo70gHI9O7v1xHqryf43LaLYm/oR+8DqgtjkXrHXyZfqwtFXqZVNBESCKl
uZ/EYTrR1s9TRuTodnT0pHJcaxAeEy7fQtQOiHWe3chbfn+J8z7EFj0457VFrbhe
bmonf0vqXtbxgyexUaDnP+qkjts4i5b9KYx7vVT+Fg2r29dQ66h9F4WlOppOSNoa
Iwi5OvSqHG10Zy2a7YwuXZZZOYDXH7J1CncoLmNnwHl//0FIKAOxuqFfANGI8jlx
T7HqA6cQ6Qy0pG7mJn8ctoJTjzkcIkoyZmfwKyJou5s+MqKW6cuA7hWUNfdzR4uK
6Mz6fCe7MEzNx1slE8mzF8Xv3Hg6Iz460GwwajmffsJ+BuMaVh0WKdQv1RjjA3rf
iO0tPxoC/RvR/jQeDiNN4r5RjIJ72e73p7jETQgAblekstD4T6NiojqRkZJeXt1j
CYia10gWrUnwdBjiqTvVocMX8dqeim1CPaf/YJRMQrOjaDx2toVU+wPpY9efDmaV
D5PJs3jn521o5S9Mm5ecJt7OQ6B3+9HdLcVtTdjP2Fv/sQqy56BkcYjR1TES/rsq
W3GyCer2ZugbnX8muEcM6i8CYsfirSS5oNCe7sBCbQ/NL3g9zbRj8UD3rKt9zAlP
wjlTHWopTvoooL3p0obX09rKryYTgsrWuMj/bJUUiRLll+oHrSKzJCn6NzZvmjvX
w28VGDvvWXVIUgWvp5KQ6/SWwSyTZ1Z1NGOP1zgIK38ZhpF6VuwYuSUzxHg16cSB
JSw77H55Ny6dZL5j6QxNcmzZaCAm8coFzZhqDUwXhUW2dhBimiCfaLsFNx28PVGF
4CYJGRoWvXp8dZThkeB6Dr3OoIK90A5C7ZSIb1YZzJkbve5ZL6kegKVIidmuf3Q3
RAU1fsBLJ72AdaSxsOrGOVCdfg5CbEu0jeCMzgOnwt1humELsv+6+R4wxvt6EH/h
xjr5pZpVJwU2R98kBKfilmKMHOZVRygr0By+8vGXtrBX0pwvj9sQsVhRikiKG+0b
JjNOyT4MUeyiENpBhaxXAUKW2yxWHCEI6xs4d7+BqqvbSxISeE/tIx2qH1K7PGdM
A9/+lHkB9syvlHMJMm4h0qu4A0115A6QOmJ/XA6SontuPe7to+IaBaRrleEtCRBO
0A8zC5vwauHT1h8hgTgpmUWKCPYeTzLnFNeoBURp+QwADFVLngv1vemyD1q7BsoI
68Z2t1xHoBAAH6uAYw/V0608bTbfwz3+SbUHd2AxYBj9eCeqCMrGz7PhJIf498tc
pgtRYZfZcxqQFruwUHI09M0pDXAjj6mAd1YUrZWqPePLHeTyLuYiNz/mBiozL8C8
mys3l6Vgxo+WyOBFsPYApbfbhGGFiyYTCbjF8UMLMrUL8H9PCcM1icvnRdK+IZZe
UOlEbWtFYS+5sqMW4slI3VW1IhzDs3oL18neRybRGQKoOIv9xINjScRGYRlz2p44
vjjB9lyYnqnn5l0sCL7ezdhN/lYDPbVDiQ9etZ7xjdKWzRxJnnqQ1tlpm/F+i/AN
JyZzDSYOQr9qjZKpza5ualg6HTSGcmA7OHhupIijuR6PmIw4zibpEcxkt87aeHLv
h7TuOdA8urykuoPPStf/kK2MJItiEC2yF/CIS0W7iPUZOZf1z/mWV/bF2MwV0n1P
quC+c+AkLevaB/tiGl1OYWdB2nI98WiJJHueDLnBiCc6knga1F+qmx3P9zAwKLPr
IVmHY07l3LqcC87TU1HEVLNBD1csPJNka7BaAiDHitRV9EnoUTm8nFYDny/UUIRn
1GTwnvsBxO13ovDA5Zyh/w8WGMZ9GsxV/QCsavZarSyG4Rtp/uLN3K3f7/48TEFc
wHes8Q88tpxBBI+3cCON0F3Yi/JIk4pbcKMRIBroJd/vHSJAb987smA64dhfWR46
EtBJ0fffCkdZ1nLLEMYqVxvHfirIeIXqZJw/G+UAJI86Hm0NVoVPZMrwqv2nbfUR
Pn9Ejw3f3T2U4seIwiNiA8IqFBlgnVKe7h+pQuBLOpPv1y6g2dwwauNOLpBLqxlG
qhiZ9fA9+9bF1x44LmIipG1bxt7sjDr7wcTu4MrAbDZnqmWV1wJimCG4lsi2NWuW
zgTiPT0u2bH1cfuSf3J29ZxsWQ0XjyGbq8GSsxDmHMphKzulL0et4UlNM1JX6OiH
PbcU3JEScVjjxaVMPPhvdnw/U3p5GN8OqMWw1oDknSeF3grmsmFR3d2sbxCEsNf5
Sw8d770sbuHvWqnAWMuu2/qvp1xryGMC3kgdEMiunfYyOlp1sKg0rBcE0DJpSjIl
ANQpRNwIw7eUtmuMAwNLmBMRvz841f4NiPF45o/FeSmw9PgWiMg0IArZAmd7XrnN
1DSiNVfR0BTOBRgJ8amqYWWZz6XL354/6etnQmJhoG6hIX7Zjbz7cq0QTfFqrtY2
5eypMLw8/Dx1uRVFz/M1GQ1qY6Zc79mplOrcAFC7pCymrRPBT0N9TjnnBX1P/fVR
cecqHWGaHwLNT7ZlYojHLZdpsbQhluvc9yWRnvHv4f3jjFgnIJ2WpOl/+WFCwqgd
bIlkYNBnwEPaPsjLUrBc0Dn+TqVFooLzA9b3gvB6P/ePmK17SStBh7Xw9o1y3d36
/T3iZmgv2pb4TVo5/0qqvXGjDleAZI22JPKMOtAERGfktHK9Z0VGuGJ3/MLud67t
IQCV/HOZ/BBt6mPUsZl6o0Fi+B4mAb0B8/OJ6Bafi1DIpb7rjhUiIxiu2aGs7FEF
UR6Gc+UM/W3F2LeiQgUyWemAzxDUrN5hQiAgB2FGBrb8+oN2u3tZ4cC3fPvMp9Hv
Z+KHF6kvduc4aZ827wKPqUYZxZeTCsNl/rRSJRIoEiqQOWydvmj4CRvqikd813wh
u48facjgZGDCP+WyVsnqwRGCys5N6uFDFIPL2arJawazD8rvmWc/h+0BJP4DVUSJ
6boqJRtmSM0Qy1TOmn7cktCMJVEczcmQGVD6aYs4dxdhESAHINRXKRsa7Pi9JHNG
GSqMhIUBjz0nH98Gbax4BLMfBOlli1XcxTAqt1zWhp1P9PCMgnaXbwK3H3v71ElK
3sALeq7X3dfAeEcD9oGjc9pg4ISjzh49uJQ7U81pytRkBbQv58+zhuzCH4XA556J
HgYd4JuI9z6yCVQpVg0QN7sLn/tAgGRDuXjYViCsYCVGCypEQEdFjpKWP1HnLEKV
OUV1wAGvs+cTVoXUkWrp/KK808IEXssIouEtZ2H9YT8bQ3HmVWCsQum4jKCcR9dN
Dbbn7iWi1mFT2NinJixlEX56Zp6dI0GY8EnQq1uJQIdcbtB708jowz2DlWudvK4h
TrzfY9r4rGM0YSSOw1sGAfpHhaU79GAJpdYcdgz/twcQv7j4lktTyYYG9tukOOO1
r6HrW07TQ1EtMv67DOH5ke0SWoqrT8a4jsoMxzvI7cQLiz1tPtPVzXKcOTvsRZb4
uO1tTl75FfQFuU7ZZWoNbFYTECaT4ePiWySZt7ofuaNFLiHHUg/n8bHwOCyN9Vfx
UVfx82bOFO/kNh21boZyiMDQ9xCvI5SOlN2QrI0gJGwjKt0o/Cyyp8ZZrLPFmfO4
zyZOGSVeljs8zl9T9WccWkAoWufFLF4GX0PiaFSipWxSReQ1xWglYz4cB9WE4U8o
1ahztHfjwtpmYAZMqUFgLpnPZfcDYm+HH6sQJ7n1EJJZ3pQeOFSiu9KdFSJw4kcB
EZCkdgBIwREAHtxAhKVoohRiZKCAyI1kYvIip/2miWIfAWRkOe969G06FuCKQXaE
P9mgUHaKPnzWzAWNvBMQ2s2VsQsJyJClObZiRjDWCCbYxMTy7P6uveaDp925O6LX
fXkj9JVEKzsI7LZZnLs93YoyXctYAr9kHKDJeaNqU3oIEEoT20vOmsBaLw5hMPBi
LgoNmgdI6eW6PffCqmwlNls+N9/6j4fXRlh7yPIOWJWhrv4FSnt8bfbrTMc2yZIr
Ql7USNRVotEt5kOZu3M1+GWjOZoK8+D5E4Ri9+3bXghi72GlxOep6tIiqpgoZquF
6+wfc+a08yrrHhMIoi0d6EHgaCj931r8Uptft3k7J01igBwa0Mjc814D8pmyN+2f
+JyIqdT6VdjRweMx1kv1I9XzfZiNQ0jNBB2qf7eJEhsUcDB2diNC1ezrqFqNyCH2
a7v0m73rg4WWcGmYmAkhuzQxm6r0ZRDSX2XZfQ++t/k7jnBHLAWPsdYQ4WP/zRr1
0OuOYk00WfSuuJvXGP4wEJtbxSqzWLOVs7lvhenK/IuQ/KVgpgldyEQkJF2c8S0/
KkUaJDiSHbQ1+5jGHOXvQ1F9j+5KI19DA1nz2NsiwCpp9VD+grDv+ACE1Mme1a4R
B4Bu5fZ2GEZcRVeguBrwLYMyJ1Rd/kxQ/A83PG7gbWLyFOQQHnx2tszRnPlCt8YY
HaeLDiFwqEVNVWT70+PkWsE7+beyF6j84aEWMu+5kYRVuFYH6XBkQeyE6cjN1oby
NHQ1dgyZX3sd3sGVXjAgCEPkfr23DoDlrTOApZS8sMM905QRBOVj362Dj09aO4m1
Rbqty25V44Ds02SrPJbwt2iGTuvB6yTOQISfJ+ocK2h2SdJDp8XyRO0y1LQpkqTM
M1yUttjfKoSQ6ruoTzxsa7Fl+/qM2D1wYASon6czLsmrD/+yg+muAImKkWL817XR
fg+QwzBlzpqP8JnnU9LqkhiC+Yb42IZKfJcIabNuqnwGKC+fOQNS99OHqoCXLnrb
c+isqPEJaGthL/8/ImOT8QNkOvxsijV9p8LJWMenR9YN8UBuxv9Q8UoWgNMdeeu4
JpoQ9uK8HTPP8RIRL7Zf+i9J+wTQxI44ERDF87QcOkR0G8n0jiN1UCBXzHj4u83R
HvA20YH+R0kO9jwgyHyq4Kzf+WU1WbiZs4L6ELq9FeY9rtDQW36Ssk2ox7Tkz8TV
QXwWVlTB1sBOfkctfbZdRqyL4xMr9eA6nW8o7xOqLIBH8U3YCx5P7aiWWDhmtiMw
+aRZeulT29fV7lYPAvXifRwSWYh+ZPtkgG5qAAAuf1iNCOogVVnvoH84itZLomTF
bYOa8FTYx7TWIZHcFwYJ/eyTU0+S+g38T01ImB9V2bbyemCEQvtTjE0cSFxz2jAS
6yK5x8gxZVxkt8wVXptYDd8KTWQz1PCuJphMPAcIBnY2j7Sen6Gp1cljCf7rVBNg
5HqKPf3KZ/Lx09D4Ul1DHNzXGi9yHBXlRbzqRKf3DygW2ti13O/Q/tFP/w8ZARVK
Uhfhh0Dms6QK61V1B9jh2REAcDK3EJ0tWADWkpI0AZxVkwqOTGTGuCI2aGfIPcnS
ZFZ7FonNx56xJDnozH/9xlj3H143XZKOiCE4ZP5Rt6R6ZXb9vBEyd0iWd6d4kl1O
aduUhCxwRrBpvBbcejduShlr13RVbbCq7O/b9n/1tP+ErbyCHWau/7Dh9RmDyCv8
8Koofd+f4Kx3uQDoxefoylgAwcIasntGt+6f/sBOMKqPUTJ4iKg/1a1I6Wog35Q5
V5FDdYYXy8JdxJq9cBL/r1HAubLP2FIcGLalCHcM8WOtUbHEqkw5N5aM7TmoD55E
9x/QNoXxIsKZpdTD87/dFk48e5Hzf6dWokDFgkBektkhADomEZJo8pgXfns7Ken8
DRYuWmagfRApYwl/FRkUJoIEtfQ8qGAjp2B90DlTtzkDMzbkUmcgo0mo0vxuXtiY
vgNT7EFT50Vrf9DkTDapoKsWAHMMVCGMud1ir4GZB/C56NSzL+KCkkqVlJMyPVJC
zIaiaVbGsCvNjRBejRoA3YYUCDoMN/9ii+odQdF0NIsJ3I4dQ89t3A6HmXkHaeLf
7M1fNmiSdiXLbWCdS6w8qRcRkbdGEhVYlrYmorCFKeX0NRvnJy9lsO6DbpFofQtN
cF5jVyx4JJmkfWRi7h5wIBxuLrzoZfbgrT3lEAJv6TZMz6iqk75hNUWKJFoBvHy2
MD4Lrfngww9/n14n3WunJh75vwjc0sThymmiwLaJRIfVkDozKJb2/IuyRsQ5e6Zv
qMobVWkVXi4tF/3d2OxV2KJynRodb5Oow5/4Fb+G+4RP1EiTEc9coOkdFq/OeQOH
wbakUnY/ln6pm0l5rEK3hhaVB10laz3TOQEJIRFSNzvSBU5HHdi+M887qo0yljQM
gHdkD3q3CGOBc5hVYUCt4BUz6jGpLYTHwKYkCjyPufp8oDuswvYzAelK9sLGbtpe
rHUM/YRnevraOlvc64j2Ms3mz2zA5PEpf7NdfncN4lf/4WuunzcpGuaLyMBgeYc2
vhOFgE1xhUJ3bGS5E9uqugvALayJPE2lBxLDg4CFZi5VgZLi7OZCr8+ynxetR8KX
SgzhBF//suf04kARP1+SQYDidNK2wh8jvArUU4qEdExstRkMH8M0ro9feABP+d1R
mdolV8wrTWtfxaoQDSWnzmqyKdaEAZk1Tst8wTJQVEpHPDcksD1VpVxLRIB75ZRi
lOPaF/Hb2OKCdfRkhmEcIsN9fe6Ahwv0zwshjaQgpqP8q1d8kZDvYOyVhXv31Ahk
FwsMXI15RTaM1JxbpaHDTnskazMMMP+6N2xXPfi48wvl3UHxlZEPoajl/EL/8bs1
elZmhyON3EIKDIbd1fJLL3TMhaienBkpoAbMg+59lqA0vvfRWZVk60Fc1Cp10yb3
jPnKFU0ZjLNEGXBOfwKf6bLYGdMUK6nUG5/Ee+0EpdZdqy+lmwjUPZKiLr+0uBE2
pZo7BI1IBvywnJ5bj/Jq7lNfoO+3EY/nXxMNff1RfeiWWi3xbLtKuLtRrhSm+iXA
CiTJVpmKH1dCfzgsMO9vqrQ1DCbrbr0WZssSlo9Q8ROluVRrHzcvSgdCVGpUtUG1
0hgaqLhYpQDeLg1u79CTOYQP9AmYp1VZz+J/o5KcmMd4UQkrthQnIa8hSReg/A2b
C0+KNf9NDTNgdrT0aCRBaiQp3FDeNUjv87/HN4/WbvuAYLd2gcwVP6ONSYTwABKG
ajjnG5m/db6UkXLOVBSNNqFBqj7r1FqY8VPOWpkArUf6wTf1QUjoZx3IaB3qNI7F
J8zJ6Yq9egPH7a1lidAkl7DBYwWADLNlKG0sDvbzPpWY4Euh6EfejSS97Lp4354N
3+8F4aQLWnQzxUAghYv9uRhj7WvyCUCigp0dffmgGKO1QGtA6SQBImFBL4EGIetq
Vg/MB8BSDrOg3smGfT+8sEXInSy3R1HehqzAOXKq09jEdWkVS/tfdu3FOsc+iAn6
znM//Q//xFxYwY87DXmTF+OKR2ANiZmsm/tRuD/ZfFh10IfBahmkg3gf4W+QjktA
8bZ9K88dqh6HZZnvE2guFAP464TTr7pP6DC42Ly1GFfQdLUcVvNnA9fukBjhIhEa
jt7Th+W1SnsDB45622FmMxtOmXongq52jyAQ3tgUUHdLkANYd6I6cvUXHmNguGrr
ONR6jEXkVQ6sy86IpE1CPnMCBvwOriVh32uXwOuAT7qXsoKlB1RejN4lqE34x2yB
lxpnpWf0S2XjTkKuETp0Iz4IzJzpXtHuO5UQ1y1K+OHjCld9QJbguM05tBt4apwa
Y4BpLFYF5/uYqMDwszLp3sNYfiKyKDHfZFKPbjUVp1Sr5JIKEKEqWN/i6Zsn7jK9
ESetKPm3j5mULsRRzrZzF1OEpap9xcNL0cBUoqvGaqa/ntcW0U4cjdzdVZ4xzcPw
LLoH8xzmfNOH2ci20LumRPMC1VQkjKxipQHBesYREJFjrVoA+MtXQKbRQPue0eBY
rxfBVNixW0r5hTZRG76zKdNxOYBultUKxLMlIRhjPj8h1yIT3gC8PMjpeDgZ9ybV
chCXqp9Vc7nFgC/MZhi0VXiYjOUTbih41tGBHzBDmwZCuGKcT/PEX2RC6rDtloL2
MzxYuka06u4ebj1Mmapg9SATZoQXtrWgcPa8HHlEpTDzBB11+JeepjLTUr9kV7Ue
cNhMitbaiWqJIEJ8CtAhvEyzpcQjtgxvKP+1okiXHUn/JgkZZPhs2qycWOxNvl+y
SB4zcGjCY2qtbvDBaLLE113Qc8/oe+kwVbN95iPLXbe8dB5tLoKY91G5T8skIZ1M
yawlAnjm6jPFCEpQBajNJODRO3R6EWIfzizkvQyL3yVZq+SuKO//STsYBS9zwuN+
b84+kd95oFi55CToKXgiUoIJJQles5PaYgvNge9pX00kPPGU4mIQG2mOHMui8plF
p1QdTW8L7SHmWMmVs5tBDoWqui9tYBVtGTGbITL6XQgqp3U2wBrfVVSETE2Ghoon
5ANY1r5hUkQiKyGFsdQhW6uwaelEUSTCOL3Ta/5teQ82577LnGs4LrXlpG5OeZf4
F1Bjb8WqvACSLa9EGFP+FMUTPNjVASvR293PqFFQnyaaE4iXRpfxMIJY8QHqFjgw
jPAOPd8Cxrf2HkT6awAJVl/g4ZVyAMcfOOMOrUSbqq4=
`pragma protect end_protected
