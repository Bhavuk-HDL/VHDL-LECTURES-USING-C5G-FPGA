// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
GiLGIGRIl13+37fJg6e3YWIk3n8U4uhTA2LGjNFQhLJ1Cvb3sZjs18Ki9DqQ+BUZ/TVltNW/41vH
/g9beyfBNxtjYkMzRbI4njp3M19Af7t7Xr4zbHPYnrqLySWmm+Ln673uoZmiD6eufG0vcb1essA+
0tfeczKHXf8hbEfkockOenqxxuH0DOx5EDRIRx5d9XaGpS9/VHsUBeeknpmsBUHuVqiNp/pi4Byp
E6mHgvqmiK4/gdr7JeoLRhVI5dImHOQs1546jeewx+11wbOxAOk/b7GOrysMqgzrVZCBEcckigVh
JZshKT/+F89CecpBNOleKnyWZ9X9K3PIDb/r8w==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 30032)
IHio/R0a98/8Rk07xAAckd5J9l+i8E2Q+4cFb3/wdsyNFFF2UnPxvGbjquvCug/ddzk+Mxuuth67
PyILPwrYHrqNxZInQt2j6lFb1xA9kWr6beL2qegwTtUjQTER7d4Xsx0pBz1drm7SiNVni7zBhh7X
pLSCVsQtDG/JJpSkiv175FWHscB8na9cVEBSg3pbyCfadzf0PqLT8vVE+4myupJ5mSPDJAwz+sg0
USglEb1W3kAW1Mlqx+EG6QKqTxRoUZPPEOUxKEcgp/q+bb1hgyvvnu2b0w2A4hUDufLGNPcG4TgM
iP4fFGB3ST4Bvwi2G5QOczb3vhUvPHWlRJxhxotwA5HTgVxdDczJnUuve4m/Ap4FiWGEa2hzGj3p
G4nKqPHtS1CCUXQJfE7TJ2daURq2IWkPEJ/PjsZpCXW531mBlOrdXBihcVVPWa+8A+KK6EmOlVBe
PcE0I0drdcCTq3rApRnXVhx8xiwdDrXsJJ10VzU7IbgUkdpZwkHkBt6bdK1naD1QnkApK6C7Ycea
3UtHKkw5qQywHZzr5w73XWKC5gZrFc90exagSWrPqDGiOMpm7VmbymPQErYDM6OE2YqXAI+EMu3j
9zHIxWxUBdEvYFrLbMfz7Kd3+t1ZjoIklFuUfDseciR9S9oPywwnCzSI1kyVLt53ZFucNF1P6orm
/SFTXwC+J16v331YJ2+stGE2soK19t4kxnjOjPLHXlHwgAGx0xi4BMHxAKeFszJ+CZ6C5+FN5lnJ
KRnkIw3FDbq1jVnpU8yPw8gUUhrOQC5sUHzvEt7jrCXdkFLkAG4AIqQICTEJwnNEU0gg5rXuXjtn
/p9DcPJwh4CuQxihgOyt+FZ2EQSK/PWQFkKvtjSp9AhCe/CsGF9FO15a5ZQreP+DQlLyiVunUOaI
4E/yDZvj+XfdIsWq8D0+3SAi6P/sLkAD5h7Jlk+J/tEZf75kpCXeWkPnR2VS51HvKMsmx6aZgr8f
DJHhVywZQ1nKq/gorJjWAmlLk1bqFfuuLt7QKO0SRdSXx34EA23HBF+HmHUVg1UrA9Ymh4RCgHg9
c+otmddSzDM78BwWhDSWhwHvYLI5M8RSH1yk482IvVQK2d1FiN4/F9FIor8CZYOImLstL0wRbB48
k1ED+6h7hhyszuhmX4oT50zstHjA2N+nFeauqJaNM/eVFTMnCi/+zzoBsJsBR4uMMRSykzg0CsFU
qCYTE5VMuu4Fgg149zNvPJbsaAVGy3XxW9jUbdZT1g4X3diaO2bqw5m8Kw30LwklaphlLcCQLdkU
Ox+1Zm703uppUEww0FAsGj/aHfqPVxztHElUyiokTCWX3piTJ+o7jFmp0N6kywclZ5jJonDaSjNt
by2TM+vd5fNQbWD7h4a3o8s2K2DWBxuGWBc2+cfdrq0n5p3viskSfKNOT9c/c1p/Vi1SOabPydxi
qAvJZr3bNCSWL6aagPvmjJFwYixbz/2yxCsay9ledL/wNhPD+6CtQPc449d/b4HFxlemchF8uZ9p
72CFsgk/etXUJbQbNOmuBOg7779ihuFoakAQ96jQCwkBoIkwdUzH1BaWf090f1Duim1S76tAxPeq
BZ2NHx82b9NAncZcctUBuXozomAYLdwQTohHkwcmCiygR1ogDCIaQqbre00CvkDFPvR8Yt5CaNqI
stOmP08NwazR1Wk0pvzdm9lTwsu/ZTtnTEogy6ot5EhMOUVdA7Akp9lOWJWHuU8OZXWaJAOm/yv1
/ctng6ceEoncyVJhM8JQFbcWjOxkGg9mRl8voLLc+a8ZDFW6BjqHXf+THAURKIgF54xFP8aGGMW1
1MbtC2QtspfIcKYBs4CA2QvnGo3i9rRB+uJBqTwspUMpUswnyHzJ3vSbFCh3K5rkeMB2NSziOZQv
d3EAuqpHFARg7ca9rDeyBcaBOC6uAjln2J7P3rWQNPZF5e8nfsODPAEGisvoaxXRUj1UekWjZ+NY
/6wYZq8EK1uOAoMqJPKgjnAT3wCtZk0ErpAP1EvYVC5TDXudQU4v40t+aL+/ObtdOO5Cp7SFXhZn
S6sem08wvI+uGW89U/VXlURj3ZfS6301OccFt2VZFw8gQii6VsYM4xjIeEN8BzVMnBtrulIHr7l/
64AhFooipfpsYQkCeC+oz7ZxWDP+aIEwnOzAJeYSS9k35I6X9CKuyIi7VSP+KbohKvy/Z4sDTfwR
aNOnDOn/yZ+8fcT1fbGX3qn8SCHcCsvP5OBTDX6gN/NYD/HMuEoyeA91DK2vhv9cPHOTeijiMOrl
wFKS1LAVjMyhc3STggYZXApUABCpL7yNVhBIAq/WqFaBXSwYKGV3vM14nuEwnd2b6l4zCYlpxD+f
nxSfj0ee+imbuNJvmVfiq5VrJChk7v7bd+F5ISKHc4FgWzziknctuD3sMThhpOw3pCbwCIG5MHwM
wSYZDYQGxRdYJaUIqYyocaU1MG0w3wQzjQYo3jQPxfN5RBp7bDghBAVVSc3nmxvZKheVzgjZhOuO
DQ3kzYRFYpZ0/Hwl2uPwg2E1XWBcy1MF/tuTSJPp9ZlvEspZqrX+BbR2KaSrMf8WU//Xly8iMtTE
nIvvgo0oOSnNJfX4kljimeMz+WLXDZB1EyuLTpm0wRq9DKx50UHP6/r+BGOD9ATp47F9Fn3wl+an
h9a0CfWlGNhSYhxpZqbH0+6GfcBxl2ndvlIJ1iIfU7PI3X69InKKU8U/+e5AXijtU94PqhEUjlNO
ayHikegxd7q8uyviMWfFzie4U0BmEF5aUR0bhIBfVxk9yslcA3BcRBHFmCwELSV2yM2wy0Gbg7m8
6ztLEJFvzq1I4IbXxSjD1Op9yywyEOs5FuX9KrJ7MHYrCGeWAfrhcKtVTjyxJu9bmjbtvochVmOi
5ykQ5B7CzJIMh1PtIkBtOwWYZtEzvRAFDbK1Xm07blgYBP7/Wc/lQA4kP42SgNmdlWNSizB/D0UE
+xfgUC4Wuel0f/ZNxxfk29soZmRaP06AUqSwARbGAe5ycyFNMTMq9QdkmDpaJZtBCwFZvtTcJP0Q
OPnGH0RBErp9ig6AlEPcWrKg5Ye7b4B9Xw6IZ4GV+h2ddkqSst4ZJmxquT3SvevtbH/exs1WrIGJ
FCSzVOOqyAWDTpUpm9SvHt++Rj1hjWJYjOgxuVF6pMpSPgalTw5vAwhWcXTHzcRW4oOrc9MGvFbd
u2+iY3RXfIozq2hhTygDgu4DjmsYzbzgk/FwrqwuAx7I+CBanBPtzrkPJGzpuzqGWCQvxjBRaRun
80/fuQ3906HhBWa1z0Zap79gK+asWIRsRfb+nEWBAR+7aLaUPxEZRGZDml3ba4cIYFrulsreog74
XwW9LATA/Jo+Eq8jSogLhGhjMTcTPmbfG80YCMyDD8ev1B1Gl1aT7Fj5/bSMjITLiXOOtUvIYSIB
qXW/onEspVd57uXP2R7n4fctmDoV6Nah2yTkEoIPVbixqh4RGlgxpseAqYhnX9kct57P+q8rE06X
GsbwlYltkIEcbn1a+RXGMVewiODVGNCHLOxK7jbWOYxV1hSQM6umT+yv+8GNqYxjZPylKAdl2llX
xvhO1IEgwTw0HO7mGdPD9Dvv4SbJEkqZwiJ3ZxriQmeNFmAqiBqZ6ODYdypjUyF1gDKvv6HovegT
UDugUpSwrEgqymve+YM/a1dR3K7gdQvd9FnqmMk5XCiKd/jvvodCjK6abxG8ziAai4E2jV5+Thkr
pFklH/DO9JN/uZGoRlViXsOFsNRn1pG9/bs2kKk3O85qWdgSbb2XNI/OhT3Y9Mn2DwrRwTgGB/UL
NcfejYydYIUmu0pEsXsT8Ps5i5U/FE7JvNTEyN3muTAeuwSKk/pxkxKJGfeijwTHpvTFQK9GZrfw
fjaILTT+lYmiCIA7fQ+1yHyKrC5LWyz5gG6Glos0l7ZsG6xTfjun1faTPGXbW9aT4GwaYaLOqviU
yi72QJVYgwulO89xgjdvtIJ5YC1zFij3xzaR0leJ0IRn7cXsLrIWH4CpBHOhoW8ycE1NQDssQwu2
SOWsibWnECSzl0ZT71gsmT4puK/c0mvS6H21UKJ+mG4Lz2ItbDl3XSTb2wS1wwFjGsR8n5YyiStj
PuJ6VkoYefF4WjfqlqknsoxTDmmbKp7hUnfX1KO+24fsNOqpeSvp66lyjsuVH4eIgxbiTKMRR6RW
4nljGL3TIl+7fZCSSs3NNGmJzO17Xc+Pa6fTICCA/mOLq7VHdklfS7niYLXBA7uL/2X+/9Bqdew+
BVi+mqpaXrmG+wgnVw2i3sTk7sDMstiUiZtXsCKOpa0MnXIgfY/ti9hILdg1KVNXYjmfRVjznkE+
iDsrcewhahZ92UhBT5Im05qpxZk3JLtSLdFIK+LrhSUFFCtAyQybmMAcaK4DgIhEQfjVsVYe5v40
WTKq/O/mF6FjsLZBFob1aBbtuA0faizUBACnK9Kl+2Agac9ibpCcYHnwNokZB0QE6znNhSzd7PBb
cLlTsZqiXENQzfQpDTRkasv746m+81RJQ0dHqJL3okB2h9jTeOIIcCtrHeTh8qN4x0Cj3lPEuF62
8qguUi05oazNk86XEJFUW6VIfQsUGBycbVIydRV3uwppUV8IW4OmKizXXRQMFmk2O8sGk3KYdR8H
WoGSonNI9gvMgoRO8zPx11FohsL9WKFV5GWOxsfZXDajHauSjqHKoTYnCXejYrM9ydIrFwvftmZS
RAkgNXUPIFtW9wxbKvYwu4v3Kfr9RKupQ68yOl7IuBvsZFLfs+TQCna1v+Pab+kyCWvZk03S+YtQ
OO6g1PrzO3BQ451kX+pZzJxBPDL+ayNjS3rMWpcAiB4xESgEhGsvq9J57Qo1ajbFS4RBjCXyrwm9
tPulkioHhpU5kqCp1GdxJI/5dGMlEbf+glmTLpx7At77WFCtwKh5dviqbblXGxBkwZU8nzIrxTcx
hTSYckn1zrZj+jMe+hnoNGZbRVjyMSiCkhtnFPdapC/J6bG3v2tg+rWOA8AxGU2gBf0ktim3rwdA
KjrIXKlmEYOGRhC+vhrV3tNSr+PeYh7ftcRFw+fsEcybhtuj/fxOnDcaucRQgyLB7030MxGa9cX0
JYcvPA6y8DmsIm4HmJj3aLT4t7MTeeKKfGRnMLqKqbz+a/sI382c1nueeSul8qxm4fFIpxKYVMn/
+Q3SKCZ5NF7LaprcJpm1LrZ0N+mXDAob99DJuUB82ij6FspZVpG6RXsJWRUQSMsE6JjLyZP3EMf5
0uGP9iCaf78MKmzt1Vz4FLLlajXYcNCln31I43Bg/QtQoMFzhsmPlWC+c67UTZyNn/PvDbCvCFQe
ew1x3PEpeUynjcYLKJqkuNhOhl0S+no+APHuvrQWNJFeBEQcuEBpw6tzgPUdw52NGA552RN2QCtM
7AqIyVx1TzuLKHbf3/bbx6jvo5R9RJkE6R3e93OlgXvEzXPd049jiAedjX7CoARDGBVvb+9Klhln
Po7h6n0z/IZAaZ7ZaBSRzvEAsD1LrHZ7rf1B28Kt8KwqMcwXbkz28OZdyX2YRBVRWKGw2JXpoSnF
Gc3h9zT33Zm6PSSMrD/3I8XRq024HvBtbOlZl3/TrfBrbHlxie0dqaDCGYesc29vXafQfGIU9Qby
WXOHXIYwCw3PYe2vr5gckR4D7FWOYr8Rkp6hoNMfw9+ZAMMPjjXVFDGwkFtye47v0rt7pSQCWEDI
YD2rFByUwMeLnfJsj8FesK/7B4V8ohRFEWBGDSWyvUqNUD3qvFNj1vNPgNOhMRdxgwVv2W7XwEyt
YuKS3dhnbU5J2EO44lPF+UUxRn4xplTOXT91VT7yn4mKkFSFlOI/mNzKVBdGyRb9dHiQ0190VzEZ
SUdLM7CpMorQ2RhKalxuwE8tiesQ4mx/u7ebQNS/a8f2BK141tZW4Wzz34mFbNHWgDZEzRF/nskt
dwGFfpvBT4oF9pEbDUlfwMkV3NLFq9jB+QAkZYFwWsEkTnu03bNG14Hf7Fpui/V7j+BmRVl6mfjP
J5os8b19lf+c6vPzNPnbJH0Xk2U6TKITWu556NiwKGnNyKXQDz0eWl+V7tSahxjtaOhivmmRAyEc
MSNKnr8rV4tVeUCgpZObOHQVxYf6pC0xwBfGjuPefb8eL+W+nwZjbiqSVpHuGIPlBTxvPgWTgNVT
RMg/KNLqOeT0SeiYiH0pHQGyKrwwNd22d3XV6r3yZzoUcPrDkOxkwB2VNmQ/JPszv1wrQkYISkJx
pakndIcVPJpgTbgbeW/xAc6XWen1yUw3CjX65Ni3E6wlVn7ynCUycuhNgbK5jAGeTbzYA2g2Ob4u
pqaXdrOMkwKah+Qzw1Moty781c/5A19IDxM6surEu+x8zgLR+3Y9PCa6QAYT4glFveHEj6DjnZ8a
BH8ldJFzxMA/MqRhnV4tbErRJoZn8+nXiQZjvrJEP6arLuk9xyHtwkU2gnCOODfzSANd1AIveYus
neVvUI0QHtbpJnA3N/fbAHKrEVkG14DSibGOodu/rueHWkGAFgyBlMNFYcQge95HEA8K8BCBk+dk
2R9LkiSHrxJ54I/fKbZQr+EY6Y5ARDWwH7ALsISY83WYKreJSH98in52kgL0dRhaPkTHyIKbdQkL
k0h+p3Yd7+alCKb67EG7p+Ya6DWzEZR26VHA+gSqqXzC2JpA7H29L4/cXoVQVFmNGs2SH8A6Psvd
2HfFydqXzqit9eyOpVDmAn+fAYzVn9PmgB/VJ5vAdeqVW5eCtjSbcWYh+2chYYjp4pFpkO/vWp6+
ztFoZsGhrr6CXWrk8cKaoU6qQBp0N8BYrV6s+hKserXGHmISgLcPE9Cwr8gvwfhgsPEzOafHH2bo
Comuvzeq6YVXBkN2UDvMfdcO4aL1pOQ/fu2gafOuMuJqdK0vvZvg66b3CaCm0Bz8bsQaeAhQO5JA
A2a3+oYSWcVG1shjZorWauOyZk4aPPddR03LVBqmJX8dBYIVWP9MDhTk16VLpWIJDywR/8aB9cvp
dtu4Tlw2bGrkIFpNCeQMaeaNoCKcBiBSQp7c4PtKUG6mbJP+H+hGPzxBsXmtSSEDL9LB78y/rd3F
rSIAikPmkg/fLyhJuo6ebhecsZxlFPRyaZsLb8lHzzPVh8A7UyZkeIHvBFFXiYd+JV/GTNkyypJf
JowQyDS/JdzA7P2uIkkVh5qwmRASpVZm2vrxN9WNYhu9UwTkBHhnzzTvlRb/aijN8VwoLKYqmauR
ECgnKQOFuJr0eaP6qhRwkN/S1Atue5zCMOIn4Ds+BXkej+rB8GDLMWCaeynvXTvON8A3gtDmhYba
aQS7Uy9aShozon9183FAOVCGxai6kyN86jUj1n4V1rrXsww66dPnCEOEjXjNhRMY7X5yvpoADtli
7obIiCeXHKIZlq6Mz2ir6zbdWK6Zd2MTrScO4Jxb1FcPEyGUqqx4KLYXFit8ye+xunCtZV/Zf4AU
YVOuHa3mAEUu0UuFw6gFtjAZ81mIQ7+5rCZ/Poj500cQKPiSukoirRVFaIrr8kaseBTcN9d478yN
CgmugfgoNAr7wmTpf+XpVc1pY3ny0kKQS/LDHe7+uyMwiismdRkZElshR6dPkDBJdA0cYJP0k+h7
dzQiVt+dee7xzD3FmJCKCef35HBcWbx3b6VvMhh3vNdHGLpB/H/nugQszYGenR1HPeL0mM9mC9Ch
08q9wMRzYnLUdbxIWOx26PyoorKKgu0MAxfFu+v0Dxx0aiWYcJc1jNLQI+RKeCxIHymkYe32KcLe
CXPdPKal2bVhAMJYPLfYlfhF5ohQRwpAXXMgjSwKu9t7rpu5tr2HsRahmR8GWFSs7coEZf0WTWq7
12chg5TTsoDLDXijiAAUOFZ/LA372IJYzJhDB6rYy5S9z9C4ozm4nuSfsE6NIZSQT/ilV8XXDXey
cMDxc1qnzNlh8GRgNnVnA21DoUIfaVGWYMs8BxI3nh3O1ygLoYdqae6uARf39+YR4IEHkMs2U9Q2
XiN18npeuXxqfL7lW8eptJ4GWs3cyREeQ765Ro8AbeSpRI+ixFuymMQpFXN7P+HzdOHR/G7d5gJ9
44ul+kT5xkJFy7vwrCRHFBBDfGnhB/Ecy8gljROiHZDgzcMzCTvdfaEnGRUe+o97MpcCzEYgP3L1
kFqujsbGUnZe1t9M6cOI+PgqDIxldBS3oF1q3PpAGm3zdXEpXLDUWYpvH4EkGFkmp7Nom0Vhc4Yu
eJP6TY9kamkJTMMpIyFFrsP+0W5v0jk6QLQpNwfR42qE9PZDoUQc7fi1IedfhM3iWmKFTlyIedPg
qkn0APmDphwmWciP7RCulKpZ3JZpWWi4q3V/6G+wU8G8K3YHvVeLmzjPwepbNU2dU9ep0Nr070X/
pCjfwlUE8wCeiJKqQas78sjP0i07FP15BRWV1d1R5vQ/w/LggvS/x+Xdtfynfs3ci/ZyUKCn9r4D
D9HNurMlu9TLssvaV2GmvqVtF8J9oipWbSl3MKAEfU/M6H10jHyhKOD77yCC9fQyvvn6XxCV1N+b
tXa//SUn5ZzIEbKnq6rln6qpRsjbxL1gwMrISa58L77dQxhz/+3cxNI8HgNTFDNcQS+1plWmy3DM
1JVmsayRvyhehMiJ0Fp5y2nbDEqiXPQif3/HitoMDT9fqa6I2KLOfltisStmc/z6nsJU4AdY3XxG
wFQvcygQXxsxAdz9/0JFxB4T1AQohWnPqE8vP+HuAhenssZGDtdBIXSLUw0lo7uWUVLjgYMfoFfF
FuScrbAr85TeeRCfkP62Y3w9VKpyWhEGEPiy2M6prWTiRuCoHxTVZRhKuHyoXRtLCS7g3hbLsBVl
J3wzLknw7ilX2TH8qKjIZQN51bRinO0KLYePzRQ9AOuLdhV/PXExRlPgrDeEVELgktKd8nqVPcrL
4wVnU7jFINmoeyusRrBYuYGAF91VL+lJPmxeeY0Pfx+IWbDGwFd56pa1pcYpNNNGhtEYe2Rn+Awe
lnFnJsiHeNdWSaZKCg8TVRq4HaCTT8NWmpB6Dc+qa3C3yl19TkX0OH7hh2qaKc/2OWLFzSr2YxIy
K1Tplkwg0QGHuou68wdb77JnFj30l+uEExe7qER3MwGXu1kRDxn5s/DmgNjjvUb5Y8Ra/RJI9YU7
2/6tHk/tAWdj1XsUDnYwnDNrJRHrSkz0ZmEEPSrWjZcaz3N3ZphlBQwbDQHTiEfQoTOCDGVDP1Ls
n7bBcUtL3Hh347Qx6aRIHozD0HfQyq5e/kBn/BKWji6B9ysYZD9PyiXHs7wmVgibZV/eOkwZ75wn
KZyT3r84/n5ZveUL6UJdNIEopC5ItT0F5q/I630HF1hQIt8akbpssjigw0Dv2+ZpSjYWPM0ZXhrU
P+0GGdcAoqgUvQ87K2cHZRBDgjYR4a02nYvCblIlIRXcxxhGYBniUGfElUuEj1OIZ4hL5t/eY3Ut
G/Wv0HpCbuXwwAA1Xwmh4lOAZ0QWrMBhtCCpZseRCTA/EtH+gNd0tGnL3fyq1Sp2PVNuOeWMMySs
7fdAOMmDAdfadBA5yGTf3h7BDe1iSsAFF07nxTGYIWhfomeaC/nfTf0IqdjHy+co8J9gTBW78lFE
wdNT/ttVcA0ohp+sViMoFPF8v7LV0MMU1c5gyUPv/i2UkQRWXZucnouxYXKNi3ucsc0umzouealK
kFg1aEfLSXNltV8EXGejYCNCWQ2wGwnoObYuY4qKIv5RoTkU8hkcFmOyjp60+SWIiHLKtO01l60F
92qoZvTkAxeo/iqm66YtVE+meBrFeKWPN1JsWvd0jjXwk7nbllgSC5X13EBcItQ4hLEnbRRenUg6
kIR7lRIFd/X4GuuuR5WdOEQeonr47zTnrbwsKO9jMyHIK6Nt7eCVG03ON/CvjOLQ/Nr9XD62lpGZ
wnENko04cyVCaGKeZaoNySwkcHFwK4xmiO2qFDjVThgU5DNWXh1vqkIOW82Ltyukf0aLAdJU03vd
RcGyPrqRfM//o6ZJ65XFH+2A34GH/Ro1r96vreO2xWVyP5DE16qlocQf5mWEBRDak9DZYcnlzXlL
9LBAmilD8Vq9K/f9XY+w8G9ojpI4F5XaVqORMfBnLiaqzREx2HHN+WDzJbD5I5/zTWHC4an5p9hw
awbWFrWKlod9fbav1Cpj59fy6NqDQRqwzQlmvP3DrfpxM78rwRALM7YDzO8l2unSc1qjmiuZa1G+
hCbC+oG5jcp/0+geG8UQKKlxqGGcgrWGjgD9SzBVykU0J6dVeum0V5MR8iujpUaLBinnddTFyc+6
nDbEOV+41W4Mj2iE6qFVSbHyAwKLEZFj6wFvg+rLAQYsef9kBDo5n7alObYoNcBAgoczuqIaAA5Q
S7pQc5HhcwiJFyJk5wvZkO2CxMsP3vyxeMHasyjgBK3awP0OSufHddrxBgeyMtbsNJ/kf1j+CNLl
/v67sk9KRj/RahlaRHGFDR9YF5dbho/IFg1DwaMv2dx71V7ciXdMp22+7UmxTcKksyqblbjA1ZZY
G//UbyxGpoMUSqtfK95/Xsm3cdIfRqpA3soV3Eu+dKeiDk/HRgBOMdYhUg1vKwlub6ayIlfyuUpH
Zx113NwA51Ub4EUIjVIXak4SuvMH6UWTqSrzqaAtEHPv28CTrHXxsV5A4/j5WF82A8ixg1XE9GpD
dYqW4i0QFu+LxYXMVuL74uCjaVLqqCQ7J3zC5qSp7zA29XldP2ItsYANlmo0i+PkQNbHtL85ySC7
y1/+cJ23EJvxASJFvjN8kzXM7pjSYuUYti1Kb2/hyH5sBnD8nQai8DnPFFX5FFdA1VZm0g0Xpn8O
NG4GjiujPMeeQNieQkutVP75DgtXhJp/vqD14EwE1Q6qMIndlDfIZo/lqkq8J5hDRA2fmvPxH2dz
kCpyX/STtslooiCqO0E1cJMFS48Dn+8LpzNye+z7d1XWX8A+qIWW8ULi09UZ17kHMLg1dAIfkXsZ
u7oYz7dnSPu0gBnzOtj7c0XxB4BM2onjzffM3vzhMgu5o9sUQfzXl58cTa0yyB5x0frvfTaZKYUn
lIscNto5S5qsB9+FTI9yYTEAPMA71/MwXMVDJtzBaaOSBIr8F4Q1TIBpX8TutD3BXx+59LZHN5j8
yTmKjsn1dcLQGHyfbMLPjMlkRL8dHcjTJqQLVMNq1po8xWRIxDLeEFG5D4f6SNsLO7MLjlbqyJCD
4rFqqH4h4acyWZzp5lKoK3JXwGbkOcKuhSDZf1jIYX/KJYWIIBcQclnzCUBJuFjCb+jKPKtbhD1+
/3/P7KWa4t6UbqgPw/kQXId5ye+qr7tbft45ZmDdaYx7JIj3oZWB4OM9Hu2Kw5YEr3btb4rgrGjD
3hSbK6jaiosm2lSTSqKxc7yI9GBMdpA1aQc3Yv81SgM6OF+4uA0/liqdjdjhdrHjX4StkSOec+uA
wPOWAgUglBicZn+YXKNCrA6ofImEGnzMqMlyrVyehQLNhTgWPqp2xYeUj0mAeiOnV3a8WQcNQZOP
tdKCgISJwfjP9MZCQbQE7j+TwM70rzpvrjSuvMG7fCtUUys/Hyq8lGmDnQ/yfVrNz+wre1yEzeib
QRmeZ78SsHUuRVMicf92TO3evepCoK1IJE6/EW042VU7J1owl9moktIsFJxYAt0HQNBiCNIxbOCs
OO45Thyl8DZE1jaYKFJwa1XJviRbefUGizXQuoQ5L+nMyZjcSiVGHLe3scoHP3W5485WgAQKGCqZ
Z6GQZb+ITbC5gQFa8aMchKltwVv9ZbLxLSEfvk6YNX77D6zQ9gktdTtKMjFwyR2acVhVlktwHED2
5rSOMjOjYbznACWk03r4uM75+Uvqic4gBpsSMNRUlasABQTzBWDmJtEXuUEHzDdz9A0CV4FOP8Hg
V1uvO80YKhXKXYF3EBuhuFnCuNENuSvsQzZ2FmOS87P3GCFjp5X808cmLJdpVJpZdjOTT7XZlAeL
FP22XNoHIKvJTvAJlOPjnMovOr/azQBC38DScK6l64eHgRiL2JE6tHCRYcY2UZQzZa9Xw6bUkWuc
4xDZTR4tpwVcZuRnvfR7vxGTkDue7DZy+3orjQDldk8t6DvAdqpD5UYlB/own5HYSFb8eZi22eOm
BE8qcVUZ/kHc4m9dZV12qK6f/H577xdADSCZJqITYZnxs/dSkPrDcMkFT5eOUF66oE/7vxdmnR/r
nJA/ZiUOqqYAnHQu7QLc3PlSrWf1gHBdKbOEKU6ffcpnfj0fvNiMzm6gvBdI9wJBo8y2pjYJTU1P
FOWzPzDEL/QfnLiX1/DbJJCyAt22eyhFABRczce0EZTBYh6PVo2PMs0rQKP2yZp+VVnqifNsuI21
GdMiKuEj4oXUtynUk22RrFJa1VsvUnFrzijlHPyQtQOUki0L2FYzA6X01TdLVj38z292z9sW9J+1
1LWcJwgCHs0T6PkYDBac9XpWrdhFLQDFYz69h8fsXuCZElNczJRx+1uDjND11Q/+2ZTFwUHcyTrr
lKo+4/an6naKCl5XeaqLcp+LmFJJH8iOAVQewRtJKM7jb4KxnZG+mPu8XTrI07ieQHqrztztyJ6H
4zWSxpmXhK8OdFftiR+2l8jXb0CZe3Re1wu0Rz8IW55pUF9dtXkhXAY2GQHoBvUCYuIK1u3y+F9i
ws5qUzCULi2R1NUMNtsKuGsKHShgRp9Rk91pzdyu4bNRiJ2iGi8IXeeu7eVjmqDNW+JYDdnC+Ql8
+eC00mwebPPENofw+sU8DqJfE+MC7OazmQqXa6pBb3Rn9/0lRZGmgDOqzpGa4owOmj/Hrfug/QFt
1RPNXfMA1xEtI6jS5c2rj7g4aKpc5j0BFiMjxQO/AhP/tF37TPsY2BXbLISabvZZh96IrHPWgWBJ
0hqeS9+84PRcYI72l19EVHSwB4r4S+qzFaWupTjukkHNdVZntloJG4+fslBc9Ll97z0up1XYsSae
lxEFJH5ePK1l5PWmdcxcr6JAIG/niHqcKU9gmJY3mMxGK6kh3zkY2ZitwPI5Kq74jL8HbgGn4vwS
baF7Db7c29wop8Fen0pdFIYZEme6NZCePKZAPh1Iz0MeMfDiUpA9/GA0QDCsGIBn3bojYXIoPSre
4MZDoFvytz1R6cbug81gasf0+b15zVBzpCqQwQVLbw/YQvHZpsb+YlQmWOOvFoJJ4Dl6DQAPwXCd
6mHHg3ZKgekeRaM9VnXFblj0bOIq+efEo8GS6EwX9j23IM3UO517QUBfhTDS2ts2z5T77nstDkVw
gGRMOVN9IHaEHgj6X62GPjCag1JKuV+v6Zip+e/IDKDdaKCzpp9Z/oalH9/ttI+vxyBsjaS2fDqh
ZDzqnu+LVym0kUme/7pLDgKssnrbbpj7CYXCjU6tGJYSMKeOFNXs8I+xDnflUvD2fCY60C8HS8HN
T2OvSFpzdmLNaN6Fa9sgCH4QkwKVpulLIPAHaTj1qCtb/0nYBGJeOMm8RjFEjHCgv3KYeyPLzBTN
VkrpNKbFUuYGC3ZGR5I7rM9+wV+q32esgRdGwXnq9hnF7cnS8nGYbMjrVg9Crqiko4gtl8qJvBBV
cCbBd0FAjHJxyUJvGjWTKAhhhqAWwYHLBQNpbQSofdvB/onsUCimkD9jbXCIDYn5G2sWdek1ArRC
PY/LEdWyoX2f+tUtAjaillXN73f4VKDhuOEFoPkpbFam8dcmGmPufzwpIiisPDRsRVVK9jFgpNwR
lNkbpVYYP09jNflYbF8FeyksFHR+220eGT93tl/DMnaWRIvRyZtPRmplNaAdMxruceMs+NIzJ8Vr
345ty5odyxwjjOqf2GvPIV86wN+hyZmuLPUTZaRrO/n+xaI4I40ErjFrZfNfa/lGi8+oa7xEGtSr
7zTIyIONZPKaLQf3Uq7dk/9wgcf6Q2FgvjootDIrcjwHKu6hXg1NCIjXDxuw98Wct3rdNdl/Qadr
wkHPOy4Q9TsAAAtNSIjBaa+fICBxVhFaLc8hA1MP3P9nD4xHTL8526OWb5vr5cdUWfQs4NSnplkZ
cDKM3zEWEoz+VuMncC2J3d3buZF9pxDfivfl1+h2m/SED4MlhpmrTzijsKWKLJmB/4OvdeV+BcjB
1QNmLuwsPcyu2bLEBPiXUslCbFURq7BRc1KRWzjxPn3tpEpBax58Cq1hqr64uJoROkyMt9fE/Vr5
1Wwu/CuD+X1WE0zHnBeX9/RdPSVmVhSdq0tKT0jHX8ErD3hgvrcLaqZtUax6Gak6xLfWN+2FRgxl
6JEpSn4MS8xA1tb+FcXqdLfFxZaiho08ANCxGjpxJKfBNmDt2xbK8zPGNfZXV3MxZktNaIpJV2d/
OYy6cXdJHHDJN+b+VagKXu2VSRN44vthB0dYKcVpjw+tiN7tSL4kNxAiNaLT+2qt1tZN+aPeUOk1
ZEYTisR67FE5hsLApyFqn+P8dxCnJJUKREg+jJsUzoyuTUscd80Qnyv+Jgv2F7uiGzi7zjTIllP0
lxNktZstLPGprFiFY63FtKYRfu0L8mFgffbLxbXj5i/WR5SoBV+HxakIIaSyiZkq62gkOe+oagt7
A4Amd0q+gCOT0LMcJwLqJ/hxUkPf1Xvf9fm77oNClYS+PYkLCQYtY1cY1ST9opmBnWdPVREq52/f
OwHqAgDNBW8cWv6TSeO6W9X4zHbe5af1t33uTLWFyKYPssc+f5q7lzYXT/Mdpcaugp09MoiaKgGV
I2IRCjBkQAMApJjP4YGKgUbPtQpdrrgXCom7JIA8AxS4NfkE3VfssoAyKmvGtUasT+fi2w88NzcF
+lKTlopftAsOfCY4JZiat1fZGd56zFs0L9cnB2noLZcam/vncZTAjcfYMDA3EVW+G9QpIxW9S+lX
K+1ASRD2gxakXEXFhg66gI97nB1L/ST3FKWIIvWYGlFxIRxG8JJgaF4OXpds7p9iCeXM000IZl2B
1mUwjXe5eOJXui8m8SatMlyoGyfOdL+Ls9Rp1he7mNEkJZcFaLfGb/eQ836kwQLNeJxyM6SYM+dY
Rbn/L6c5P8dAxLr3raL/mQMr0DHX5Thr224qi49f1rL9HsHWH19ptYnk7eZQfYrBsrFIKzRNycdC
gmziHeWlE3gnqCfxc/0eOn48swPlG4ylwXqSE3Cmi8++KDICSTY584KlOIBgmLZ720dfttGDjT40
k5CiCKOi2hRAJojjY8vTyxSeNilbhvFlDgKOCJdQ0h45SW2FHb7K3f1G9WAO3nG7GqAu8uG6kfiu
uUyY7mJRc+94svLiJgA2808z41FLh1s4D13ZftzklIpi/RskcChi8eoHCjyd5LqkNgw02uTAlQI6
UFyRU+Lh70B+/GgoxpKsScjOyY3jxdpTKzfCg5jNPFzWEPC9Vj4FwpNfqwcvivGfoPFrEs4c7zcu
oDETMIyfgWi/pPQfjv94ppwKLywXAh3JQXkoXQ3Xo28o+S9yxdAeUegCMhg6Bq8YjI/9QQ152va+
9bVDNx1jaANL+LmJLYwK6yCtzoXB9Oijh8gDgyor+wsA3PGOVbSw7o5rHKmZqCIZKSo456DgjAz8
Eln7kCM4+0aSMGqUEjflQ8sYUE2bbKS7NnWMPmXSwSP3m25M57LPqrvuJzyEDNxfJkz/l3Pqq/XB
veqESgb8h2CCo4HJZmFHykfbrZQ9j3UDDT+5gRMgHhKcbZlZglESDdLQNko/IoQAEC4+rN7hAVx8
U0LS/HG1wnsbwU1FnLfW7+rFv1u66ZmL75yl0ESoE8wF2qjsk5joW6xbJovq3q1O9vZXYhZLvBsk
KJBtyyL9jCH06SUa/u9WQUhm0w+kaNyE71j3Kkklg9MBPZkQURStr371WWynlbs/+mxzE1OoZoVF
LwRO3tBRzAjxPKdqheRgIuIoiZp5GgaqHZgfbWzwfiBezG8/IyWTjD2j1aXcONIbZLoLCWGUKcf8
M2JJQTj6vRcMDaD2/uniMZcyQtWwXz6jE5FuzpoflqsxILIyCWGZz/wBao3VLT1FRm8V0Z86kBxI
GoG/o5TwF9rX9tHZKL7FiYa0yLqEmGBv815qJmFwSi619DHA4o6zmF4g+57U3sPfl4d9N8XhZPyo
rQ+J9Eq2WhnMPBeI/sRYJ+vYLekamwxnBCHab+HDED6LyD3VOTuhvfiOT8WkleTOoRfloE2QJoRk
Xnu0SLyR10tcD4120zvFta5hmMBTfJNX1l+UuRDyKsnrw77ethlyYUuNAfD4rk/vYqfDVNPFPgPb
QXLwsH6sP4KpcUIJ7HhulMsfG5MPatgb+9uDOzHPgRe6RcSWWenYSh6iRZR6e0yJCU/FiU8hDQvT
vKlTCDCyaoK6R/F4kKBrBBZpYfXzg8u4uZvaE5lqgbXcwjmjPG2Jkkbey3P6qwArPoMNtiZGgPNj
ZOy9fMY8F3DL0cpmW3avYYc5HSlJnxGdNNpNM7lybUgSQVt9NUCjjrmp/a1eWrWwxSSr2VSJJodD
FiQCgvpscpyPsVk7mHjQGgxWZQa8vWQ0d5oeLVWzCpnLC/kBVfT8BCSlLWV31l/lwF1r3z2+SEqu
KbCAluImrdadEqH9LrzrkVedcsWkM12G2ss9UNrjCAEsLVmEs0gr1LoQ1KYli+NMLJ8BHQ2ZIwyR
4hfeOa8wouuLpoyFWY/xJbelun8xKmpLGQjSg1Tsl2mkeEn6FDe8ZnGUB8H2x/rZsayZwu5eXGhs
/7ts/lDmF7d1Zau/ljGcDkHVZNC1xJWE9r1fXLyaDfpUBq2cr4iCy1QT8txsWJshijKdtf6daC0W
SNfIjAwVhHVsFwdmPnk89+8EFUIiY0Uofdl1IkkQsHJc0mYMeV0H3qls8PiOl/7eUTbwfljxVLqV
gZDcvU0fm6HM6X+OCCIiH22Z3fokZKzV7fYyKFHiDIGjRT+UUm84ogpeEUxFdp1ijf4JVOsJK1tv
1RVHoKbwYoT9YQXAne3GKT3lO1+L5rTcTkkbM5aJsjgSbnGKUh0APPM2+S2DhRRT/nAdAvqMbteE
BtnoEuenYvNYEHqoBZh6rNkg9+OJXr/a+PTxeryUrjTbqUVqMIDhafJ+7tdem5G9boV3qDvYPVZo
Aq+GjZQ7j2FG2vkx91hFBJcLgw8wkL7jD93ySHyonP68G491t7sfu2Kdg0lzP2ES0S0j+bpIfx7v
cyrusfhmlJdVXQNxeAIAw9ip359ou2Z4wXO3SpJTsO0Q9yRPwh6sPigDY4aqPdWIyNcftK2q9Vhr
4f2z7uWEOoEB7rMPYYxj0CZsUbK1GLldc0ovSufVOgAvRFolQ2R9AuzW6UhUybpA7dDs17w4lxv0
w2Iu69CdYJOWB5XQgUvWKL/gJ35NzkO/Bu012OT2CXtD2UhgPCFKr5VUxqtvQXhTEKemxpu9OcDa
cXNxRXzOVyIpIiKMMHPHflEMEmVIhdAfAESwZM8cj8J/hDIpW2ilLwf49uU6ew80LjXROq8npp/s
i5fBQJIZiEZyJFVzjIgkJvm5Xy3DC4NyLGNFP7kT4nUcSYQjhnB+DVZyk0Ak2DupCzHsrAT67mBN
/aVapJFdwKHm5cRLnFLfN3OSCA7USkOrDlAPmX4s9/ei77ciuvB95qrSaI3UZwjUOULVdJjrRXKq
XQDgob+5AAXwIb2H63A42UWA6hwrZUzHXn+FPwO4wzpNmvMb0dgf/bUhmL3WNMkmeENntNhHIK01
Xzw+Nw0JNjggkNrTHY2KX7DFs0eE7oblpaTnyg5mv6OV2GVEG5/FBCa+C35Xwvy2mqADNuaF7+Ye
U9PVT0Jj1X7cTs1pWxA3wP1X0SZcQ+1zCSGR9BNa26aFwf/fzvM3LlpFsZWeE3gBpiNJAeZScSPp
Sm8PoWiWGs2DrGDZRGU+6K08BsZYZArWfvzxfysbPLtYt4+oN9CtD4nx/4BsrHjcQc500dlr5Uvf
spZJAgTvnJuBE7UhjSEc68WH2KXR3K6Q6oX1GdWBfBxflOjEF4ev8ASV32gX6cDnJK3dqlPGPxQI
ls/BISGZqxPptV9sX4ybO9rD9X073v+nFrmZm4yb8+WxKowHaUnX0nQeGo5PZQhpJWO33tD3rZr5
2GDNcrPvgJhR2s6ExaB/9qNZBDPqL0dLle523cDpoh9V0XNcJtvWx6u/n3K/mWcUGQnjQRN/N2uy
yXBjD6kDcAeYTOzK6rs23uWhP6W2fNoMIvfkNZ032pmmB6uBllKl5E8Dik0zLhheSMBIjsVxUYUF
7sGwr81ztEIquqx/w6etWkOxD6n2J4AVia1AFnwFXNf4IGGA6s9cBE4qjFY+id+D+d1W5ZJ1aZJq
UoxPS700k5JZzf1G4oGGSDoxFEcrw4DFeEjAN4fTQeK8OBHZsyW+Q/8q23gMFPLiSoaKQqitCY9U
vDpkMh3xnD6O+rdMKmN88zWbvbdWsvpnZLiML2VsaUhqAdcj/emvq48AFb+roUOA+C96budCt8tQ
UOIU3jQkR3uXud+iZ87+T9feR70CcHJcZqDZHce18Sbn6e5T6pOqp00J1MM5RC+M1D749lxnZsh2
FJRsvn8IeFP/ULhmxQvB89r4S74USUdyqY2K5hq667NVPJ6kgFq6zb0COpzRyDzyTTbUp+TclQUO
tnkdPEZXi9zvZdtIkd5wGc4ouNq16phwhD3ASDldVZ+oMJWLhcigUxVoynf4vr4ZbF0RKk5j3D8I
vYzF4rTH4LN/BxIkFInJe8qIYmFmPltUWjRQj7qBmEl/yPu7PFJ6Ebv7i1nhkauX3MOm27JD/KIT
qmESs8+PUFQm5HO8S0oy4obVf1BrsGTh7eUeR43seJGIZLiZDGV9i08BqIP52oOMwbAf7UGm9Eu7
EC4EdvWvYA0yxvBkjpwvCcgblwiqx7maFWrpexR79mEUyBpLQTuQUN6Jk/N7fBRDKXyrXFZdNoku
gg/gJ7FZfvUn4fvgToJu2fbEixls/WS40U4ibOesT4MG5dqpNc9clC3sak6BGjrYEoJPtQEYKOaX
yxO3vCdxaMbrogDuiyq9MmxFMN0oXxwYQ0EVEfAKvm4iXFS3+W7AYlHJU0AzCsMOUnuQL3aJZilr
mNXcwrSlkUDsjmfmWD1xRRfJUoUvTQNGNqRyC3V5JPKQpdRhctl/Ppbqhtk76QVWP9AIVKBiavWS
iUGVhviFWJnjee+eS94gwPmfDgboGmMKfDx0NdYzM+BxNVuQPeQBRF5CNj+WB0wJtplkzwWTsguF
XeF/lGx2/R7MnXWcqBaKHLpEMvL/JCBo4uq/qiBUp0F0r9Baj4EqT/8a/hsiBF0dLqBYModXOiQj
qnVIq30uFnNuBHjyZ7qEnjLjK4NyiS5xfeP3O8sHnfjMbNf/c5PcOVx+RTic2wIiqygwxl1DZshf
QPGigxLJSH00ObKqxF5hVlVgJnbz5mtL8B8PvMqWsWNlSqajGqFu+4TzuiuQJVjeEl9yYHCv0j9H
CoHCOwOKnXcR6fO/lqWorIdm1v/2QlW63Zytl9YXM7vK66FsNNRolYvLIcE3HfIZ5aZNVO67zHMV
PZfwIZPwbi9vUfFnse6tCCpMUNSuQaxW1AmmiO2gJ4hZH+mKqFe8A/WtizXaTVHodYVQDS9TLeZt
MARCclq/zaGIMTAJNBcfXwwJhJ8FV5VOdJCXb/uqLhYNxsZXgYX1+9rzAwMb1gHPApYJLNxyujCp
uFJTNnjzpyZIwfeqlUQYUCYop6R4rnBOtuhqS+9eWw5Pa8l+GrdwCOga+0IEhXXMLqB9NkhUNts6
t2cn1a/MYhkPlNWmG4XjXDOFkj/NxO4ocYrc/uYsSPR01BwTLItUTjm6y20GSPhOlzFMtfMNajcF
SB9vYDoN2L2YZK0GOwGIxysnTshKHNdqvh5tSlnZK0iwDc6DcP1axSbAQRJcoskSkuzmzXlMYmgr
2EjFx/HB3DaNCcqegWcQIwOzQ5/ox8uIP4jCuQ1JosGNgtfi+Vc+Ik4kYpQH5IZ7XzPOWqIlCI4O
N+NmOfgc3qQ8cXJ7080yyPMxm38hvWZHrqtWnGfcxRS6CMBc/AU5rskLOzH4SWLOGlEaNf6Sqz/M
7QQ0Xbq7YPi5+88Hptdq/cz2CAUN0OeH7FPxSqefgREZ6qMvwUni2EmmullaHOKRiOQoCnGiMqcv
Vn1pmMuqAOvlA8LAIXqp4EHfHL0LmpjxnaFytPo6VgfT3VaVpn3rlkrbB+QLCmNZ5vq7+PMEls6m
bTwPzMUYfCXS+kE2pLyxooAnfg2z7ojE6f/ub7a37KuSGpIZRt36/CVOwyrTFLuHNA+n3i4MWOHf
nYU5Wqg7oHsVuR61xdlZ4pO37Vidwk3tRpMTTZK9ST/t99TRHL5tVTMJViatIOiIvkVBHhtyFjys
8bPc6/OjCVWJfJkSAHRbMDsSHDoCoNTO2WBN1PJgvCKt3tcKE43hvGvHsIaeyIH8LxC8916nFWOH
3OEzcFxQI2VtqZDZfVe1Dv+qHsYtI6lENu9F3UoXLbZTEl3x7iAOazNIrbzHTQWAMvmR8NUWRmNV
VkbWk01qwbVPxHYCaNegcvyuo4KQXAoX6Hqb714uC6wWmq3enmmtAJg9Jw5Ur2ekRNWJCwUEiepK
5WgPsZQrdLG2sloL7cNP5ZdE4oI+BfaWqo1F1xAR21kG8BiE5jR8u7G5OtWVoU1RwcD2Jt3rKSGf
JEOPcMPWf6Wsm/PnShebvidiVV0u47xeF69tUV5Yj8X1GlV9Z8eCA3jWzGRA3N/kAy0BpZBAKxAF
+cYih7j8RUpgw8GwJRynGcy6Z/IuPshoSt0qdrblbIJPhBJA+D/LLfnakNQFTuOpBngCVJPxpKRC
9pMMNFW7WnAwogHk5a+M03THmrtzgs0OyJ9iWrNTWv31mgxaERVAy5gMj/NPs1nf/IWdqqFq/ors
Idbnpl6UCIJR+CIgl2xAHGgdkB8eQ23yMuaFwyeiwcSIPHqjVVax+2V8a4U1MHBknT3EJTMpt31t
RxLumA/iBMizLc1zTt6w9egnr4TAB1HUyrWi0HGYO0Z4wpjDBzAJtQ7enhCoqh7Pp9S1v0Gy48dQ
gYf1FL5bDKFMcx6G7AJbwn3/wkY2n+rwgDHqA+riHRqF3eA07gPd4bDRh2IG0SOb0zoARfBOA2LL
tBAJnB5Bz5+zkO7CaUz+zx6R41yKEmLvOefuO/beymhsOL8iaY303zezuH7DC2zvCwfbLl2Hy9Dd
n08sr07+VFRFSHBP8thZHKJn38HynUOVCep8KCWQ2kA5NghKp8oqP+ol7quMSVHl/mrVS9+O/uye
lH2yyON9KfSjT5hxdwgXuNQpVAp7by4nIoX6HxviUAJuuMdBXpPDukLFaM4PmWta9k1zgBOf/kmG
ez8TjojqQaV0Q4+lZaZc3cB8CSXCJ2BHiobSjKVF6sRpaf2yF6YfVGxY1jg45h5lPrVHDgpBR1Q/
fynlPMSspUk4tZX8OvaXUhJNpstQwLBx/2EhkENYg47u6i1wpJjcWRpO2vfJW55QvgrZA86sOJSt
36bGjfhrrN4G5Vl+17ftCxHtwf5xmiV6jZfp1gGYm0TNWH4d2UJoHJgKbVNHsDU1DzuobLLUg+8e
MeCfQGkPcPuJ8n97fdmzZz+iAPV3sbuL6l7yzpCaVEYuNt1ICl6S2O0pqDRMF8fRv2t6G8oxhH8D
Esmjx+I/vJjl0Mf01W/imXy+dX6i2I95tKyg+eyokYXHWho/irnGPGgWCFLy+pOerWhTqC1rsZKS
V9oLhKMAVBz7p5/HTBXYjhA4Iiw9hfNPGy0vg933n4jlQ/dx2TN9W6Z97Cy6N5+LMtT+RCru8O19
5mTh1XN0E1Aaw3bp/vTTYdWhPRldj4dfJFm+YS4WB+bmX9rbFkLGUYq5+uKjNhsUA7E3Wc0bxu48
ouFp66tSiS2PKldUTj+Pyt9hhmVBg0PN/tF7va0Z0BfWFpn8D/PYCsVz7y4M36or/ObA7ELQCKSU
krWFMGRsU71igtUYEjrZchlMANYeC/kGRYuMgqhCnV3jRgM0GEGVdAUPU97eNUtWwff6G3ZiwwPI
1jaN9NXWX9lDrFeOSB49Ibaaul8mvsQdTuTkpt5ueqc1NTZUFlgbNjZVmgyl79MPIFHmpsSMCAsE
/e7Bos3wJxtZBIA77lUCM9sMEfdA6VEYlwD1yLvfOVtuXdtD6MvzirFD5XfFZtOemkhPPLUmhdir
qtICZ07XxiHz7/sd479hdLdOhMunRtZhChk/9DTkxGpFY625RYqFJzW+NwSWMO2/7UbFASaDM9Ud
YmMh130NxB3dsJf0TgrGJrDPMYV6VTmnxMMc8tOu/A+hO0Y8NvR46XcEgnrqw4VfW1TfoBQtDF2E
APeLZw6/gYBPOw5JIoPyFJcDjC+2FDVEhtyN91dQLe95A0WWysd2RuENKFVh+FzzZrRY1vF9QYy0
gsBE0l5snawiAYiXrKGPUMJKtMUxGV6RXZ3mi+f8IZ/hWjaMYArokLkaNzm3xb8Jmta2AZfBNDqu
jT1RxYOQQvg13gHBGmzkE/LbzYCGT1rSflWXwxh3aHRUhUMUfH3tE23y/4btr/SDOts5SsGATyAO
InCmmsnKrI2deJm6tFfEH//wmu/cw12DOZhIyAuWOlci9MWyoOcucv4o6penMij7uSOL5VoVxauL
zAjeDQ3DTgMThssc8ACxX6Y9NLUIRQI13pU8XCij6g7+0fZPB6M3M/sktGFd1e7uaD/LLmlRaSD1
lVyrdLCVGhtFo2ph+9t2N9/usGe8jxepVmcqLTVVKLw1XxZ6XfOy3GA9skr+Dyf1cifO5AGFxQv6
MV1lCSwJo3EUjYxP380vXDw9bu+nPw2pXi7HWZKD896GK4K0kEBlOVdubQfn0t20vA9PeO4LWNs0
rGBXOW1Fk4kljmHu2lrr35pzqcEXLwRu+1fvU5cv4EjUpf/nzScHx0jOgpoXtGGGRcUB0EHVwbq8
kX4tQjalK63NpGUDp240ltlHLvOwH2T4YpcFlaHUZfjsKg8gybyPjqpLmia4zzfxBWQLmrEkdA+x
sKloYVwW+DWxwUQYL5zaI07wpjTkmJqaUQWhaXfNqjHsd3Ylrp7cGR3Jdh24aUkt55br54TPwGmS
DA99DRa3pLCNGvjUbHbEqttL6B0BuUj3nxVq9HjNgsck/7aYmhqlxZaKpM3WjJmCbSFdEGmeo3/s
srii5wXxP+3grWlPFX4JSqoca9rM5s6+qTf/LJ84UWd0AYhE50Q2xlPA3E++7sDY/0pkvxAqsbJe
a1oadQ3NQRTvM30zgsnuNnHpBkOw84ZC4tZBqMmK9qsF6Afbv5AFZVsPt7P+lZ6ELUGHpzE78Sit
js1hmTB9vwodnyF7sO1wtel9W6Ag6imPCvI99HiF4autYZyaqGPpQzm2aiv/ApbOB/p9fKahCOcI
/JVgLt4JPglT0NM3P/pYZ10Gzk/DcFyrCcLCwcizsiyk/cWX9qS2jiNivJQ80m106d6b5K+7hcdM
4Fv+jkZjd1V8DgfLeMmfYn1ed1I4XzMuBAcnXQHoWdmE+OOr+vJP0ljuXCSQqwSHghaIMCZLf6G4
4C0NBkxvEwlo3MQJCqCR0PkWFjQik0hk4xZSVqIt80GzRxWVkruOrp2mWCbCXU+iuvjO5r6VUnzD
0J56X8tpW/aUcyXcfZBJBxopk7ZwCL/3YvlHTiUSdpkQ+J1tGkOA3eoUyVV39A7DYH5SKQM6rSc9
0Bz/LzvpUdoA9mk3GoSt81DSAmuKh+PU5nrPIBpPAx8VqG3+e3LlLa/Zrml48dsGRDsy4uzo3orL
Sfg4QrwyrKQBuTtXkXdQrjfzKM76QaWhai63nphjdB5640Lvq0AwiD3YEXX4OJkyJyeaSw8wVum2
gKrZrSRrR+LbOXROhM+gfe75lRT/E1kbprEypJrSpDHnHSdo3V1rUNHOTz9ap/wtO5oCFAceG8CD
Pg1BoeeMTr0ZxaAcsrcSL8vo+N73NpcZltZlTUZBE+LnBii38ItF+QsR66iUena3MbHTslRBw9RJ
VLcMvMd0gk+5D6lccXfBvm7k7AWWff7pddvX0tAgG/6MRKZ1tV2HKjCbh17sGYKT/M6EWCtW0mYl
oHxeWOr1GTSoc0fMdZeYMX/V7ihQ/a6tK6z0eIwEXPre3IkggMrJZXhCz8v6RQKVP61srMlYGGYb
FZdaEXlp07iF5GY1/5/24pgsD1lAnFDS+lBOHfHa3T8ah87JxYuqJZBDGNXUlo7fY/+zK9YKE9FA
XdBb/Lab/MoPJVh1atGkPImozHEu+yKe8ZC//JcMvnUD/1QiTex3AU0YjeDQW8dzcbGwz9MNLicK
hXoYvPwSJDB1PM8YHGwZh4ofceQXgshgwi+xOb+DwEI9sek01psi2oaVlGgSb/NQmStZ9jkWUoMd
gxjnZck3+5egL0Q5MLJFGbN7ikqtr5viOJ37DoV7JQ4+feeUJTYlxQ7yS8X3dDRtMlsjAkodExHs
pNmbxAcYHFaIaFkRiZ2btX9MsZBHt3H7U/6BWFH8x5HfU+7FtEMTNWZmSwN89yCm5Jp/tnHf4ZMt
iRV/KtHPag2hCgu90IjdQ9mZsgC0F1vtfy7ylJEb3KBvpstkrwmtw+glP6SqAv2+keXTZ/cWmn2d
N8d4NAsOsSBzmTHoQJiKyuLi+705DRnuGyM/kmCJhYhZkEirBZJWvNGLdW91/sL77zDm6qmAOh1Q
wPasNspTnodw7KPWe7OK1iVkdLKCw/sUNRT9wzw41rEzfMqa+UeA/XyeiaflafhRpdK2pgNYeU+O
3b/LjbJ2LQK1zHBWcah2oXhxYwLoTfQ83+Bx9MyTFe6hBwjlYIiuE4zsu+fTcubWF0JzUmqcJqmf
5xpWbgfk2HxUJGTwl+HRIZqGwYw8ULj7jPryJsS3L4Ih7mKfuasyA2ChAhy4KRAuGqK4AHzooeLS
3ONJx4vtgjX90BnOyCw4CDQEuEvgX2c7vun3+QFWme23qtgtPPlLRTNJn2GalOqtrxpVPDoKt5WV
jXdDgptKEDO8K0UrlDG1vHUxEsLG6+dEP43JXweVt1/nOownKOMqGnf1dVw6xQU24TAQDiLJ/Gb0
BUm4lluO5CQVUA9QiUotNbC5AK00fOUJRMOBKFFkkKPf0uKmQZW7jiAoW6uel0o7xwzPAuvgyI++
EX1vX0vso5o2VfAs3iiMWp0fsYVjnf/kBxck0+OaPADQZNMyrtmz8Xgu/LiyKRdPG5frw74SY8f6
E4hF0by6wuXGltbDbKzoo2onP7K5O45JWqf5wcz0JEQMcHCeqWXxN0ZXH81RmqT2SNBnDyq8OHey
Db+Pfr9i8k3nAs1vbKfYGp0tp0Vid8CoFeJcOrr4y8ZzAXP1lEGN9v5SNUu1nBZUs48EU1P2KDVN
fbjNc0RxXNZPVE5sIxF3ic3/7PDdX7LFyU5B8UpqnZ3S4zQIZGAb4Xs+wRz1G9EpMgf2YRmdnyc1
6k4ou/53fZDHaboeFCZTCfDU+PC6y7CiYgUUzbwrkeOyRThYzNXV8nD/+JHX7ScaM3Z6QI2LzTRP
oFQenaDQG2T++mzWNGwmSGvJBNSi4x1d+DEMt/5bbJuDXBy+qIGcg6r9EqtqnstvfL6c4korQuMt
6eYmm9IlNCl3wmixnx/iCuzIzI253l2ikNoUNyiJD5Ml9FBcyT72uIB3AONYolVcza+j3x4aOnN1
fCM7Wylt7BKzPSiMtGlIGvOI1skN/HspN30s9G0QoK9rjoL9uS8HUWUQfaztJMCW3WiJNJjj4Iij
Nu7fwntdqTYT7IV/rFFFsU6EYapHBRWMxwl4E3GgEVIptMu8UDvvWNzRU74WHTWD4Y4sz7zQcBkk
gsqN9LG0nmEY6eez7Ww+4nO6v9NoDmqdsTyPgxbIZhWu0qHDkktaySAgI42WuD7A75R0zgGNnQU/
FtgxtDM554dqTKAe/Ikpl2NtyXLqqduoXuWw87dPTRMuv1PdREVs06jZpahtLONSJznhQUjDW1xY
t5hqX3FNVOnLlE0H1a1k9mthubaEPd0gnQchEd12KV2IgCFoqGMttaoVp3CH/jxmjPrs71xR7jMj
fDsgzLZFrj80RtR9pa8sAqcSsuYQ59hmoKiTZN1ViQXhExKm/K6WWKfJfG2UPcfRP5Uh5VRTkdn2
CwmkBkjYavovUORWp7/yS47f9PWEPPuSP1tl2kmUn/DBNMW6OnvRWYdBRTyLBgY+mCk+T3WWRIhq
oYEKfFUby+YsT4ZJsxixRPIkIdYcOn0YsKuK4suK2PrCbNlhSlCknRFVZweIq76OdGjwuZK6qjlA
8a6bH7Nqp3/sFX2Cz4bhHRtCRIG/bkmIxWWmdBISgxPF7HlDRjI9ltNicJMftux+fXpuZYK362/o
EqpMdEI9XT+XPkaHmiYB2lVAUAkW6wjPRzN2Y4t29SSXYsl9yAutA4r3dCFzl9F9tAg07NA+o2hQ
vwd0aiXEQKnyES1CcV1hQAlzSaqFHAgpF8zNxXdwtHfLCDZgO31Tbv8chq1BUGyWyJmA+ICmFhec
3n81p0oZXuMyTTdaMidixGLQ9RHXOOxxtFJbOlUP4gK6Y1yly2yn5Av9h5XpFWsJUEVgzYNIa5s7
raVVwnS8oQRurtKmAkP4WnokR+A44I4cr8fYSqAXxdmC1CuOAv1pebcc+jtLGNFCUoajgxK8SohG
98pAkOEomNnvcUi/6aDNjqrn90j/XUfuwGKp1PMw+ZGvsWISKhX7l1lgMA4yKMzxaY2iFzmhs/xN
GWZJkW5WXzFjlzLtVoTy2IC3zk0WkGT5ZStHQLtjPgiP0YKRdENlWVWwJp0gQ7F5HPrs2mmt8FCI
GzgmKLFjF8BsgVnJphJdMBgmiAr1kCIRg84zsDGDEXlB+54RWKApR8Pe3gBs59tG9l6Ab7YIdMPB
UG9UuXr1vfv9xqaof1Ihfwgytf+PA/r93dglx3IoKEzl6HtoC6ZRwR94jqavmMod2nZe8Xd/W092
izDXFVoZbt7qelyxp7PtoDAcfHE4wpi1eSDA3I1VNdlO+AIYCfG15PEan7bhhkNcRNxZ1vThzeWS
BA6G+P6+f4C9zppnDoGfipkw6v3ktW3wj7GWD98DG+j75yeb3cBil5IuKjmFVN9P++CTfg8CUsQT
Kp090Bz6ngoosA5sKeupgmCytbMG96SmcL6wzq7pF5hImmr4+tSIJIWGPxTlu6tJ3fNXPXW4bLv9
Knhxg6F1MqEa28s9GsoXRmtkHYcLHDqB6x7s7LW2/Vxd8D9SMX2Puzorovz1NhWHjMelR+NoBQvG
pmp/gVRLzlLIcmlhvZZtcKqTBs5TolTqUy9APnV9rZLv2iqWUfVRQRoKol1H3BKd/GfqPPs5jrCZ
SYqoOEV9TEQxUH4jc7rhdJJRCekKwtc3D9Gsmct6QC5hKCiQ4Qx9MCbBFcWTSW09ZceuWz9w7Wl4
vZk8yLco1K2J0b95jz04/jyjwl8lgJzB8Yn8ZC0UGD7TT1pTu8mKCy+gUClVECAd0g4xswldIgm+
FjuEamZwDrUbDKX3huBBek6CoMS7Bf5gmMtI2dbs3jtTB5fG1PSJY+MbefDyE5jA5iKy0gmILRmf
+VrDDIEuCHOyJEsOZKF1g/4Nxnx7WHdm9NDxFFyCgwylBgexEXGfhCuR21VlcUQglOICT+TBtVzw
LkivR5tvN47yHVeXDNE9RsB9MROidSGrIEGst7jqwqC4i7i96k4+spBPRGMl8e3hV2iWuAqU5TAV
i7v5yquhTw0OpLCQz7LxUEgi1RHM/aDDyJC68Xyd3GEqJ7eOT5JLtGRuqkeAGe5NOT6KLbsFfuXT
RVGazr0t58iQHMdBXYgj+Huk1NeNS8Pk6ITnsPmkiPipOJk6Bs1lhOoNzjD7U12IFcN3Le0Od7yk
4C23dVmyK3fqUzvknpnGQF6DoyuGV81zY/43Y7JZgt7I2T/eiJl+K0Zuy2zMYOjWZciR+DImMTAI
2fKH7qygxo2KC00Qbu4WcDyCUpY/XXYPSH5S80bCfSAQbxEu9X/pgeKo3LUPZdF5vWvpMUWgMhHC
nXzAuZepEv8tFSEC7LHm3qyXN6TEMt+Fyp/4mxlzJBPUCvpoq2Q9Rt6lyM8iCU3SHyGujN7N4rrn
yCeUfdt0W9tgwHVQ9lU0Ea/lMrYAafk/JyBcnaYIbTA30nk4GPIaE7Lj3Ai1QPXU701qOF4uNmio
cFrmV65ihQfCxYlgaB2CSO1U5q8Q8nMWvQsAX5hGbLVQjQJ+GBmAbeFd+OUWqHHkQ+3w6TTd+Te0
qn5paRzt1pWSPEePna5KPBmE69SmtvYAT+96jKJKfGncZlU5KAQOcD+sMVHTKYFoLfVTVh6zVOZ9
v/4v7Tf0He5cLGyyNdX5OJyb+xJn5YYe+GsJ3I6PTMxse1iIudyhgLvMnnQDgmhSS+SkeUQLr5EU
wLUjlqojE1xsn0+QA+M0ndhvEH5fER78Gcw1dty2InPQ7iZ0rt5orZNpoxQFhAd/PVxcc3XgFyeh
HmxG3lQquxHc6NJY1eh+U+shqR3eHFKBPLR/7Eujzc8t+8V8ycziABoxwLeDUKKHWO1D7ZbCwsXG
uST/uggjelU4GacH6B+DHETvetusxAQ56WnBMRz6fmLxy3iTjcsVkPa3fiS9lSGD4zpRR3fkxpgC
CGG4EhbB87+1ZwuBoH0XQrSpXSwjGllj7N9E1jHIi8TGUkqWiCzFGeWUbDy7gYre0JMBbVfMB5Ha
wsFQfwtJjgEBReMToZip9ipP49jKc8Cg6RZhHOl5qVfWDc7OQrDOxDhKlZ75DBik4pqOhBU5RbBb
TmgoZOF31q5QAe7MZUf+xh8dakwD0IZhBXdrH6EMcdEcwmPqKcWmoEP8F2yXRz5W4GW1EILadxT0
hVclTrQVmkPxUwtS3StPMzsqyJtmcLbJvfJtj6sYC61LGKXOg6+vaMjlQsZYVz8iCm/RAQLMrSvG
V+pwMst4FXCh0ZLyc6U50i8xg/UBWomrPo8q3D5NoKWr2xCz2v/LSgmpxxBFLslGKsLwn2rQWncD
DpEhR+TAC+53f26tT+z9NQ0WCyuTHe8ilepi9DBamijz5KXmVJbVBkn3f+uRaYKW7aAAMBEh+w7O
rRIF6ekBR4ZGNL3x6BL2pZLMDsZ+aIJpMDhSUYkijmyrMLBwyODd9lyRPXXiRbYOFUqsBf8rHV4n
a3ySq/MU8LTacdO9qit0SGfnJWol1zzc/oJDjety/2n2ddrHwU9upFwjZ59jPiZqCkjnqxH6OBKV
IYMN09Q8tixvl6i0CiiIMoNoR4DqbX78LvEXXdSYlKgYvfmp6evTJXS/ApRHapplD3y8F8xnalu5
WyVPZMfOt7oljd4j85VmU8P7LBwFuUsFGnmuAGhCD907nacXMT+IA0prg26VW4cIt1KnJexh7sox
4VQy1t0wMsWivY3izr7E0bKYbdi3szlGrBlWPl5xVhEKuJlFr0GTKR5qpjfH6IOK3Gua3x48L8IK
5sQWOK5dmXYrhjMQTRh6Y2uFRUZMDc8PiFHtxB+HAxDLytrCEvC9E7UhJ/rKXB9nIkd+qsaAdijd
Qz1kAHpHQBo39Htqs7b9jUmq3shvjAQEU2cB7994rTqquacxzf52dBBzh6RSZRbZmyMwcDegD0vE
elchTehkceIVHHrEq/ywXS6liWni/n3oHQ5ky2QGmPne9zgktnHJG7f1pyhRcI6abCgvDfAyHdhK
6iOBjoB2VG3gKvtn6GK4uXMqurXQ9SHCm1UIcXXrJI6Y8RC8PMTfCq7bPzaEjMm8V4cFIEkefbeU
cHyrgiionV3hUxLyajyNAxzsNZd5Z6qFQNJBoQGhxKHUwA1gMPhNlDDy9mEdsmoK8JQZ79PN7/bT
OQcVnBtB34f09oWaszl7rYkCRWV92eBvNum3CBSSIV0myejBrunMVbkojtaVi8avh6PGJVMjnXKD
gpbES2pdRGYEipqYHk//t8p9ngqPxhIOpj6XAnt4xCOGJKmIm8GRLUggIGk/ArNSnZXm3dXvrYLN
nGkBw98wE30p1iui+Em6avdGj12MGLEittdAzxiVGOmX/4u7HfOKNImWm1M8C/8oiDGY+ywyY75Y
G0KgMHTkdl5bxOMAGHdncGeU3QfFY26fPbOU+y4T9XFrc8Lj7jTd+d/LqwL6Zg1s5EiHhn0J3X1f
C+7/thuCiEbessLcFAsRztyIbC04saYp2CDyC3s4fW6Efq5Ozi90ryOVvp7P4ETjp1IrD/JFoFrm
ZHVftpm6qqPIBgr4H7klK2Uh9UQ+qOjHVQkXA8v+hdkR6LxAl1z5h6IeX6nwCXn6IiZwq5x/bzSo
VzNcuZnUY/W4Z/1GGH2hjT/tOIBjbgXEEDWPj6dUSK1JVXU29p8IwCvpm+caCLDLgZkqRUZillBA
D50DKZVDA3yDhtQdo8KAnMYrkCttqN6CNHpnjjonK4q8PgKQdjCPGdAYlaHxBi3Ft8+gvjuhtP66
++KoUdozTja4RLUeRugJBKvhyGH9QGX+bkGhf+HWIue3io0r0pp43baG2ojqKbaSg6DpbAQCfhev
vu2tRamZL1em71gDPTPu0VtbXB61HW1qDNMujmoJgGXK7yAgY0DuKR2iZdAjLb3cJtpWWy8EEDAB
9uGzUgLocPFm8T2sfygvznajAwWplFA9Mul42y4OUIsTlpUndimG5csibeLzQTfklpMQ73fWOe99
N68KGvVdpAE8WRSGbGIJVG341wp2dBGbkYpJtIIrLE+uCBrN4gnoxuqpdOe/gLbu3JKfwWeAsXZN
uuoRDeUNzr24mMt4lvDEh0KqXJ9BshB8We5RKNpAvmLWFLOntP26zQKSlpm2fK2mgUI5CljNk23d
Z4TfEb5Jsnd0MXDgyqz4pBjGBQqQJjSAghq55Fu2DwwiEP+u1BlCKgdvYyFi0jVnew6lKWZEZiul
QNGnwLUWTr9e9SOj4/+ofqSwoh4/qnJoHET9mJbgtBb/+RawHWlzP6sSxSW/6QvB2SfBE1/PmylF
htkIQDPZs6455iyTe0yiEC0J33itHXJj1hBwibKBIG1SwdmVBAybteWEJqGwix9qcGzmyoQBosLM
EAxNLAdKHC78cvGqNTVUAOQ0vCByAVf0OEn7oSLdPUSrmQheCCvGfnHu9GflQIHeTRnFtMVEWj1j
aEeYdIKuoPUQiU7/3whMU51uRq/XVJ6Z2423Mn9wtjNfBVnJPI6aEfG6chs8HzhCDh0Dog6FNKIw
2Z5CJHr+A+i5b4nXv7rn4LyHmxTFrsTGFzjhCfpBoGiKhuUBRWIWfMBppFlZNKPjc6z71PBwJVej
T+Y0WavWGdFA74jEjoxgyz21SIRDJ+eJ1XN0DTxc9+0gefJlF9XbSFEw6dTVZV2Q2ZQ//TVoYk/+
StD4qwHKB0bS5iQSKEk8WzRl3kg/BfRDuCWNVCOQVeKtXMDVNjMT1QaTVfl9/3Fa98AuIK655aSB
jUK8wtRNzGeayCVMROkpeP/P9NiC/Fg4DMfjVtQqYUqboW8qyEKm/6nMthVZFzbSj0G687HQNKA1
WyvGRbFW88cBc/jaf7FLqZdCIX1jdvIaPG4OY6bUajo6+hzgyDcNC89/GNSF0pN5JGNdPjM6INEX
ePOOzMWdmRwt2eYqqmH/+DrHwcLbh0AbCLN/Z0avr2Ct0S3tAvoEsGgl1qE47lKQffNkKcypFNIM
vOin3T9SHXL5HkFPqE9U485s7k/xTOJr8bzTeGwKJwy+eOuFPR1BP3PIDCU6G/RF9U5freenyjY8
jBM3xkq6j2hoi+QAuKRXLXa7i/e/AJFIqE5mAR8x5SWoawcLRYF6f2bOOixloOMoVrPa8avWZuha
XAXmLBXtln1YftC6pRPvjQM5MSvrblOlfDYh69b4wNAX1blSaGOPaYeIkQhcQU6P82k6cC8rn572
qZt9sL9kQ9UTLMBhXmzQjiZZ6xUPLJ8WtYZJoECoBCeBLqdclCi+ddxi2Mio7zp4av4XyLNESk4X
JjinxJHqe+BU1nlKs4J9P0wCPp643ov6bpw8s24pm6YKex6n8Uc4c6HVlqo+j+Yt/wOiK53WLwEo
tMZ8KomNTVmeJG4Vl8IqaU0OsodBINRYvLbrijcV8+ySCIW3xnktF9SJk0GNJ8nlCgiWddxad/dw
t6IWkdCHYFGao4x/bFSN2QCwR3juvgVrFIhS2JskfXfIxHgU/iY/fWckG/c0GKSdb7SHY0rmA3zw
0CDbG1zsYjZRe/2ktO2i/KMj2Oe0wN9OYCF52ck3s4JFh1pyP2gT52IWq67hFjSzGyCJo4fxV9/w
ISTY3a1jMBq3kKqHHRCuBNllAh7EADFmJ1MAgAeDLvpatAnuqCdXzYkFTnFBTfWFQjjAkMkrIXpa
03JU/WRmRNTeb/PJrAm7+PumHf5wSgXPZd041adb4nBVz4x6PJhbr2VJ0nxSDt72ZJqXKpBACJhS
lGVY1kX54KsuZ8pQBv5oWIWkO/2AYpUbzbXfzgCJvGj5npcvn0P4X51fy8r+//Yl2JLj3ynIAeMk
NN1aRFiXdOO3wdEhtfIs/MGL46a6diTt77UJ+n2UeMv/hGU4JlI1qXuRTxktyg2Usq2OYrf4tRbQ
2dkdznuTpRHKFSz/PukO3KHrzVU/Ng3Yu9eK5zlPmzeekRaJ+3vThIw5K5q9hByogjY2cPoSUQtF
Q3MyDyT6edc5K8d8ULcrvNpzZxD/Y7n691FO0YNIEoT+ZCyLCQbx+q9VeDvlg+v9BcWzJ9Ixd2ZR
akQZmd+gnV/BhtWVpFlpXF+TAop14S35+mcoUqGMoVG/AawMVE7f4j+dp6qFXowgRkbonJJ4tpNK
v5CG6RA7+iKuOaKg4SyZuuHC1LMCoQQYBL0hORU+BFbL57MRMg6zKld/fHW+JSaasCqkT1AqlesQ
3tzaH5FaeKDME2RHtTzwZhlIEhhmQLqbM73KfacXy6XMLbrbKzpOVs6t9gZUkIRsdSAO6IanHM/o
OQu35hB5P3iQdBgVmno6MzKJv6a3+IUnGAcBtqPhCPf4qu/ZYGrGWt5lmY7vsnaMKoqhuI8zl0Do
jlsKQbQ45cVUGyJRyos6DwD9ilySckfDGugYTqNyJ6QvfT99gQM5m+hrKPVwH9/GYQJLR/5U4PiP
ZoeMpSH6pEQ+d1P2FL3cq+rEgrRlWntBib9PIItBFbq0JGUS12K0Lqv7GHr24KPp0ef5nvsyQFWm
RQBmTGgq4r/ff0EsJLzEdzn7O3rgJeFOW5cdd8hsiMHfQ5+qXdHEhBC/GFBPUADZSJ+3L6wtfnAC
12Z33NSvzxbCcMsTXd+wgLfU9obQ7vt96QMJWYddj0OyBBdFa2Xh556N58LmJ3oozzU37URJu6MN
QGN3Uy835IYzT5lXOQ8IfAT4vbta1GYhaa3aDbkJdSuZACYu40KYVfxfLR8EfvW+4m1cT147gqTt
uRKM+RfgfyCpWdBIb3HTFUti+JuwOtur5tpoyiY+bvRmKi7Ov0lCVbfJ7US/Zo3phENMIdCl4/UB
WLL+iFpiJg2lo7k2oXzgvF3qbdLj9gob+//9ZRLNU0AmXS9Mx3WKeMCjG870uVAflW5NZ8UOXnTD
dRJC2txV+kLhzjMlIEa5YTbbj4XDrHsyydB8jsXt9/RZNqcd/r1G6dr2WficcGpYzIhVG/pmCikz
VhljWFndS1d5hMVG4LUEa5pVZQ7P/7u17pvQ5tMI0XXf15z6IE+9aVI8E1a5u9mvpUMpfTxBMznt
JwO0g+TVjyfMb5TjxBJzgkHAvXIUOkb54yWMrXTAj5Tw00TSIUf5zwvrPmbO9KE8Qx43cZTvsQ/k
/Gsqf90eFkyElf7TtIMqpKK/P8Qx599HcPuVfBk9qFnU8DpGGBEaViwPbxyGmJCzSX3jtlbTTGBW
+scGez4Xc2nZkEG10n34Wcwo1LaB37X3xg4GmehZbDXt04+nVHicTZeEOBk+379hggrlZyz398G5
7eQ1cmu+IFBehpFkMpvx0iAp8IbZqQuwE5oG6EkaPo1tdXMMcq5fQ7XK07nVMf0jhy3DwMbqdeXF
MuuqHMaKJcdC3FfFMKxvFRx6Ufn7P8MQaEYJaswek8QPl0u4/Mriyj/XvcRRygncRZbHtB0Qg/x/
Ev5P7BC+xVri/I2Tz5cVoaRCNSFMAGNeAxk+ivQ9PKZj2ok5X9LIt7ueM0kikBQzjxzQMtqn2AzB
7hcHHFRYV6WNLF0ajPFsFUkqbuaq+3pn2dq8TcbKniUkVK0G1P/pITEIaz09rz3yFgknil4iKYWO
QUHxc3X+IoM/AogwKbAvDqcXK2/Ka7D1IOIPlGNTzL6zmK4dx5nlH/ayH7v3f3NEZFGlHxyZ2MlC
BT0hlE5SmHEYA0O2fOM9f/v25y1rP/zbVNMTH88ZEsAZSmNwsG2c4uIERIS218UUzS1tPpIddvkN
TO2qWBEECslE6jXi0Z36GMkYLwEtishRWTMc8GsFLpAlP5/kvT9P8BCjURcgBCPFYNPVi5DGtJW5
o6Elj8twdCbPAbVzcCalbIbRU8oba+S15od6b0H+Ta1LGKGGkCoWTOdVk89lB1x1brN7YQ262xy1
h2hp3AR3JrR5l4bg0RawHFk0swYo1kp9DyI3s8gTIji3A/EwA621WHDy2PhN1Ecsmi1w58mu4JDL
PrM6Z15YpQlPsXKw4dZdHbjY4W5AFwikKzIZLRCsLDoANOZu04TN3aa8QBvIUEpRXpdLNLre1bqN
pLzpV4qZZYLCgb+CjBGsO98fW38Ka/XtelN/9qz+eVOcyPj+dLOtq7i5zFXP7ariH1fvrxGcud+C
rwLgzxZgStt2mWDMzu7utqOxJHphCLsfdr2E/A6AOeWQAKExypXdd8+aJasOb38fPLaRCfkbZ63i
baAyk+5+W+tYG4A0ni9p6WDO2yxEasSf8l09UvDcfU/gmwQWfnbsHrTYXimRIBTuVOsAARhC+n39
00DeaNUNb04yFhsHM7q/EQ2Jsbc+3S1beUS2mH9FDUV+OBI0p2OTXba3jR+B1venREdztjMquQgn
7oIhKdS5R0GQ+/7OHDjAsa/dSc9e8H5tu/3C8kvVFeDJQ3/59NGSXMwHhc6F85ibxgVblU71Oqdw
XzQIucR7QygR4o5w8oHPfGGIbcMsJJn8cNfQ5NSMCWDjltY3rG1VT07+ts+l2K77edqRGrX++zZ4
QU1NStyPNl4ooPkqA3jTxWzoZf2MSCg9AaYb9+58ScELEMnRl3KC1lZK8bQo7CI4FlAZVBqgZQDp
A9IoZuPWZKcU+giOhYY/2xDVGMZWMyb1loFFgwiF9xRIuGVTbMyIFxqXGtxHuGTdYem/IUWZxiAN
jKb1AaXEXo3knk+QW9W2a+xRxRV1vLjSZIIggNTjbCC3cl4gkx8O8ygjJIj70RNSFKwy/N06jJC1
z1NFvUhwr9zQ4KaOKr0uHtBvor9pISN4DQWa49D/rSvxQ/crsygviiS7b50YED/X3lDoLwJFhmHU
ELsrCLOlMJlKr0ps7G1lvcGGgX5dcy6bPG9wGWoe3odAlLZQbbrk/ZkL+iyMtoX1q0odFohIwnG4
3+/TMR1Z2I+7PRaCR6G3M3skZpB29Gy8Nm5OnSYh0+apZ4zoRjgbjVKuCwVoIyhV51EapXaE5mrf
2+ZLnFKzLx2JMOarTKWOC0F00yvhTjf8KThyFSug0uAwjGlJTlUg7Y9J5SkTvQ9sXWNCpXpXlZLt
DsqU8vZ5y5H7z0R01CbvBNPXiowm8yLRxQerRzQTe8Vq9MBmSC1ql8fSoKsRKgFdd31axdYul7+v
oPUhOe6Uya9DjFjLSIn4vbTrIq5ENxgYU+Uvxb8iu/6mP9DhDoZU9Y0Vkhtql3mOLv7ibaPWrGF8
jaYdEnUtI5Y5pkk4rPgZf6ejfJX9SOSIGHcp5WxgMyscg9Qg3aSMlJeOH5J6l2gXR9pcSg1bZ5Xk
69T4Y7sCB4pwjq02EZVqt9U+9FCqk+AmfOr7xnc9k7LfYXySt99AjjwvydnHBT2RnGssQEqeV3u7
O7dyX2xdX3abobVeDhUq2QgrzN9vnw9BkgnmwQ5Q5dsJ+ajQterD20JEgdoRvc6KZJ35FChmhLMG
hIK3EPvAWnjwXf7sUjO5o+n+uwadgYuCkxxav+q7S14d7cJgX3Rcte7kGO5HL9L1GLvNer256mDT
MDV5S/WczUMWfZZYC8I9fh6hmv8nZ5j37CZQFa+6gsD3xkqSuak/xGiMPfoNq0q6bHkwoU6rNU4t
497SBhRWSMD/ewtgdmkgXT9MpMEBemlROZ5fKyKaVU47/bEI9ZZPwJwZIkuVqxoBi+YQx6S88XP2
WZbJA2rqXafF/lF+pnPFWjH7IKiYsFrp6mKzny6Uz7afo01rYXOJPwWgnaKmNlQUllaovjdNLULE
MZEa9gYp0w+OcUR3xKGtZ16KT6KtLYO1klkIla0A5ABTyYCYD7tEVXLtDjnpySTuoovcYZWG1xMh
O9/tt+G9AEXddDTVsfsUFTQIZnd6GHqVI9+R1ooKvs8zeMNoo1Y+Vl/vUJaehXmfl7WHDvFXD3GA
pKROYklcQGDN9+9s0MQZaVJyj6IiukB+6kKx4mRFt1zRVhcfIsvxDJk0WPUBNB6+mzx0ewEUcvus
LbvLT+WeVtNlZJUbdf9wbPmvt6a+HFP1UP51qnWSGC0h8tCiFusSIF9ZvnLpHLaE/6omRQ1D2KrW
eQawV7xocZKdeHKb2Zv4u26YABnAllQRZcm57wnOt89FY7BSrPCy0Wnff/v+Jjn5vQrXeNxFhf6+
QEE7mRoL3HSdl8HlSouPMffkXmIKlcWtGsinwaMzDALLVcBkUjZl/EIOolRTWtAumOhRN3Y+DmvN
sr9LuANQIZ6ww7miJ7kfD8vupYAvMM4kZLaDku+x67MlZGflkj42wKBOZCBIIEsIN2AvyJ2ifCBy
XWp8zQBcjVN6LLMDv3VyPc3zKPiXm5RZREQvzkGELRufDNRQW8pM2iY5ppVINatKt0twd7Auej1Q
ehDyU2ItO11gQDzFTyimWTzhNk+KJMYzhI/m7ryWpTeTHI5J03R7l7SyxMbkp2f73v+XbvlNpdAV
/erYIHC80jmv96AU59eihavIBkU4uLIy4/bqPfOVEruo6MqoC4sWj1NvsGCjDF+XieRVU1EW0V83
KLToegCRZP3xtq9VbI5YQSjv1DfBRlNmBB/q94t6CwPM1OYA+Ip/6B0g0a1uyMRmJKVuRJ1V+IMp
bvEwviVYnL5bVueNf3n6ymcEN3vVq3E6t/sFyos6wZzTOrozxnYEUFfqTfxAbLK0HulRh0fIgEW7
MBkJeM2SfL6QrTsKBLtz+XOjjN97nYsT7U2WtPnZDppXY4RGMrx/8Nmy888g8LDqdZ9UUIFPuYca
c/QoY1rarmqLwuTiSyLRMeSob3NMZyxXsQz7ysJ1MgtGgMkDepOwdOjZ7V2VbgJoTRFNmRv9TUrR
Ij5c1mp//13fevYy5NleItjlGayYqudgq7WzuwX4inMPK9uWEjmP59X+A88/Oa9IFe5wr96rFfLb
QCfeQz5fuqf4QL5Ep2HqLTT0EbVfHfQxuqqp/6SXj0+oEJGC3mtHwGVS3UBqI+Rdb0F3mtLoazO+
ZfsxotjYcAFCtG6K7KDsbGvDcqDX13xgTLt0EebxXyDBweIt7axfVwuVhV+CDLcOlO939V6uNNXA
sHewyKifvQ9hl0YCxTxApJmhXN5mDSsxGfgizYxbxqLGV8j28a/IgljFWvfs/kYbql/e4LQNPYkz
/vyiSzOzgK4BM8nK9MGIA4jlPLxVOAuB2xGC6lUXtePfJu2QfIv3sDs/rYRP7OCb08NAwjnHZ0Nw
NeSiV+cYnYwW84Iwqf1ltum1fpLHVHkD7Kh9LbKPjPDAn7IMts/PZFjdULe/C961KfYDnmrScXIw
eQ3TbxTM6XIbCXBlkKcUkIYFNflFn6ZhaTKzJ1qWNxtxNX/DuTN1eMDu70tHmgICyFEVz6UUQ4Yv
HjUm4Zy+Mw+13/EYC+EcuCf5jz5+Zs6HTYvrjfks2FZ+BM/EL+GJkIGdolklDMKFaEdnTq2N+ajj
GBWGOs2c0D24Eb+WKpfdkzENagfCIeXfnCDj7Sa7Ow7tceu7k9D52Ds809Hi/SqGB/SDFdEIa9GY
JQtwFk2TglbopKa40E3WyNFgY8F5LW2AGxcctY97Nve3T1qkIrZhaBIU+krnNz5V0+nz2bAANeLK
B+yw1ZJmb9IEFISDzAG03etSYUth3ycO8HujADhbU79xmITujOC4r2WwhMzP6OvTfFDi8jlOmcQ/
VnizEhS9z/E3gdTO9Nb9XkmaJMvlOQqFaig3vRCuUEUoHorTzJzRlmwqlo67hyAfKerps26lMiH0
4LlUFzXMi5HfMFS804Tt0rMdY5bnfWMC/LHIrxkyH7OU9TMgf6JRfSk68A82g0970Z8Of+V7mSaO
DqnQBX+2tCcO/3v9jUVOegZ2YRICboR/LBHtGE+B5nZo51yE0KoL/5k3pvEJMwVZbKgzSCUgvNcy
rCIXskVQ2cZXtXr8toOQ4VYaEbmrTHi2mlMElFkO8TKR6i4pkih0FRg+bCbopi1DVI2t7C3/IBjj
qj1aogfawynWSkCM6rp+fEmolFVbZyrVVkEpQ1C4anU3U3CSen3mtlMwPgCB8XRtzROgKFNX8U0n
V2lM7crnAXcQOWOlN6CKGv4Tnw+bhT4f9nh6QkcZbP4DSGGLlsmiEktF7yjhmdG0jKjQzW9xyEGW
w9TS1A/Rkil/ID49SIK8RPfZA+WV87gclw3kpm6RE2Nzr7co1id9cjb7Vj0itBFP8G3lz3NB+eaS
wMwHf9Nkp/UqoYavrhbUIjckXU42smdjWro2WK4st3fBfaR75lbBbD32zOAMrra6McIRX58sifie
FmnVqLymTxE2W30pnppp5GlvCcVlF2X2MSirD5GLjy5d058qiO9v0tLSnk8URhmZvWfybtw9IsLS
2j7Ns4jsYaorZl5fPHCrOt0BHHY9BDx1xy6VcuCnt95N7lRWcpFkpRQJ31DkRSosMLDNNsBQj+Ba
USNx99X4KYejjQQ611y0IP5fdFUvkpvYyN+hKHw9BKqA5lv6ZeMUjgJ9EwSp9V5vqmTMAqm/Kdj5
Zs51Cyg5MbSyU5eQC5uzYRS4wwgh0cXum9aJdasqLxYjKr8fH53XZtg4MCqybJ2bVRsQUaRbWKAI
nsoC8W4YRgWDcOh5bLGOOZzAE/rTGgip9+iqrG54YunW/0sN+aTef8DfoqmJ3IWG6V3iihtgoGrB
tGVCVcH+xoiRk/8Oku63Mw5jacr5GanfRjudUPEhZn0K7pxat2Io1XOApjIFfNBRWE+0y04V4xMk
GZ0qCv9LKJF6RXwLA0tpOkzbBjZ3X0utr15eEUadXgg0QO7QR9l/Nj3RF4mEf0dQo0tw4O4i5InZ
JEjdchTJrKrsQlFxTHDUdN8X+A2rzrkx9xcD7HwP1pvazHf3tsxz/Kh1cEx6/QcBDtlpeG2Oiv8O
usjEP+bVVeB//l1Li2mbHFMSbKrqyoA5JvIAxj52AE7NKqLPdv3zWYSWvl4aKKAJlNYf9JVpsKac
k2hRUm0yTDlSc01AAW0crvHlH4ehDZK+KT+qXQX61Wi0Wtlg1+0Lax2uzDrmxYIlo/MdnnybH9VV
tTZQLDu9Z2UhUvwu+wN5z/EofF3U19qLqpSBn5GbycHV48gLRFFuxLUmChLPVNbAVDvmbUFmPQeS
+qmdLzST9ZV+FO7MPRi29P8lfrZFcig5SHk8WV2axQzQqLFd5UkKiL45Q2AUCKtbN95e6i+8YQwb
ewmIpKP8bIhKLrBYCeh6SWuaVjpSAFidG0PRi6rfdgs4fQO5yI8fyhgjWmCIZh6bDX7i/Tw0Fwdz
CODa0ILP8F6scEhSQ6mrvcr3RsrNc4E6I2fD8sVZ5qMvKqVScQGYiuIMvp/jrzAxvvcPbE1cYqas
5tYY/yCpb8XlGfZu6FXx8Nzt6pjwmoOiWLPwlPVgw2gQ59rIX+usT2xLWXGsDV+W4xZYN+bqGU81
kh1pDVLTeDZ+CJs6EHOZm3/4fPQZ09SVKPY9Geljs1Q8Pdz6RHdzwaN/e5AMU57s1PY=
`pragma protect end_protected
