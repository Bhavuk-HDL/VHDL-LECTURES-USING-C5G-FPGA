// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:21:34 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
C/EBxh/9XOqFOMU0GgYZ5CH/ynk9exdc3JFlCBw44fsMBmcXYQ6hLmFi9zxl7C1f
VcjsNT91zfiwnjUvqBLNFcL/glt/74cH8al7DSnYPG92d9MGjtUq9NlIqncmYqmg
2G/nugqUxdo9OBMyiQNTH3n5xDb3whbptFE7fsT1ViI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
OuH5MMms7WREjGW6nY3/M0I5hJitfgLnZ9Ybm+oE0vOstaujHKgkmHeSjvHcjZkJ
/VR5joR2Pc0Ypa7g/EhZf1FWUactpixQL1zLIx9hXCRQCeWShw23pey7d3YSK9F/
lkyYPz7oq//kAH68wU2eMBu4DPZ3DckWgTGxSLwQKzBLw+YPpW7SIJci5G7nHcYM
sLEkHR4JnJAptbexnXLj2Xy1LkDsGXX3+C7z6/e+t4ReUd2kc1IpOa8TpXTemFEk
/dsNcXpvxLKn2dOxs55gYX6wB+LYseIEaq41o2FK4V7Fo592Bf7ilKTaOPVqIj4s
7/PAncgglY2bHDT6/gGN5bVPq77pNCOLs2N4zh9bP2PF9zORAroH15vmxoSQ30b8
LxAex+NFDOrANn2wTErf6AOavRdZqhZxWE6C2xgI2ihSV6rJKF1DkILJFPPcWgxY
LQIRfLWpOTPhruO6BpWiTh+3t3VzpX3Zwp5PHonlY9Ju/an1OWKaEad0JfqEJ082
URCwjJ99QKdeCaBU4oqNJlu3P+0dlTkRPORS4yq6WCXoHQHN/TQSDJf2Rks9Mn8U
bUKbpZjwdRjGlhahPyBHye11KkenVMR9oUFMwA9bI76Mmq3CtuBUK0jaLDRsRnM6
OGsLf13uzKCjxIaHcRp6Q1qOsC6/jbyNB/c0OtimfFKGTTHnWi9m10dkmGZ+pGg/
Y09vG6p/whlcr6JN+xV9EmWugUOocuaC3waPR+WaGbT2g2PU9SKFZw41wxouzD/8
f2Gs5ANUDBetJxH1SHzGRzGqXp5k8ibe7KgZwWRBKiAuPJTw088VaCThaDNshuIz
SG09eX3zuOOmBk04bDtVh0vGJvCPeXtA520J3bfV85SF7Z9fFBZUhLGlpXzwd3ax
ojyQ6eMkqyFDYNAeNeraGrPBQbcuI8bTrHPiflE+ApcE701BCHXDgPsuHz8pV8sH
IqOtfFDpk4Qnl5zJdR5Xz3vgasuNFgPLXnJV8Br5XuQR+b/ZMH9FeMBF4tyrgbda
laaRPrHa5jeLvq+GaPBoLJOvEoH3c8J94QHLN+pBJ3kgiq40bc5dUwIJj3Ll0lTw
gkfpV/5Id97YrVFXJwDQLNiLKIVo0wO9ivLbj2IFKNt1hB44fTAqYhW6+Drf/L8U
EQxg/VBhlQZ43NCFZJUZLE1HMbqzy6BXzgQtL3RF95pDQ2LJ0+ikuphRCzVp2n5x
Ch8AIEEPo93QjGB0oW1H8GIqbn1PqtuoiaSdSd9VKO5Q1Oxxb0hfGJd7T+AK4+TL
8apJHKw3rn+Vtnd8hzr9DYH72clKag+W90EIN1xdRPU+mJD8WF7Y1M5nHtTzPtgI
zVVdasfw5i0GMnzIJTN5OFfAWA/gnFKekkjZan9jvsGflx/1appBKTl/vsqfMIZY
OJ6nX/NdDGKvNfRhFCvc4g1J6fMPNRnauXqZtcGVu30kBg8mMQiBoQGQE96w8NBy
sZHgXGNUwTuLL6oOkQDTyihwr1fcRAS6MD+xgauhAdmiddGBhQwsx4xkByFwFfoW
oHq2/eElRMqSw+4gvU4sCj//kalSmdm1BQOq9+hiEnX0NdZ6bnMm3pCIEQszMHez
us1s/BvXBWQBlmYw8rV7JD14VUFGT12R54YryzPe+rEMGEWezQ9ZEQiYO2woHCbr
3HetpsVFzdZjR4EafW/xU11vceBSiZSjws59qmBOzEtRh571ZE0SxDyBGWdkbhRW
Fm5yQ6S/ws5E1z2lZoTHLAPZbEMKs3CCrZy2CmwpHD4ssPAAu2IxJW7WmW7lIwX5
6hnxI0cMzE3oiWTAUYWAiJoQ/8Gx7vs7EhH3dioTKQDbKJ6hVuM0X6cRZVInEr4v
99jxRqNpo9255kC7FY3Iehw3ZMRkVfMb8SFXfjMfbJQub0PzTPmHSXnzqNchFgpI
8tJPPG8zc95yX4HdN7icFmKpGUpWGisvkzJhOfkpmukH71GqaneQOZZmTgvn85+C
egcpuHNv1ITuxqi/QjE9pYgVQGK8ftSYZFrfxj0HEZZBdV3dV8nwVsBf7V1pRbfk
M0LbOiSD+MHE67hOkc4mYVMvAxp64Wt2Tp+JS0A3Q+EWytUhhs6Y4efSgFDDDtQs
+AY3Swl6lBXm2J5LHqpBut35h/nAOKOq8xeTpNTF33bH3vNEvHJpLVPwlYVrc8xW
6XjXpqtB83qBIQV6w7i6yo0DSOnvYaJKHTZqyTzatittZ0Wts4KZNbNUt7IOP0My
wPBFgsIuVm14OhDngQzg7EjRgAsHYFPVYeCAOjSllM+7h4qAukVB3Yd7ux6ylTJO
k9+r4TBJOwL/sHvae5x/NtQF2u8uHLF+9ElLj+MRCBbH6CnBorpCjETtCl7VXFw0
H0u3OJ4oD+cAXQimGZ8hh64yxB75DN8LZ0fpVmaM3+VeikfYWAIgeRfP0SLJyFEW
kMwosh/+iXrT6GJwvq1u0SJvry9CWH6rI78ZxPXQ7OIp/Jr1bwc5GbshOW9AHoMN
rIlJ0aZQGCAEa3Qd1k+acD30cvIdRquFdyI94pS7O8vQxJMvGJxnQkGM8LoWXewG
aIEseePMwLu3fbjhfQS4iXApHV1BNeQm4uArPSxF3sgB58iDtvQarzQRx6OsNJBS
RCqP8yS7e5wppF/LC6OedmDuLddCi+ViQMLou1mLq5VmG/4uu4YZClVcTju0bzrX
FTqVMBceSIpUyUCunwV8nbz5cy9XKwXqYmhpn6mRmNmB4Aq/sBVQoZQXBo91u/pp
4A2ZHHGrt43rDxeutk3fD8GgCcu+Fqf2AOsW3DnjSr0YZnNj2I0fb8hzkMqgh6fx
tguLUdOP4YD8kJUyl0wnzS9i5wqKLnMPKqffHj0KdkBOq9XWYOJJkzXq+2Sg3baN
2a5xDWREERQjUQHQ6J7G5mxnE/w/ZD8UdA2kX035/Z6nkB+7+3gMRrkq7Shvw5B6
8iC3xQnOr/6CytT6l6jK5WkYNJhy7CAjytmsnuxTJjy3QbvZ0QuPWMM9f7/hK6DI
S3X9OA42hzbhUR1UXx2hUEnt8rKmWJCQj0/zSuiZrOLhTkEfrAJaRbhZi3uY3dI8
GuUmLdxQqRcX6XC4gYEIlFCXdzoaSAmP5c+iakcaU2zgUWC1Anv7Wccw5+Ku7cyz
6EXM7Y2EZIaczVdp+hgwmS9gZvzVC+xxuMedBLx6gDZvd7YtADidwhhHt1OmlLFn
KxK8OwLRWsOk2Tq9jjgbCKMKvLcdL3plF3iUAqAqeAxYHTzmXcjNj0SxqAkGHexI
0HN3FUTfXcx8CDRznwA3ztzQ91TINCTO7zpN6LQq8z3ChOUN36mTZo6LxidZf/QE
JP3RBLFcLQpXKwcGz9rl/PcKVgNcjqQrFeIyDNvU1YM0i+x+oiJlmTuo2Q55fQtC
vDc5Yr98cSJhItYcK3XuPAawsyRulaDkvWIJCmyuVrCvWumoYe5OwpDNmu3+k8G7
6z+m4eIhwFAxkLz9v+745Wutb2NdmkrhiPECuU2QjtluBgjiWqrbuUgCWaUeajfd
40IMbPaI5JN0XlqLAeUA41tJ8OvP+Wua8ingLQeG2AhdJu1ewuZUWzhNz4xOgFwb
TYTDSKq4P8BqzkLbQZTIAsUULCChjAaec9yl8IBrioXKBCiYQL5w41FvBeoZO6Oy
65qolQqWJgPtiwlszyF0IDRvouzIzrhcPeAlrfAv0MrJu182ju2KnrRTEOS49VaV
fTpZ1s3aFM6wSgJnLjXYIcRmGYvC8FwbhvgNhJAIeHMkL+g+BZJ4IQNiNRWTUgZ0
htwhyTeHBi3ZTwhkj+QtPQwgIer6kfe4XzNqhETp6GP6XL/BCSeeXx8rSY59r4p2
OYyUS3ZVkyENPkFc4Mg2yYaqQ9zSQLYlAvtfz9azFn5ZcF/DiTcbhVOGE8cB7o9r
GrL4ofn3ih9l3tKHtvo76r1JNF/c60bjKzPfpzSOoyAHwi+l7ITxL+gJZaQ8gBNd
z/nxFIfezqaY1TKc3zwmAhQr1VhBAdo+d1C0aN66r2E/mkjs7NACJrB80HOmwYWk
99IavF4L7Ixl3GmdvPMdI0CJ43cRdVCetcrObj+mkXiSXRLdSc+ipqS8+chMWxyl
SBr5dpPJHnNg2m0zWHoLNXvoPayT04TKlvLealOXD3kbGQLsHMEkSv60ktQJmqVE
NtBdsAK4XfOkF6yKljEWUkt3T+enrmBNopz3dLzkdfTmBL/k2RRLQVZfoctypr98
RAOpH+BNVTzL2mY+K+8mdGBNdmShDsxjGbKHrEblEKmTUjO0Nv90LuToMVUq8KKQ
n3FVLKaqNgFMhDPXsqN14TA8Q8lJ14hjmcPMPcVeoQI9LG2nvyWqpgJeMzFrkqGp
Y8xR4pIEXGKsrABmb7y2auYqvkcjGu9K7j4yJFhfEHubNXbSlZgm/YxTMkNGZQrs
zkafaATgdGmoamydZpTRyzn2Ux5/DQe1ds2AlgYU1+nrnqCk3oogO/fhwKicevnp
scJRZiewjrnRYLuJFXbuGzijeoG8axoaBr5VvEL+Y+rhIWTu7OPow9PhtDq/B/bW
ve7ZKK/qdIjjsXNNmcJ2kOdLvaMcPRvx8ev3KzNo6XMsGe6lEScLRxCZWtVSB4p4
4Wj/8utu7k6MGRoiMhTtQhyCBHhJMzGUs99YuUIPyNOCc0pxKz56QWwZFhBcypo+
Z/bpxudOMnbqR7Ol9xxnKRODnv+4IRDioeeGzhgp1UfvmpkoJvaWR7HRVtA6XUOF
a4Yx863GsdfFdcvnCZ49VG/LiKeeFlurTEIIyxDOCdkQRqbtVUQPy3lprGEH+aTj
EiI2MZ0Uo3DPwdE4d3edwbpvzZONnH+Uz52RU+0k8QRMxPW1FUJ8gyCjOxDif3ux
E1mHETZ/IUrnuo48a/FnRI/zvKcc/pq7Cw1AxRPL1j4Zd4eLTjeLCO6MzrKNOYEm
QifgImfBeOtprziE5ngU4cbbrVsTX276fD4HFu38iRMFj4XUw2aHKKbyyl0ZfDoW
E4fIxdg8VuwbeMh15D34V+a4tlp93XEpv8I1ETWIOXx5t/j/anxq78FTH+8Rccaq
dLYJ6urVErOYRl/3CQyVXwUlbzeBbOX5XAQRWzuU16gjmsxBQPlclJd91uWV2ogm
UQa6w5duzftsiNMvZtrpcqyAoi/wrGafrbawC7Rwgh+GxIiF7Z3q2PUKPDP/ZNRI
h7LQh0dMbYTnjLgnSso0LhC5y1To+7OmSlhfuHbghUJlMTVprgaL+fcU7rT41KTl
gXHtmg5yh0szu1Fuuf0ntO3jcmCZQDsRRgn/uBzumomDgjhvrK7dqoRAHVCUB66Q
lEHQI4N8NWKehScHJQSBGDDeC95VxIx/VkrNlX3UREacgfwXlHDTlp1d0UpyvzbK
sNTTAL4jjT3c+4ETcK9NK16ldwAe10QBhzKqsU62mInBcE7e+LPDp9/tBZdxVPoB
HrMnTnZtwMWP91ZegKPWeL8U28jSS4/vCVrEHWJWJhZXc0BTzxlM12XN6+itfW8+
lwGtww7B5HPMcAsYG9ujpPVCGj8E4aOrxki8vv4AsSRUtVVGpbHqtxdGoW6hZKN2
cYHis/TgDTRCu0HPA0dIhlEqbIVyMjeKFhlmzcc9VTKVmLy27/KCeJH0OATrCh0j
iB17cGFhSpPWLTVUQrWnfTz4ggJcq7QyrzIVWldivoOcB2wIKPw1biUurZZesucV
/5QyCeC4gHbDaVVlIxTRqnud8IrL+44eWvC0inU1rPnrrcH6DNd+rDKUfnUKzsYO
CsgFAbxM0JIkprTNZPCRgLX/axlaPpgRZRLEO4WgtpOXuNpExN8OvBUGRBeRcKD5
0GydRl+0PtGOSIF+D6lSQlgfbPVTkUlUdUeydlL7Y8ilX3SqFSHfYcYST24qqTEQ
Udm6iXPaxAkt6vzA62zQq4d/8E3Lv2v8c8LrBZS5L0lNvZi+urIcReP1SQKxHhnu
DJsVhCo2FoZXzX6m3E8a+TDxvo6ZrLSAXEFe/kOOXN7amUygj392q7mczb+28/sl
V3avTcLGxnbWbYtaffPkenM/wpp2aheQQk04YmGioRsXs/3lfpy6hj9c+ihiEoNJ
at7Iy497i+E5uV+6pcAUCLZ4p6I10wPv+t5Oi7iMPAR917mcOhDxTvySYbS6baYG
w3AtDFtxcI3CcOaQoSfRDgT3Krm7IEKj90orftpNFsaL4os5oj1IBVwRdK1SNKdr
hnmAX13gIYg1Bna1fIdcYbFdKfkwXetzOViYHLFatYzXrv7Zo9PgSAhi3EZ0mjuj
2cJnbCyHYz43P9DraodnpDX1J5Dzu7xcykUnNR94nQKE7AiEQr68WNpK7S6U1a0R
wTtFoRau/b53XWo1J1hHITUauZsG7Sq9DuH6IKs+XTu8Y1uV0eahWgARmTIdR82W
D0lQpohMA6wXIebfaRy0c1zriNx0etzfhN8sW/UqH4Lg4Vj+fWi2fpk8Ei2Fz8Ef
dPGpG7TUdn7TfXQXh4OePZHrVnxYU8kAeTtGEu4KscwP+fU9788nsy9+S/MHks6a
9S4T1+MQjC5sO2ANoUCBFoD8UTEapGF/FqpggeYt+rvWjPhSr8BVa1lsQv/Uz4Fw
SDZvVxJPJvrJSm0NyQYBdFnRxB5TxNBZMmbCXFn/hsfAzUN2n0/A2e+Y/TvgpooF
yU/t7hkrB0VcGGG2b25Jv2eOZze8omPGi72gIRAGD7/vsXHu9rY0vSTT2W6IZhNX
fK2QKTtSabCPV49hreZLr5oC/hUh45vy4BMiitBkPWVqDcMyt0w2fOEeNM4q7p0d
11ry8cghMZ3Wyq2/8UagxaLnzAGisYfpDvDfiArPRHX+e4PKf6qIB2Vwod3KN1//
+80wl+yUhqHkjIXd0SdV3H8FpkIpda8zst9tsuuFGgT16l796AGPDNfNfkI8kORD
ram2TqX7zUHjgtWjdFeE7ANomTJrkbAq6nXx44ei1oFv4eEH9gV67KjpeZCgJ6BX
NVHKKJCzxvpAR7q7T1NYxctw3uY2S+iqxNASJN9JnwZBO5nuORYD11UlABPufbh/
u7J80maKMN72kCxUTrqocnJRA1qfSXmyrt5C5+xCQaIQ8bjZrbVXNV+YWNDx27mX
xy55WJn9f6AuBdvzBGaJ/K27L/bOAP3W/11oyadDxn9pEesOxXSZ1osJTr8AAiF+
aT3F6SLPRgzI+57I6Nxz4dyTHa2F16EH3KKoplwqCFdPDxncolW3sE5j2416l3TZ
qnCMnlLSLviy6zqUO9l04JAcZe1T9JK5J8H7S5bzeTxHGWB9Yhg/ddGuDYGZXPJF
Og3LSk1xNtpbtWSg7bDG1oLr013ZyEeqI0YrejwqIIh+6Q1o/uDfLYkIZwIu7QJH
haUCTWw/cjb7+jfiYYpRVq/l2bYQUkNRvGsMIIkS5ucOnmeV0D8iJepzcGfX+HQQ
PRf6AplOv3WozcODRPt2xw==
`pragma protect end_protected
