// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZCTIi6PrvLZaMXId25eerlRnNevHuQKw/KxMekndX/JhLziGwksLflopP03nwUoc
vs1+3LH5EwcTgAeX1Jyww2z7evWR0w7lATj2d/C1uaeQjD6B7EIj4HlEbRxUmju/
Ox+B7vF0SXwlj0kMbauGzoYQtDytkMOdhCUjiVZ2PlE=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30112)
iiL7PEIlhjSACtmfewCXbyhWuCQ/BD3IaooosNO+krYW+E2h1CAJ0fobsJitJcSL
Ts8kNCbOcleNLFOxeMOCtAsqdbg7aU14q6KXP+mqNqXZ49f6TpyYdBxpnqEVsxRd
NGRCxdDDToSNO6J2oSxasgS3lF001/oqbXxeuO/oHphNLX2UYPoKYlZyBRX0/157
kQ72+VlUXSZy2AE2CM+7g4Ti45tw/ZQg6Piv060B1tyixXFyR3HxTRW3WkDEFHeB
+WkOZ3g4t/b3gKxx6H5MVszgHxekOcyGDL0+PabLrLIBUv3YC8+E9dLenk/sAJnX
Gb0E0E58tVTiK2WPoOHxUAu90i6RSIb5e4NVATbD2uvBqwAbOngUb9qOQ1N2jtAn
83FLpJomA+xVO9TbmqJE5RqFAIKsN6O/7KArBExtVF+ykD8q5QvJwLWbbhpJuhHN
GHAk4vO/PFacX3OxFOrnEPNy8UWFgvNHaycEMHsoYODKolm/InJFSGaAO0nohq+G
ZtPdIO3MSXY0AVpwlh5DefrHyVtZovAFX0/RDQOwcXI4FWJ89ZgIdQqrjFsNmScY
xZwrsE2EybYCnUHXDf50eEBG3SQLes25zUeuJNf4gAhLs5avp/+qPWYd6pmbjRwV
ujJ3dCOgiRbGqyzO4wMVnqxSqVzF3fRZZTRLqsarY+xV2kb7y+hDNAGqTc6FU17Z
AufxgS7VzMAeUuKZt2WBexoO6gCgBoTkvJ0kAtNE3FHWK29qtg2p4FnQVdRodGyG
flYnA0IeP4xi2wC9Xej4ydExYTbgVFtp9dXOfcRIFVWiEt2Mrt2dmt171f6bGTtG
fZZ8UVO+oXn2vLWXbE6og8j1zmkZPH5yzApM1trpF9EFvceaHaskVJy0MUciChCf
145ZicJZuo4vtpF4epaSJXLVCxjBryHFgrjC7Pay5aBMzjS+i9LfOyBrVPJS7ihR
EEciSiMnfZe7Y6xZNgR0EWdjkaHHcmD0+SfLLQGeb9L4C7b81Dr4NNfVPSFjtKBq
pNBxfz5lmtb2Gm1LTxENvlj7hBzykyy+75EY1Q6GLV+6lBs57gfpcDFhFyeJZMV5
J/hl6tvYNsUHFaG/CbxN8Ew+0jhXc4GoWveFVjxdjxwamvVhxwM5kglp9mZiTzsY
DUKWUZ3OEZRBYG7HpmJNxrqBRN2pfBqxVo5IZQJK8P9L5/ZkmJGi2G3eKvUmUuT5
u7RoILDiXqU5H7NMf1/P/YVI+13qyGD1fz0JHbmHIsKdhAyFWOQ12XkvaymVwZL4
EEFeMOIoTE7aYiqLwMAnjopp6aocukO/XOAwZpeVhZKlppDpnT6dCSCLB+wFsMzD
GyEtgRKtDozhRDs2kzSi76XFF1OFpPm13XF5w3O6rKr5Tzelq3CchhvF401H4Eie
OL8vUYgHwanXGrhY4+fyqDdQWtuSYzH/x+ZkTSwCE9u2Rt2lXibnayeDK74+0+0e
qOVW075TzYkkSh8Ur8CQWnQncBE3j666cahw/DItwCGWp/dbs3W0OlMCjfClImEj
ZcUpiOxBSsLPK5f7Amtz1ta+B8zbvZh1sJGl39enWHjGLIXRluYMhRlmefzxvH3f
FIv9h5rmC1pr7oMhnElrwThPhHWv7tgnzIUqeWPqhO4gjax7lfeEwJ8XSM5wDmPc
W+Q7KO47tDN9PgZKkS8cFO+kBkcgoaPKxBCzNa4WOhRhiUmvJO5fYF0VabuzOhLk
fHVhYoU+bB9satbB0HIvSrrBBfCuMsc//VHyx3c50HcTyUMIsxbpOKayh/NLMsqS
rRfC5d7iS4aYsJcjbNYwmvgGzr4YewkwwaKlI4moy9xn0emLGeB6jWQdA1iR8Um6
LUe6dAKbY+eqagttxipRmlYfANLmOQSBv4Gs4+3IZzy0zQrVpzNP7V1LoTksBDQT
koQL9tO2SQkLrhvsBLtOzTcCCLQaX2nrefa2HCPAOLVXK/uMJK2eKV1LYs0TNCtY
OmGlGqAf4Y2V/zfybyQ8UFLl2FkyrBHw7zZtGTq9r+53sPP/gDdpKdHkHgR8PozA
avLkMsDbR3jh6xooV5UBFiAGUXZEv2tpGL9eVEkhLjt1yehY3SJgZGUzg5wsXmqi
2OiKxsFDqOJunNQlud7KXz+uRDv0lRJfhhAXVeQh7RTWm5i/sNz9UdbLcI4NImW+
0A7KC2kDMlckEnd02joG3cVo8fsvIb3Iiy0EWmSwwbQ5apYkDTTX3CxfewIFotiy
wY6I+uuvJlUCzNGhMgp0O6H3zQ87Jxr4Jp+k2DY8DnaajOuy1405wnxeq6qmkfSz
ZHd9I16vefwePhGejRenBVopalMJWWZ0b74e4yRrEU06wZBs3qGmLydV1pXCa1y0
nw9pQ1sGEFjikq3iU43KkLAo2O8FW0NxtZ99fOAAVE+Hd4QUO7aQD5s6oK1WSi7r
NqcIXyFqMgRvgxXa/H0dua1WXp/Md2pTYg3UdKShC6w3EQ55WyCW76o0WbFHuTOT
eFMqGMJ5y3XRRU/os3JLaejJ6RvCgiTtNSO0+RWRHHtoRDW3AiDANmqzaS4BTtKC
2ygTDT6v5+I/vGUzdSs8De55Co74drvNpNYgpKY+oidDQ8LKDzB7wFyHurjCEAqJ
o9HOmmLfG5i3okg06oL3tszlAQSxyt4OpZHNQhIZQHFq0MkDeuzWuZLVRrlbymFr
qjGVRTvhMlE2dCVURUy5Ze8gePT5JJINEmpMXYSqnmiLQrtP3rQwiDkkjBW5X6Ob
U12pYC3bn2GEAErj9axA+/zXVGfrm0VmCWdmcF/iDIP8VVZxQxB42svEs6oPLiVI
7vNCDwakdNtgjBeHtsWPqWJ7PahjiSTRJXZK+uM80lB7hX8we5kIWdR8zxlKKZAU
TkZgDUzF4qKlUHxWfRwkvObXn0lJ21Ym58PSvf9CM1Wc2LqxfO1F/0/z1QIx7uZA
xmc83WM2L1tpSH69MwP6c7rN1BBcdpubt/WQ0ch/Ek1T8nQdN+iVfCfchtx+iHYt
/zimFbwnGW/l5e8JxsoNDRoshx+m+m4yQLzMT3XlyEq1dqy6sf9NzdXEJaF7iOvq
GpnxddQXw2nM2oS6tCK8u4HhkjZT2SSSL+JiL2/3Ib6Ozy381gTdcrKAl/ir/baZ
L9oXRP2BvjA+P2oGtcQbcRzB61G1P8lbrT73/NBWx+EfnYNgbEd9rlu1Cq8KugJY
jC8Jk/TCN/pglBdEK+l+Zaa4V8j4hJx4wC2nDKUPCrU+HbbhS0xVO/oDvxcABRDQ
KrUlHmly9JQNAG+s3tdIGpdw4MTWv/1RaleSs1wVsEvF7wH01ZIm8hTf9i1vGmTb
S5egzzGueh3bJD3ViOtQy6v0StdA8tEeQ1c+MrTMjJbzeeLS8JCgZL0YcjT4KTow
NRZeyPrdzGbA2dJx/I7xuFW98sUsa44wLTET4RyFniqPpJZMI/w4AQMOt7Jvu223
37sgOjwK6WANnQSszOq34RitFOvslcTbfxJ2ldYzbhLMrhgpo49hY4ExFovHUZTs
MfE/FRcr7auaQyDinljdSkg3neFpqVA0ao+jkgDS4GR8IPowduAi6MI1iAYWrf/J
VkwM1u/J1dkhOAuo1jM7kX5g+jeTQeJ6bMOmPqjym1RMW2xJG0DyPgQ+Ws7KShQN
ltDE6a9dNB6znI8I7HQKwNs1VLP/RKbB/kKVm5ON494U1GFGt5ZiIcietnbmV9MY
H65PPRyaaktCj8oVBPHR6B5rd03t9aydwdx/kvj46eo2N9aVUu1jzjxf48Xx4vGY
+MkF/aeaNi+KXlkiMCtwS3OIu12xSLLykx8ylnaWWABI4AURY3GmK3yMWUb+zNVe
1qo+Fm6AdVOJpaMQZmNvVszCq4AcSYXJYMtnvsWpzBlvlzKeMDgMk2e6zP19qNBf
rKHAluce4/GIJb1JEwmNuUOlfnZhSgZIvPCXWh94f7ZBHNL96OVumyPeHWA5O735
Sp+SajCPYl4CLPLdZYQHjNIc6z+ECo+lh18UItFJbCnkbFdKSCPCmjM7Uh7R3UMq
fJZZ1yi+r0c76bg4dujZwc6xJdBFtrKLWh+6f1EWDE+9BrY10Wbs/n/JXJP4nvS1
vZZndN/rA3M+1+r+0L6jclVVUMWLdT0HKdj925dcs8f2inG0IguA0q8jLt9Til6e
/Gj/V8f+mFodZatbIdLnQdv+ifRDaqxmecd3SoGrA+MO1MfwzxEs3phga1oJahPD
zs9PoZUtBp19mPGty9rgKATyYsgmx+yuU2M5M2iUnIufIMoIvqRDXqs3B+ZF0I0j
b7K3I8hr2VYQTSGHfQrjuo2ifplMRZ01/SIK7NUbsY1jMhxOGgpi6tIOz45SZURC
T/xyv/5wZd6REZI9NjGdXYvEeDPOWLHoX/b75wvVG7t1cq6QBYx2bnvxVRl+W6ta
Tm4x7UboN46G4JoEndLrpETcZHyAGbZ77aLATAiJaYOnB5Ab+gIBYt1FFSGyEDTh
bVRbPJeHL0F44R+jW4qk7NQcfxqVk4wSJeflAwERw/8IVqzD4v3qsCCWAIA2dm2h
RY7CBCPL7nVFS1ufgren1PT8EnFTpBi/MOX0oJ3ebEIphCnuxV94PxNb8buJo/R8
Ylg65gjtZKNDVHjlN+68G6PePZjZPhmEB6yKETFIUq0DakuGYOZJn29vlFUPYfhD
ziixk1Ag2kYlJZGnwM8jOyyo2oUrPjLe2V2GxQ1bY8FsOC5ZtfIoBwtPpc8hRiHx
Sa8gDvZTYLH8UBrvJcw0UUK9OjgH0Ne4yEHhVzpyCtC7BYRs36IcXUpTIDJvsBrK
zk0g3N34zOv/k+2Tq9hfZeTIX4rn+D4XvnIHMG9KzPYoTgICyeWnVQFEqCjz3hZq
RZhqvNI6U3CF8kJaleSid+paSBWJnWD2MraxNihg9L/Ksn51o3BkcQok4TZRJMBx
6RmRgShtvY1QJvVuDN3gNsmQD08JmiDq0YdeqdxEpqyeKb62FSmixS6fqJurdrWy
C/QqHDbCGfow6TO8NEypxgleuqb0j8eRokw0MjvGA8xsdDLphVaWNKZEuHbadh8h
xlkI/NrPFLiTAkKwm2nM0973r8BmOqPJAP5DrNAcO4CqPSs4jhRKm76lKUasea9U
6iulvJyniTS4tOjE8TYzEE3wwa+lDCLxHsX45HXw2oiIAFhuLsdl6W1ZoO/+2Q+x
FcghxIdpOg10YetjvyjSsnKjblNbhS260DvB0bVe1Ype2JTU6+l1SmiXWejL57ue
UUjtTNFy1VmpyElJtoInJ8/tjZNTP43jAKiZ4RlvTLmZE/4aeool5OLt+emcKqc/
rTM9SKlaJuw6RjhCUIWsDlODOG8ESTwGTMcIKcEEu+divMmcYH6y+/JhFtKTJtz0
+wu8eF6DsoAJV0F0x2iIZSq68cRUFwkHSY6VIlceAazYSnm0ozW1ss4UZB8aakr4
xLScG4zCjqK370mKq7JwGKEFKjn7PhrsV/h0Z5jWjfAB9teFSQ9zAQ0dgH8/cKhk
HUtAo/SGoaQ5NFKT6XjiJpJtIrO3zyLPo52J+tSHQMMKAKyF7gGV3HDxkFr/5Vkr
zJXZGO+/Xge6ncKtYdtRZRtrGQo2zdNrp3iD46D6N/VIAl9Fc4bIM8EVAydwN04X
1Efw1YMakM03QMsLC7GsJwP0khgnF5rfoeH5ifc/GOvqTeLK2KQ0EhFd1wOj+vWl
UqVLdzTCF2H4wNk3OiXHqzIGmuPu7hnoYHHULNkcNKbQ+RPtepCiPcz9phZhiD+2
0UUHyMqMKPbUDHuvoji1NK/A9XfAwRwcXfTITSbxtXzav/YlXUc8A9KEPHFpPksL
vOM0Xdgytyq2Dw5Zgn+3K4bca3g25VFerH1mAPGDiZbLrDcNsIevVypcUzocpqCs
L/dxl7ZBCKeNnEdv0sA6ENY+zhf1nyxprKZ2GzQN3r3f9QotXVYhD8HJpLHpVS5B
ODYGXj8KUo7GvHAlJz6a369FptokIpqNkbuhyqCaiLvMUI3wxTBfhwInQm+4gj+Q
Ba5OYB6enNN3fIjUptwp0JFRs4AtPvZl4UQnCGW4KPsOo5BHWEw7RsT1dPkMUN9t
0PIcGWVt6SwyfoChfC7VKwKn6PyPjp/vgjurfC4gsdzYjVtv60Ixt+mrK8zJPw4T
2OgeMP1yswaRnaMbXT3oaD6Vp46/VsXh888wHg8fUe7h80mYVzbvZkB+QptwYrBj
0jKphCo3hO5APXd2Ckp/8lBrWKQdyPzyAIg5JTFehHSOMKASgMMdiSVchLX1+/A1
vRx5PeuRuHk8RFQt2ziP8WCJQroRF/cRqcfGtR78dIdCD9htfChsAT1L4cEU7Iur
LIkQ3+ePWHlH/JJfot8vPICi9p8MPUMnUjoJXq7JieZI++aU2SMIDO3dA7RxXd/F
2FZ43GSvPtHrUx5kD8ZDPeoTCeQBN0RjBNccidp7/xvruWeEgvMpM3p/sT4gzPHs
kIbKoeaXSaZZrrQHFUJSQsVS68K61HiA3MQrm2W5cQUDM1q2760t+Hy39FbLrIdw
qzbjrffOJQkYkzjE1FZBsqooth6pbo6KQVztfxWWvzs7KSh1BkBTJZy2BruKtjIe
biiEZyDz6fsvLWbwaino79MwrKizEEc30CMNc/q+ZExHjc93mPXdBVOpyLCAzoyH
zwrFeznRLMwp6teVqXLM9jHclXbBYWxslUKUJF4vRxpcpAA1uR2naWvHJW+vY7cm
O2ZA2OkBLAtxN/hlL5U68/9qceS0hOxc0wVyNyscxicAwcraythOcDG/oh23K3If
sKSDWzrt6DwfQK+DhcA0wmePmdV8bLYCjvP2V1eN+8YdJwaFxCdVkYS9LvK1vm6G
ha+2CABjDOpdebzNgw+7SCIgAxFXif7HdgThZSxIP5mfVd5sLwWdfjwshxOIBWHh
1d27ILAKDydkUzHWgxwAiPpmskzmbfRx29vvnJTTbtNNeX7EkjQd/2lBzhuRVE8v
mEpFDoszz2BIEos0HfvsV74f3H7vdIY8Eah3K9cNGXxq1cwHUXAe5UVXcJJ0jZgW
x9TJEs8+5gteBHxVsWWrja3krFuOQuKc10Clv84aJHCRDTXpO+HdTpOOAW185r+Y
yw76qjf48Z7Qc1GVfchTMxZyhf5ETNzw3TS0Hgv/AbZgkReapU++OXUJZw8KAAq6
zEmekzJnyWPPa77x4NO8O9chMBJbe/NkR0hALzNOp4vdoepybLEUBBuiKibCVbPG
0Y518kGznuIkTQoLXkbSjcXxZ420kVEvvojaxY+R6reLEWoZHyuqZoUzEg9NA7Af
DNn9wgFZEkaIVGrwL3BAEmiA21yZPmkqOf3FcbqyBfKMN6cGcbajDLCUrTTJ0RJU
UJvcLylJB2h1fZlCq3uqMcXsZ8X8x41Zb52zPCTpDdktmI9HjXK8QW/dtY+E+IlS
uICAdvAN6KdjpoOcX7H0lyNn34gVmzucNBLBM2iAiEA9wYd+kboS+caQMIB1Ytzu
9sabGI79x6eQnnA+JSq4Tl3K2fIvayU/YbVWqpCffcXyWvo3KI5T3BCCMXRsruOm
2rQcF5461xbq+AD6fI6Eq7RX79nCuEpM5bOmhXWBNjBQrwXKCoCj0jEReTR+PWEP
sHvKglCeUQo3nWQE0GQA2Qrc4UORucFcLzFLItmfMt5z5qKMVQJnz9XsgJ6HAdZN
fTlAynxdEm9l8mnbiWJKOsgxKSHJiQY7diWdc0WYfYQi0HvVKITfFHt3UoeZjQRm
lrrS31z3o3VM629PQ3bYFSqOPTXFJjZe121L2zLkvOox88GgZtu+/Zoqwth+qrP8
JhSwjfj3VMi9VJtuYrF1KrTummYe52paNHOqFVnjxCLzo+5Ur7HOite1uI3naBPU
QDJ09D5O53t/KfjiuOInzmSho2GjcQxWl6OufhDVzOXZ1ebXOaQZUOaM9/lIQiiY
chGdg5HH+ngjMLsEX09pH5TN8gWm7FUueky2ETBNreoFlXQH1RSoeTvnZa0kD6hZ
9+n151ItUA58zVLBu3BpXxQguncUid6oMKYyJIeO/esBpWLMaDmxHfrWgTfa+FO6
0lBuRUxtaeWxL4u2/m4iB02TQKQw8y1fTUR4S5vC5JKSIyX631otpcW4Ps7qv2/0
nqUUFHjld5jzFNoma2miy+C72x+RVIkewSxRGV6N9PnTXHa5BqWujKg2JajxKrEI
uzwTBUmBkcqla6ed050CPG+M2Y4wTkzLT49fTkYNL4D7d45ecPJu3MPN7llyKor1
xxKrqekEO5cXPEf3PrP5IcCgzX2pDrXFjnZ2SGWGVivkwgZw4jhE1nCpg8TWOPgU
ylfr3UuYBu1LtLP99F3MzcxJK7hl+rq5YlvWN+8ErxIPa6By/9nqQPptYIFgPxju
+pCMdD6rt6GoWReDgc4b37Rg8p2kUml/gfcSYEv40Z+gpvWRp5XdpbbPlnjuBFNe
e/wj5Yd0/QpoBBtFaADO7wOpsti7XTqIg66N/Sdymo7BHL7NdodOn8wxNd6pE9OJ
bdXSCP8KfSuGPaxFhEQB50BrzVni2RsKyIDYn6Am7ILP6czXrb12dOswYsCoZVnz
vQCXd7rQB9SwR82MB1mWVrjr2xUgnJRpgnTfvqO2z0L9ka8K+ikaqpCvLihgUVft
Rg2JTYSVwz6ikPOdZG0bDpA9hId3uoCl4mJ3RwDTR5Zn5xp1MR9ilocBAPeEw+Ia
zEWkb/Gc82HCk1WfMPNKMsA6FAY5x0I/hY7N8s5JRiK6J+V4658X44DIs20J5MKD
IAv38HEXmCUXX8V1NfVOs0C4ZrCeRSCTlmgkam7lHisgcsyPYKIqRVfY7h9KyufX
sfJuQT0IZCmgy+MRmGT9jYdfmP2aOvZOsm2dpQf2arrnIGGOmQm1VgECeJdud4gl
zIo4TKrSu+JFdA6MQ2/n4rgbxP/TA2aYRfzkNByJo0qmuYwEBjUXz14BZjjof+kw
BXu4cMbar1NVoo7YtGZoELCBaiWC57G+QPK0DEfiOhB/JHe6WJn043HihRctF8+i
JUW0CMsxSNrLqupkVhYcsGJGgz60eyyOOXP6/BC4/mUokQUGr1Y9N4Ouj1oQx7GG
AWyRsq4jpp/3GgoTDqjHPVh9Gn5tTV1bWAHMA9G+mE2YC+6WkjmW+8ONIFZTm9TE
3fkZsOmDFT++w5uJRo4I2btepxd4ux1tvmnubfi3+bOowZi2l2DplgnIf+ijB6D3
AaXFgoXBCDPjvDDGtRlMiq1lXe4HNIR/v8VSoXa2svoCfuRHHjLbOIEDGBFw5XJ8
qDAWOQc3c4cTcD1DVJdZKmH4WqOd0FZKPkkl2YanqaVt1AlZEM5ELpAYxp13GrGG
fQCtI+xrGoQ80wRBiUuu3wPtijmTquArfKg6VJkkAwolSziAePihAv4LBf70yubu
O8sozY6+lqwBltGqmWashcpBCSJhoCjaU8O6Osx9TvPy3nSLNOUlEd26HISgVTcV
ig6VCtlhN/lDqf1riczxS6USdAC2THD/GaKnS3ArWCb5GM2zxOqLChO6drawujNr
uzSTOCw/5DIz9fGfDa7aDSsV4T0M7Qf5qlWS3Sdtrl2A9/cIdSGiL0QadVWVtADS
VJINQUIYOBixb7TjFcVpwpRtKmWrogO6mHKMXO01Sl251ClB0AaC6nOPONffWwsM
B1bavt92WFg+EQb5qDVxw3WUB9vZ1lJoTJPQ5OqNTktNlBEVOEq1Hx2j8sQ2g4cg
6m0m6XsvAdDwyuvBmJRSMIE8vVizsxM90LHBT+Z78kOyYjyA0jiB69iIpKLulBHf
RJtL6m6cBhIWmv8ytu1ml2mkrKOGgu0BpZAdzqMv9lGGioIcdrhatBr1Ys5BMdzq
Ra1vchOR72XR8c7hF7YVyFPd7FfHvaDyQC4PjS4PdcIUMiUQ5RmgbqbBMEIydDCc
MXybp27V1Rb20dnqy+0lLA3CFEt/m2YqD1iVHJD2YgLU81cPm5ofluOUbgeuiHdy
XGtgsl1D60qGnQCFbCqboBX631SXjpm7Wvmyv1EsUQMip8rwS01et6yil61JBIFC
oSuDdIwWY//ek8vNyRlOS5ek39KR8EArNz7G5mp/7U1oKIQtzMdXU9r1xB1WywUS
A4+E+RqO48QP6hk43c5/b4YLRlOM011yjwWOL9ZDP2NhLtAcJUnK1FXpsYnOok30
AliudMhIW6EW2G+H6za33+jfsyO+HVM/HcF3HED1xa0TtAY+68JZlu9fiARhijLR
PoEDmUAZH4C6dkC6qnC6jwiwELzPGrjPVNPG0gU//682M2NnpOWAP5K+dqcq7LHF
7PAp2flRFemxM37EaAIfeoiYWLtLYgpDCT0BlBx0Brm3uKzLDShtBtixYeF+qyuC
QepoZlsM9oDsejEHGsozRB8c/8yANQzlWsc+g4nhiSkSthRghbp80y2WFZTZvpbn
crmV3en2EIS/4y74qzy0bPe/4w0ZivXDG2h1pHbV7DVrzXPxuhRkHvO5V/ByzhrW
sOgPpCynFi2xf6M05wHHc2vrVkM6ZJVYvTm4jd2Vjuifd96T7Ei+PperNrv9Ip5P
t4+wjkb16DzI1cs9b+BuK/P1uBEC4Xb6wR3Wdo63WqmaeNhUhW7UTZ/RnSn+Ou8Z
RONj14qMiO8s1koWCzbQGd8gIxyd2peRCK928BCNjXBgPf9nNO9Ql3JnQMZvGMt7
JgiDP61oMDFiOoGURf3LbkQh5TSRWK5gFv8C5SlTdQ2XWE4h4QEjN7sI7x68rcFo
rcUchi98IZdoPgie4tWoF5+M5pKkCI4CtA21mm1tIh3NR/GjdPDIQ2FEFrqSBPzD
jvEkoWxzli81ob1/+C3GgAtOCLt5Gm4Xqyb923rDUcxzRyVsYmMmYhPXMK8ctX97
ZDjHaOkFvYS5rcwPjsSM7ApmFQJRnF0kXt6GkINQSB9UZWbt9a4ueEm3Y/s6qkH+
iY0BcZbC/l4lJqp44LN/E1pNkX9RnEILjCea0kyZ+2XYsti2CiTp3Vp4x15k63Ja
QNk0TZGWXKBtc8kU5pTorvH8KylY7cVqt1GAgcyhY0+E9ROwyWshJJGGajyilKaX
VNF1FyeVde7hnz46f1x2oUmAjrk6FU/hm83eohU/8VzouOLkKlkQJm8VShwNJEn+
PhtOHMV+gT2ydyD8tB4LM6CPiivOXPbii3XMG3/EwEWaYF4gqwPRuGR+1l3WXM2w
5JT/s+SBZ3DVxyQrJODshX9j6nTvgqf5U6dkR5eajSub9nvRYu70OB10uqPgzuFO
vpP7ZZS9EIdxckZkoM+qBHVcvjhzSQTbbXgnwoslePqSjYV5IVtk1stZUY9UI9RL
LIyshpNqdsOmXd3pPw67FMkSbNo2Km4Gye4JU5Rb+HnXmB8Rl/NDQkDrcEJs8Oup
ffZe9HV/935IpUcKb65IUjxrQbxiRKuQrBETO6n/RZ8rmGOHD+4bzhw/Uz9y8g6f
r57trvlzQpf2PyyCWnUsMVigTZLFnbdxM/QlDwZD2g5eWZ2fLD2v8EPBclMkKDvg
a45cMVlEEm6X/EzXzW4AI0La/Bg+5PtTtiTF8LtKKP5Sys1e4OYYIb13XxRCowBL
scKTZX1XVJ/co5+mJu7t7UaAFEG0GwnMcLF3Cgl2Uoa18H/4tDZzixdTJGmCFmOU
2dzOKD+1hoZ7eSStD0zWlMPwMOPW9egZIKuCz1+8KSAvr6f+PLo3n6Oo6oiuOCdU
zWEonNqbsUYafbeHLB3xTbdhs1pUU7yFuxSlSRtsr1lX+c6LU/R3DiPwvHtsYYTq
GvY82Nzn61AdT8jwtbWSAalcCUykmldChJLHRFAyNVTPthdB+XTyBkOmGVecE+Zo
VIzaM2mCQlVOdOFAxXNYK39pYD56N0wKN1UjWQ3EneV8/RykYImsV19H3sFUfthj
fPDppSjsjmJaTgxg9bnP+GSGn+uW1Y4zwvB8aZTuql4My8Uq1aMtKdQAD2/IuFsZ
POhfg+F/6aRI31Ewspk+p4fH7Cd5vuC0WuNOxLDCORomrcIrG3Vw+aI4motjZUQt
UiRcF6njYpkveSZhkpuzoZ3RkAwKYoepeFwCYPMNk8pWG1xb53vwtWu55U8rWxDf
Lfelrulx91s4e2Ko6/90ah+gIx/A79WlWF6PW3fqWO2vMgcR69WwFPXhymQgVJ9W
mX2m8EOH3Ykyjns4RX8RdQWKF4GnyLKj02UkxfRY/99v8phF7/xjWP9sALLndduG
OSvHsT/QyFmYU687IUWe7ZzhDQ2qHo73yqJwPAIi0P4nWGvraxh1dCCgD3GEO9vl
jST4VpOORju62gDM2gNHLPZx/PZtdJ712Xv3XZ7JR1PyjNQ5zyxtTuHXmwvEW1V4
DhUMtSVXHnA/Td+Jok13C5h2YsTaZz0iynf5+q84+oe2vdd3bQYFN7kr3vtek4Zf
VuNKNtU5TbR9dHZ+H93jwBp0rB2LV1vysbELDFNSnGITYNY6STUGzJuO00PvHvA2
188mgP3A5xLZvsr2y8m6T5jpI9wZ7FEdE9AWrlmncWr5GvqyWlQ+hlHltHn6O3IE
tkSzhsYCwPUHEBsQI6sFY4Aefrv4lyKL+ft1vvJ4jH/8CdbxCoJt6n6M5LQSmINW
auWY/K8gdtmma6LbGdap9je959eV9OD1rs39NLGaeIOQoqBfdBjTuU193U0Pypf7
sLE5xtAQAlJAB5ehsXyPSPmyTfZoykoKmaXp9Ts8SmHSvwLl3gaRoMQIDKEOELj7
EpqU4RSxJLomu5YWQQTasfjqkDI7oL9pAtWGoSlaqUO2tua3R+bCYaIjJ5mExLtu
BFvV62j37t/Tei6ytMbqijiDylmTf986k1Jkd/9UkrGb1np1P491vkM33QxYKzxp
iHj+m0qeqVrPKpyhcuc9XFJoKaW542um0dErzbc9Tj0/ndIBmnJZjMUryzEpg5mR
ALuyW7hq8AiPLmNtxQqBKynW22UIypQqS/BWe2FUrmuxPUsMXkfL7d0eSGMrWabK
rFfG7VLdJC/0Q2IZ7exVWd7kHsJrc3l5o9Uasy3YjKHNqZR4Gbt1V5h7qZohuQrS
wJIWrXqEBIvOemI5glZf7En8AmK67hQGND+7S81snvD9kX0c+PrFzs0RggVeXCHn
vaTX1uwkyPMH2f2QW54m3pBeSsaFaQ4T3ONKfGQebclGcXp/uOsUVX+CgKThs3VG
mrZxCApoSUjiai+FFt8KoDJdV7JOfMrwnGV+44AbCER1cet04t+p6TQ0gHlI8R1C
qKDJZkXASxsO27/M32gTClJ/PD19vmnCxD5XBhkQ+GzR8hjqDkUIstqAGaOweE72
DjFIUGbg060gpI6eSRn0plmpEuhjP2B9Hms/XLF5Ye8olsZztqrjOB/KXu+Gzk/c
fmuWJoQ7Lq66yddc9G7yqd5ZPKBiCeyycTEAPd6VZWU7gO7/BPM3HefPMTkSUAP2
K4X4MVRq1xrP+z/n7mIhXtxA2dtiDSh6KQGorWCcutAH6YlcNcHa/sRfQgYt4Zlu
3rCkyTP3Rxwy+zcrRuZhQSxjqYrZMNDF5fkEc+NG4gPDijAP7McnuQLak4f+KfY1
N2/9UD6yQ6FSUWs5VpgPTeZFA9PM6CX5ZMv06qmxtk6Y4pIco/VUfgNRJQOMzLZG
A1WlsJUx2T6EDb50kwLFu3/en5vLvluOv9YseIC6CzXNnsWqYt4PVftnOqCfJ6nX
3j0m7XjN29BGKsbnMhqf3ACqDlb3vqUO4966RCZ0Yonq4qiNiA+UljtaPgtilDy8
CQPpIZ+gq2yv7wAnkV3iB5McOZKsDn3WAWg0V8uDW8HnqrwFCO6eoBrUouT9lpBN
ndU88Y9l7+m3SjZRdPXr7Esy3RfwAEhytJ1RIX5VUFwaLWLROyPF3UKb3AFQonZd
d3D8lsP1SuRukFj1/IvzBkPuGTqJeYQW5W+sTvjbsIofnLAExBabkVr9NL2ik58m
eWGwtiopG87iBJ9223MJ2MIJxY7BAMUWpN6KUxvs+wym3VqMXy9js8gv2zXJWyOk
dl7lAtRMvM3P7Mo7UOpktMdRJ5p5R00EXl1hAXoh6GKK4/Lz/8hLWVKyFhR+LzGa
rfTamSN+Vc7sDTzji7mGds2gqV4ZA0ZVydWdAlixr89Vgu7DEzXYZSWOCNOBrEJi
teqhEIU3I6U/p5DIYzMXmQO5fRf57ZAKDFNFDeX0c+mGNZvG2+FRreCPbEjX2VVZ
oH0KLNBPdESm/MrwzSsYrmJU8WUxgm0Wv1GKekKM8GrLA5diwBe9hjrCCzfrhLwD
Z6Eu/Hgyy4ggRNShTxszIx+cqt+vcBoKpUfSZ/jlOc8+r220A53gBfCq66oa/mOU
ayxBRXSFDmFLgqK+vwUo+6PXYJQZdG3UH9CYw6DIPJGWfuFbjNDgQcIftP+9sFMv
Rl40xpHh+hqAqTTbGTaTMiyvtzY27677KwsL2gkNBCCavjusqa6vZkCHYOIqfIGb
69G/PZgHfFWVZ0YQVgXCzv+O/lVHwVuUCgWeFt5NLgA1O69SW5hYtr1wDk4MRut6
b5sd1My+dbkYWAqXf8k+z2BkFSKBjInN1AIVj8KsBANylme7uYMtIFDtLySFtwxw
HhoaI/WmMhw33r0hpAdoKdzavyVE4qBzlUupgvE+bRUr9VhppqmI8Yta6J1FG29W
/+/mTzKdsK5CvaG9zvEuqlkGNHkyHwSQplmcIyIVQDKId1ftZWQhi6V36fFoz+At
16zqevOk69LGY1lf4DVBSWcHNX9J1z+S4n0ZnXEIq64I6QyQwAPmXSl+j+IhbGv2
JLv2mbnVBOSVjw/J0vF8D11/OreP5OlRpP3w/tBPjA7lNWZUu+ZhwtLEYHuAmqAS
SB2zR/oDS8oj9wQcJavYBiI53MXLZmgzjP3WkGcVVB3aJc//iKq5auoPcBIai3vW
Oxn7fQUjIr80r/H+z4fZFH29isXhR2acO3vGBKIQIkMhZEtva1mP+aSflT5r/elY
9BymjUDYVHxeQwmowfgDu88B1MsnhOUfJlrnRipVSlo1yVXPqS9X+SPnDzlIdpvz
p8Q3fsWQAw9TUeyv/MF1QEbV2UIM0nCH1hOATNmrBim/XMTFtvAHKcDjGismd6/J
HfXUrQF84t40jwaleGFfc4HtyBw4zxQSCdF6ioNsbMW/q6htxnVuylpTGfBGJG04
G5d4wmFL6H+Q8ab/VvMCdx3QmEnk/sZAa1BmQsBCPf8G40EVN60ghB1pvOt3Lgxf
81a+2ZnU73DRejvnivjMOAx3O68flATb3gTWJLX7bsADL2FBfY5HFEFEtLqeFK5f
xYfnUf3T90TxQjiIGvBr3MUT7HD2IXqApn2wxhWnpSk3+zPTEP253bwgf8Mi6/qX
bqUawe31HUnmRKEoz+3zOXSjY3epG2nlv9GzEmebY8uksEh4a7Kc+Xe2bM1v/fb3
hBzjalsPPOoQ4I7g+BqOwPiRLwzEd2ql9ZL7NePuj0ReqGvdyUSB4EsP0OSX/k1Y
HX8pA+Gxp3VSm6Fjihc51rbnz3yvPPFgxkVdaS9Y33GwHvoIGtg5kdMxkdDehSfo
wAwwr1NX/bfFRV6pe9hrxNHS45iZ0eB+adzsPOwJNXML20Mj9eJN5htnMualyx/u
PDWWGH25nvu8lKjveABBY8xhduAjakzsH+vL8h4zAKXwMKNnOji0mlbs4adf3gpr
GbVfCgoWQX3Hx7Oj3hwhhlQoVGI3ZLZbbOEES1B3urALby2+vHQBZwDKR2D4gl1L
QhZrw2NHw1T+W1HNC94oi2v7LbfDH3Wlbx/s3DUmxMjlaVvYqhenyXCZyHD8RrxO
ayw0RcsRZMau0ihQAMFZk9BzQu6oDiwTXVZ45FsSz4GP17xITGCVICd9F+2olY/b
cdtqYQAhIDiBCZAxCJhK2NXgmYxf78BZvCdZA4nQ3vqdmYeRv/T5fgMvrOGpyL2T
HC4cm1XwfnhZtf9+XYS5dF1RARUHx9lqW4MW0BlmOnWIi6KAZ+6yC+0D0zuRYmy9
Y7WwWqxAGsPAYdn5scCGR++OMx/jXM4dGRHjJhY+U6lSU12bIc3SYHFe/XCUTU4v
dr9bP1dnwX2vHsEJO/dHD9N32N+qAKd+S6J7Y5SAqf62N8nI/pTdYom+g6UeVi1H
vfsXAz5fpD5FFx7Gjv9EJ1PM2N31G6D6TXb8YgAL6zCp6SWjOTYr39H+uQmuWFPz
Lcp5zkez1+4fV2IuO5JwsfczHf0HhkFCQK2CR3RdaIqe15RIhm1nuHi/xhl14/zb
6M91KZVpQLfJ4cDjcQqHPrdXOTeU370Kbi0LruzBemmDccz0aoyjngjThLMd67op
bhUzaRdw3KQX7uUigak37pT5gE4s7J2BBIS15jFWyB6ci1l1elmRrW0mY/Q2f8wd
ooPNRa8ajxv/e+X3aFl2vaOZBluHAQldmTN802FVJEqx1lGrAXlaU9T7aegEJShq
NzzK1w9MIJNHXRLnn/gxba5N/f1YPOw2nyyr/FOE8OYgUHMQxGHAg/OswM1OehNr
0WuCZTQxYySSqJH5+48X9EprWAYHM3zmU/ehFHms1ki0Ol2Z4uefwemzK/GgTQSW
pcof4ly9jgL5oD5GkHPsiSuru+Y/qw6rHizditfmasLR3xF/XpIv8kdi0I52hMiU
0TzuPc+pwhZZdf/To7doOtaZ/wZ0X6LSg0yCSpKk5fWBBvEAFaWh5Z4B3jiuCyWi
DkDRsCPHDbvvc1cSbzkNPKpEK6QOzNt+hvs2ObjrrGMhSxgdhhErekwcyyi6DOb7
tYMl5tZu3kqKdPiQe6960VmtyS2mduIWjlBNqqO0o+O7MpjPhETFmy0XrfPG/P//
wONmIZ/cKQGAu7+109ZhVa/htSQ2vL74ANntRY3Ma7A//c3TN/5xR+wTazvKOU5n
xBKUlpdcviF3Bi19K9aFwM4uSKWyUUfnPw9zik2mwYNgvoJNXpX3335/hYdeIQJB
r0mcjjpAqCfffuCVcKihTVLQ32etzvffCxNp3dxC4DwejHnjK24nKuRTVbAE3LT1
VgMCWvJmDR1b9v1zAVhugix3TbCqj8JJInaKSP+v2jNFAqGrsWTzUDuATEj76YrK
/3zB7Uv6I4z+wFRFgDP1xV46t5uzRE65U6Tk75Gby+9pOa9WaBEYz56WKDFjviZF
5xrfGteAMtxh4W63L4SoXo+QMdqat4JdF1Q/ac3WOHTPFiW8PrfmT7G1ZeVcupT5
xzn0+QUrJdBf9axBAH3gvINMu3quxiiQziC+FZqfk7r590a+KYCiogdhKGQrAJ5p
ehlNwaHSp07vcBhEZJ2TCzVloAgNL9YJaWZRbW6OTtXg8ZWv89UKoIsBXSP5ozlp
PN2CYHe6nPT0HIcjwkPo7UgqWGB4iyctACDsrRXmo+Pq6pC5KxYDp51q4sUDKOuH
uAkpVJ89By/LzI3LR3jpSDOA10Z6a8lO3yK2O0SvMimU85sQ5SRqQIen9Zv8aCCg
6TF2s4XIyapLUt+DWTx98A5BSl6o1A1gjNvZtiUQM9gatPj53lvGRyqQluC2Ejf5
qOP1l53CZMw7mE2PdWgAEjCeeIN+YMBt+kl4gIwWv0GXPWIwBbGLFpSCbzB+j7k0
vZKmdyZ08bTITgRF8WhRezdGS5dFb55f7IsgTNj/fRoNZOb3oNz495m5R+oQZnWs
EOdEQXF9t+TIOb8SELb3YFzsvmYAkmc2wBXSj4kbNLaG0I91h+JOA6I5tPdnwMys
v4wFIqvqnEQ3M3xAhO0AOHDHYHwp+6aNDEVGCZwYUdiCkDWW7elmtuhxW3/4lRnT
eJzKCt6ceV6Rwu5RUZCSC5yw9BuCQQF4WYFOBqAsietXfLdkUcCb0tBNpQLr2lgC
SCcFrAKTDcKuaMxYAkR8IihhUpUe5Wyqap6hEyPajwglTsl5FLb07iXIa3u85qxR
OBaSJLmnsup9bCFBptACYk/Vd0kwsuRY75tbMD3mHOZBn23rdoUpojNbDGhWe0Yz
6dC0bomNLat07y3wG/MqgagJantRm4OwI7Mk2h5VdRba36v7dwFrDzcZI6Bb1OLA
Jyeu6u9kEhzzKMMCE3Ef5x72xCXbGRyMS/dKoWeoZG61gWuoWb8rd6ykx1KfnTQY
BrtMw/H0GiohIfZpUkfaHqffJzDQ351/5+l9dBZw8ETeTl8gU9eSq8tDH8TBziN+
Ac4sWcMVRPUkNTc6vDBSVn4SIFPct58B1Fbvm/rQEhq6/1+SbdeGRetS0LzXCwGX
6zFth4E3K3XadKyX1JoK4GN5Rj5ms/CMIpFKFnGjeAbc6D0fRcnLdu/TxwjnrAzI
4F6k+AlwI1R3SKkvFnfIAtIfENliuissfiHWB1cgl+j8GY1w/W3iMQgsBjzbgWjQ
dyhSPdn+nVHRNNA9HLBa+8/Vn2z0UsVCQhSpYneR5P17DmF+/Nd+EY46bsIKM3xv
DvYADW+Tk6cBSiXeBkAVjL2gVf35qgLN5RnIpgYG8N90CickTw95veIsA1DWzUNO
I4e2uxupQufpTyBRMDLLdB+NfTdveXR+kqa2C6nndHlVGOFDZx1YWbW1bMGby+aP
GlN/Fl92JzRvb0ceFVSjAfILIvZFtZPWpyH9WGLLVAtwHFAAhhqgsWml5S1/WuNd
SQQ8ChAbX18dS/yYnbh3rumh5kettAac175iAtUkRpE4jBT6hDsLKxI4/pbIs4fZ
Dcu+Wllp84vgY4T1k1tsnMCGrYuiznKjUnb+ixUr3bArmbYBTmOfQvfkD3USGEaq
W44ijvsqMKsyrIOZuJzIFYZlyIppkHfMpZ+/TFZZ1m2AbJRaZLMKRZabj8wu8unL
cok7dx+Mw6ipbjMcwJYwEVeVlcvzyoV5fDfc6jj8aUboaHy9NGPeEkbwKBC8Nz/8
zsJiD6ez3OyFjoO3Yh62/A+nx0gkFdhebj6xl/g4FIcpnB8P75VG6w8WXfFU4LcX
modsn+e5iCqdxpj0+S8SeXANW/Xsaoqo4GYJVCZBr/95IP0yHQfeEipXM0QhZgJV
fCz870/zghcXqxSs6B3wcN803Jo+VDAE/y4rifTnwsZiHUdu8hNvFBCEGpWVrsLx
6PllVJNcx4RfwtKHbHnyYMLIySKIwQWHGDk4Nu9acVcNvvrGbhF0wTeb+uJt1bkl
6DW6PdmE9qzpcxJEQUM8CcbyEN+dhAWj8RL/7xgb087Lik5c5UgZRWjNgJYW6T0Y
emv1kpMAZrJhh8F59Vb2dYnjZ/8oPN7+Fxnbz/2PKbtqVHHMnKFprCpYbLFvG8Yy
sHPKqw116OpK9UfBBwJm8b3PeiFVUdJMb4sHPogRMr26Mb0C01rMrnWLVGce+iBg
4tmu6qst3To81zLE9KiPtaND14kmBkjhEteXWRbtCPFpyLbQbTmBgao5QudP6Miy
Yz9GmQKSCgCqG7O1iQf63I/dkiFDU7wStqF5mx3yNouMVkpjE4QksLL5tAEmvMeF
TAQfMSlGFKUy39MKFwp7gh8PDernGU2y+OWIbvyIymfV2YzpUpVTK8i47PBHPWPG
cZcGP1CTBpano05iX6umaAsV8O+VUICiJkVADF2+yq59K17ucQHw0m+xowexz1Bt
u2TxQejK00fC2COKc7Djg+izQTqZ7/oTmgx+FTkeJjnXC4dbnmruFX/QFC19mBNp
j/cdXz2xBxVioJp5vkcpwN4JOhJ+ObfmzfpLxak3QgvM2yjfmt/xZCb/q7j4xq5g
rkr12T/GfHZLslAs62u32QpHCGcO9xwQU+d1UJz+YUNHioW8FHjNylGdwsJHtXYJ
ye8mUKIklh27r/zQgUWgGfYyr6bB+QjaLT2FoQr3/m0M82msTq82DNbxcUjjD78J
T2oQXvHJBemeg6H/tXqQGmvqgY9MZf3XEfmhiVMz6t0ko8Cp8ogIikXbd8uC7zch
mG1e41XgQLB4g1hmhNFJauUBzNbiGuA9kiyBycBGlm+cIHJnGshms37tVwMNMaZg
/782wv1Qi2NpyDWVQfH3t3ChbkLjkUBUZtEExQmCwotda7dmX8OTGDHA0sFf4J2Z
/VzJGVp7FxMXG5i37tBCTichqZBGvk6Bq8Py8gqVG5oLAhKwqP7tGCCd1UgPoe15
DAOL41+34GXCDaL7Bwje8+uyJ6tJS3Af3Lrs8RlBvECtvajJyyPhiFvyVqHEDF9o
7C8v+Z+FxZPSTaGjDIgMUGAxkgipZwB/zj6QIh//JFKCJEIV/b3EcDaAMroedOPm
Qut1Mx4QV9HVWAMfTxP+rWsa9UoDdJSOwuaspJSvM4w8Jr+58VyCsMo2fUBgl/gc
TT3FFPNNpYYzwkq6ZssFjUnYz9U9fOenMWUPWbeFgEFrNfH64fNvw6Y5zc4Q01bI
0QqwhR0oECwtDedAR0uXHoDmSMNVfR0HkYrhJH4nNtVP1kvzoQDoGPNuTqhrna0q
A0/t1csiUUDSZdlGZHmG0WwQ4iCIjwTV7+IO81N5dbdzhRBlVxD7uTMMbeMCwBJv
u9k06TfOdp2GRwyejEeuwDugL5n2VQOVlLXvuK2EOFlK/lMjoEatLlGXNRfMbyEL
MmPwdy6i7+i3P5hWAj1aQjZFO0cC1Lyv+Z+iRRWLK0V17p9zmeWTw5xXr+CP9ii8
3kR1lremAk0B6HPUQyrAQsGYcuNz+jgNQXYhZfyeytB827yA3DAksKIlenc9Jr/M
srALmL61TdgLFxwhqjWZMyWLMwR/7hAPQADOOzaobSp1nAzp3vcpuRXObZE3Fgp+
ziMfRACpyjssNNLixXweuhdbhon94nu/9Xv+FBase6bWZHhdJfgrXi/qst7zhomJ
dvl9Rb+54r0FfdzB/cZhGytXF3e0U413iPZ+6md6y8iPjSRk+P23xtymAtCcVINy
+2YZXjaVYnN+xGNjIWskXf00vvWNmb4NVOsaH1LkbRZmnoBAM0W/YeuxJZZvlTPA
C9/8KweCEGRxgowzzp/z338CVVQeKDJ8rU0YutCpQytnnd/APC6kNTMVYspsUrU3
fNP2iiSPGBkYbcnMyNDTXPEAO6Z5yogOJIVjnm86kGjIgVtR1Ciw4sDAHR3izHKy
Py0dAJ1WqE4K1d85CNVJSaM6sdny9ZXKC+uvcfrwXEmGR0hwF23BhE3OsfOckCqp
rqHscsP3U1XxlKI5T+EJv+dkFO7eT4RMDeE0SX2faMYxJ7Udzj5Mct5JMJrW8Rtq
zMYPkogpdfRWHbOmB6Im1l0kA3hy3g8gC7CykahMPsmlZM+/hshCABslyzCbagSM
RR1Dtq+/UwsOe6VyBrc2RjWxAVJeJoWDbiC/B2qPq781fH5Rk65dA97TNac3ClZ3
z4LX9YBXGUzEIOTrGxw5yW602b0jHc3DoF50/W3+6cM6qc8+ICOY4UQXb2zePCDN
8f3kAEie9eZGMdyWRuI0tuimx8J3HRakO0g3ljbtNBvT4Ek6DzYYYmuXiGCBGz3N
GJo9ie0AcoBGNWbUbg4ZU/EYsONw2H8z+2z9wxTAe+q+EVCHAIdzc+Am6FdtGTc8
Ru3304R5brNJgxhF+jPa2Mmjm6F72wwjNKa6iEcZ2aKxTeRsaE696VTYIlvIg6+9
X/JHC18nCxtkA/6T2bVN0us/NjFsAFko63DTjL/F+FUMVhdhC4NVHCB4kBIYBCfI
t4Y4YwdnSE3EeuRjEiAUX/7DpNSmElwLrv7DA2FgxMrSMqG6Gmagv9ZbB/UNgVh2
oXT7mtBh2bB+XrMLGzNF3EcUWjHdztYQX2L+arg19SYH8E5tyj2ktjMezdahbGa/
QVcU0CO2amXAaO6+FdodoMgzyr2sdlO9waeW+jeyZGi/bwv35azrFf6MC37iFgj5
BtYTrIQR2a17Ya8T5iWgjL5XuReFWILHgwKJjdYJ+bVTq1RWBbZq6x2g4qbCrMvz
p9IQokmgxTsVN1+KuhZz29wIVPFWUG5lYxJol1+59Q1FGn8ELw64EqAizeBfqfQr
V7sXDAdJEEeh8KPcU4K57IYuNX3liGyH4kcSweoCFYO5ZOztMeAXD3KYTCoO3nSg
yAb6GQdQndeJL5mJLBhNtOHMKvc5Pn+3ouFql4lFDRBl8GHEI/NgX2YE9ZT+e//k
vcVoM0YZldxlzC3oZrppZO2rtfmmBPeXGt2Vv2JG9DLk6l6RR6LyYtlYJXnE2di/
FK7H9ihukjTp+Nha2ERm1NVB6sWuLQ81eJENVKPnX6hwHxY3F0MEHJq42bpN9pzn
ElPlIR4uBVN3YcPYau86V4jXSlzygKeIEP6re1ZS0BM1uEdpMKUg1rwrp73WRocC
k1+cFDEJbhf0XN/XcbhJP8jelGGGDMAUgYeC0UA34RKHLsL7WcXOoVEvcuRdCwSD
5j54FuIBmcfizdCARmt4T25bu2TwEvUeFdShlkmz8DcVUpHKV+sRKECW5BS1qceG
5VohfLRW/7gcVebyVVvuiH7TyYwvyXw91VQf6Hu8jHwXkeIixv8MazV9ltkJeFf1
BHl0hCrKljh8HBkLHwEbENBcr5B9DgJXaLmG4PyTXb6cIxtmTTXBHIc3x97guUQ8
BQLPJmzcfRDa3REFBNP9XQDx102zUcqUzYVxExPj6e/IaeD97A7+OaKqVLSnhh/k
QsQBbUuCuEPhGyuZjItQMfC+Z7P4fcOp15xyAA1qNRorWV4ahviNp1rFRbZuot0e
Wo086xKZNR5yZcqLScuncP0e11OMeebvfKjR0Iu+qXVr7s62oNZfaro+znZYfkk8
RYd95h5RQDdQMZDRbSxbNmTsjYzSsfsvd+mX1aDth74i0cADXkxYI/BHhkkldYom
4tU+EU1z7g1HX37YYrfH2Voi9v51vnqAQH4g+SPUwskPrqYsN4irsyVjld/33yeC
UuY3LTmOI+cVasEKNFj5dQ+RoavO1lWy6PlanjMonM1SkFhIHEKru7re4/8TUN5N
6fL4CHtNfOTSilQVrzBEKJo8y1nFEaVocWla0lIZ3uFrGzF01cLIlfv0z4GfPhx7
PzcHtARZ6u0c5bHJbfBXcwZxj2koIj8sDc+k4AG5FZmRGgfhVDckOBFLD+udp4v4
RU/DYPE+nCMLFdttVznYvD2zOaMNJoT8DaTJ39rs4NKsFyxyA8BXtP9AtU/NcxLg
LF4qrdg9+teLcK3yFYzXT4toOMCOGAiovDaCrfVbS+1A8qygT8kvRESESNC2kTT+
g423qNr/wmmEEjqlz3ECAiyxcwcbd6kXzzRS6rzASsaOCSd0Z3xsmATlKRWavFl/
g9v8LJuKxK1JZgbEmM/94u9zDuVhRRAW11cgLCd11woeTbqKYWr9C9KBdvv31Zjr
gYeyzgETllS6gpr+yBgtRzF9LSEtXD7RSXJ+GnNR9xBVelj3HcyqAG4TAY3oKP2Z
r6vxFnf8Au8yXa86Ln9fJlfxP4lemCKWtnGOouoP9Mvy8c87LMqZEVXsAOMJzxNp
t9nuB1GltSXmtSzZr4khpfFirtqUSsUvmRkwWjzsme7XOzUC5jrz2h4/eGudlsgX
SPlrSICE5BAe0O7bqkIkXrblSA/lvCTLAtVW7fev3XNeXSP3MA+i64k9bDRYmrFE
ZjFsEPuC0gT+jCd1srfLyG7B8E9eO1AVNI+iK71lfbTXQgS7mPF6Kod6qeuvuWrk
FlPbe/lCsnsnC2ggTaVzsNOB8T648pduB4dorr0gCYMMDaQ+4LEje3OMWU0Uu/Qo
qOY9lNTh0WkJ9b8HdzM9POCpqDqH2FLpRvp7YaKqULSGzfZOa+lnt/jyg8EcmKkF
01rhZydATFl1Kxfodb5OcPSMa+V3+a+HRWS91RBlY6cYBB6mzv5OHMOdHYzNtCeE
cpus60sXH4tBpg+EZyucIe7ihhxUx5yeiGq1K118f7T1kmmkjM7Cy/+E+HKNFfZx
UTe26eXGMDSFAJP4qa5hupvUy2yHeNesQAzsH61VgDJQ8Wwd+a6ubM9lBNcQfWJh
OAFuelJ5Yqp8xlEoY/1pp+KzsXYdAugAFeK4lojug5AyXYR2bYIDzS1LXMLEjnmo
5ItIdOibPTwnE6ihyjIvEf9cHkEn85oY6sXKJA8hXKyE3BJZs4tQ5qob1oKzfJUt
FwACvpQCgeR/8VfX7CIhbu/mkwDBObgApYidl5eSsK31+C4C1+XLoyktt8ei4UEy
NH8AQ4aUkPwyYqcUrFjPl373KKw3Twd/o+L5RqwgfNFvEi3RLl18pJKG8SZil3La
5ax2AkG9OW8AQzKeUvE4UEJdAHMN7oPG3xEFFu14QDFo+WNRwxP+NdYGYNUr5kyM
2gxJbUHe8CAzD8p0wNcGYX9hVqSdEcJ01J++vl1b3Qetq/iDo0Qatc4gRWgvy28r
MS7hiHMXgKIfPYDu0lghS8AnF9IRbwFzdSuFvAS2t+YC3EU54BJCBUw9LXIhS6Y8
M/4JNACQ/Kfsd+o2xolkNBIUHglQophmZ2inggIH24BGEdqkZwNFvxm35c7MrZBc
c1nZUdVd3L7U5FpwuT+x3vU7fXh8OsEg0WvP6KHz3VV/8FdzIbsya8f0nz85epOG
twrSapZ4hJZDHvyKZCo4Ox8gnHv99j2uZHEy7+dLVRYQvoDDXv6G+/ndfdG1UsDV
K9x6aAwzcPrP26WI6K7QuRnVP2eSw7VvWsflaSvU2NCyCtu1Emz/lGlHMUHoPnA5
HV8qUfgZt9YXZpBKVZVOAIPaS+RYuIKsJ40bqo44ia2ghYyn49Car7VkaU6vpXe6
BUk749cdAbfBxfYDpeB+p8UoxCZ/6r9AJmA4Iiih7W411XFx0TnoaAj6uWATlppe
+wFdxzkoxCy0MW3efEZjZad9kfsvRZDI74W4K6ffcgYhR46Toa9epCxvqY72UH9Q
P8tDV93LLNWIl5JYkiYJ/w81FjZjnNpKrnfWM1XzDOAuTzLRvcBCDrKWu1srS1Rk
t+vdSChqB0CxVrBQsYqv2sH3gXk+iQsv+/fblIPYrqLSgJpVYEIQeNYAnBdrg8oG
m5W1PvALMDZ8EjpiFmsXYB4z6wqn6NgAwepgv8cTGXQU1KOTP4j23p9DiZ6P6L1l
GVmgikFSODcwSEwK1kGdlBBwJZUUinIMZ0cHbzFmU5kzsQ1EMNhYickw+mGmCT+X
t3gvULtCOqsP8R8T9oJ5eKNnNjIwkzw8cRCaeHstj82Xnbv36CfmI31FKs2DQMzb
B7fP6EU+aHGAj2PpV/cSLediJpGDJSGk7AcBB41n9MocnOiuaFI82WMv10E4jjJk
wSEerJh1jr6nDCuThaSYjfeuGvlGXa0hryNKyV39kHeZvlbyw1OqsVVJRWriJsL4
kYJJuzzkoXDzKpFb0n1HauQMRM3e/ZQiVlCsSAwoMAEJjnUnOWUGW05c1aTZmMvS
zJe5NFsCy+ovcAqRac9tlSEDNwydVFSfi9a3jlXGtih0iiJyBHUsxyPxRZvmY8mo
CPLxYihY9dJrgVQLAKoaSNHNBc0EqUfiMh1y2gukdiL872TerDR5QDn57puzMAAD
7MOIeIfA8TdCM2CTwQZrRAZyjTz3Q5S9BqcZV/C4iNvXLiPTg0NqpCJzEnGertty
WH3czS0mFUKmKH29FBx4oQXCdI8r96XBcJ4mmCp76GLOrhbamcPE5j480nKh3EFv
kulZhQPGd1F/v1cPixbOPJdi5gx0LzYdqsI6D6ZSnf1YBv3BNj2jg9TBNOk7VriE
WBOkiTBPpJZnXv63NhdifEBpwcZJwLfPByCJWjbxH6z2fqSPRqM/Woct7Qu4rUEq
pq9VdS7WWFVHyAHWckxuWulzGJDi3y4dFss0KWq6cyYZ1j+6NbwUV51WkPPjgBTh
ZeE9DDkD4N35tY3r+CXsDkKR8d+z7vXCmf0wpHRWdFdaT2iB1Zv58VekXEYOT/sA
TExt3RRR+6euCE2OoYGI+vivf+YFE/oYMBqdST1nltAw68zVe9DC9Ov3/3TU389L
67sB2TS/GImys7464GHfE6NCoJsvz755AL0vISdzN+xysTyKBE1lPf8nX2GeuFLU
Y/Ma8wi5iaRn0Juccn1f983MUYcLidONru4NiFtYzFFCWxpH0e6KZjtc/ypXjUcH
UZ3ssSqRfRFHqfnvFV8u/N33VE7dk5LfWy+ZF+61wqUGLp9nZJA21spTg4Ti9YOf
QwRhbqbDSli0IVjwFjzbrCp5lbpgg+JhK8bXAOX/+w1kS6D4ojC7QbzCeUW8jIDt
lDjggGGfMF9RXBuNAL8zjElwDf/tW697mgcIZxEVmbOx8nw3YfXnNFsJckj/uGxR
1Uc73xRkYJWT4HlbDgSLH7MLM13SzImV0To+27RyBfi3ze0Hlm/SzeQ1g6EhEqkx
YN9UmaF4HX5Jh1uaZhvjfJ9R+6LzrCjtvQ3oZJifayd6Bspx8xyWNrFn+G4PJ5/I
rQ02/2tAJwRURMPWRmu0sl2BGljEMAMPGQ7SnS5lDUQu/8XwVe+QE5uG+3HaGS2P
Zr9lah6fdH8tKQguOHaFg2rFGI4HyCfL2pyjVhXhSBKpMjL0JgiRykN3KcR4pcID
c3ty5QlHZWxciuSx8zdb8Hit+jK+zJ1hH6EUJJs/cBDe1FpZjgoNhyiDKtyjb3F8
zJ91pUXXTOPWzMFgtK7/pI/PhsyUQvTqDzHsX1jvf2+3wBdXL2TmpyKgShCnRxLy
YmIlL2T8Burju4Y1zlozjSR9ulAFXxJmF5yNs3H48r8TAsHHE92AeNJQRO3aUpVC
nSgGVfOmTJj9GjM46QS35ahlnkuOFhU11HAJoGSk0WeVqToq1AgI9ohCVi/LHSXR
hYOIJZLy9fAN8KfLoaD9ImUV3Emy27Dq25SY/ywryAubPbs0kQhPw4MvqlUXWhmv
ZzK4yBhx0BQFPBMcHFGnbAzkNSESDnL3POOpEBl236N7VWcEtEEDe7F+J8d0cfhd
24uYZacYiCaM578sP7bJznhNuzbKa4KSZ9CMdU71F6nNnfJHqdaYdUSIbuzL0NA9
QqUeEdYjA8Ex+rqi3kTeilOjrKTz7bZ4lvdwjZW8gEsPPlPVeRZBFVv+Ve5c5yc2
54yhS9PJEpDqPAYxWr7Cyrlex40pDzS06XzCgaEwUU1RppgOKZUEDvssAzVVQSjU
ht2A7rPe8TOWNU/lKkWECiYwjviRgh7Mv4ERZB0C0U8U+6UHZKyl/VqX0B2Zi380
lE4gzWJjjgsTcq5/V42OGu1t2O91cWyIRzkRu26i6y3oa8iKw3CMpMFGw9+E8nUx
aBnmDl/tVl/JMZ8M8ZWLVu13kjhe/08YVRUrnjjKT9S68G+CYq+MLbh8PzKuzZ1t
al9VioE0tUnARGypDXZ4C46oJWblKSH0hMKBiB2+38XNkDI7eYc+4R1QHwVtHu0g
6t6j64wBJxvtyywvpCp5MqG+/nb/ItcERtXgfmL7F17fmPJfP31RJoXI6LiFHs5F
JzL8Y1aDP14Odep9aI5Dm0YgxQZieZQ+hfJ4H5EEJNRXU6aDcRuUkFESkQEH9wdc
+UT6skGFNpBdlXygDfbe+CKJN3VD+3f1uOQ/6NgMXNTppwr8CFflee+CzXYI3s6A
HmRi/8Yjc1waKyEsYnzyVHKiq+GYfwVnJ9zEOdroAwBU1PiOm6npILlxdRvueN3g
Ncwq4tleMy90XTSefkZvt1yAyPruthaWOzWYVt2TzoiN8hoZdtZ5cVI6YcDTa27V
kv+cZIKKZyoOnRy72YVoCMwqEeuDG1jTDAL2d3a9juWh77nTHTFApqAw6JlP+/Lg
05IpDcMyeDWu1xqqWA+BnLAl2B2T0yEoexzH6tj0bvkrNWQnh9TiV/Y22+prF34M
nNQWZHDnOj5MDXj3obXflVnGkAiUjg+FCegMLbENN0HNJ0hQhU3/9tWYylJ3dUkx
8ECuSTpJajWBtuUH9mOe+aMgf1Ux5eqnehwoJOMtLvVhfQn4xbnuFdO066Rb5B4e
Zv+sOamIuXIwy5o3OLxjtTTm09uK1QHPLz/z1n8Vkouyd9GdO/x6fS/Pe+Vlw0VS
isXH2WRRTW8PFZkViGxBU9nlKuPeYXIjP46St15BnxIRzK2ks6H5VrkAByK3xKBn
8JTYmxIhJLAalehEg5LPhoJ/pQ4jOlzre/Hrm6FBRzQLVGilXTl5PzsuQiNcWHv1
RMDqL1SJMepJUwkGOi1AH3lOahzZRwqLmxPg5mtqkj6vktOVreKht5p5QYjiUKti
cZtghh+9pYsW+PjCTLWieRr2KfQr5mlo+SOy+6uvWMPXmT4gCGppI+hMZHU12H9+
0d/tsYWPa0j1LKkG6Ncn7HVdDb6gpdmDnvDlErzYN1IufUpAxjCcG/TCisPk45nB
NsLRDwfpwnPVLBmzVKPMNwWpfBr7Y+kEynnc4SzY7C9BPR7g8DzfNe038USYRYV0
eKgdTfWSEnMv/4gnfahF4e+E5a2wXfF+6rDASzwzOyaoB5Bs1wIsFpGhOmfz8O0S
YTP7PED9hM1RBN98EchycdmqFIEQ+ndTkKrW3KwfSvyZU0tFOUiHx3tJnvNdBoS9
CxonqgKpBOYsrRud5JocaqL7sxfr6kk1bSlxen+0uWMV+eip92DVV/6DnSxQ0vn5
OFCzS9xuWC47El7kiHNfLS+iSY/WI5i3WJyfufZXEqc0JIFjVOYhLYcMe8POLlVA
E4FXULNFd8zKkPYRmGYi6VQMcOTosol3DzCeSHKcLauRqUA3+J8mXGOZ/GGzIIZ/
BJqSDMV8ozIkMA/HeqwM7aySkGifEmXLU7E5DBA8M89x+O+RtJBwDo+3fCsTqV6B
qf+9PFnsn9LwqsIaXS71T2H6hkxNJnpDV1KRs57dz1/D3cwl8iHHyoKLQNrZuoI/
A5KSzUnJXF6qA6Rwpbt11K0LUaSgLI7n6R5h3BuXIQeBasF0S/0rGA7UL8f1/FIV
EdlZLrgM6NdBwjr8DAdt/MhO9zcLHtX3H1+rgPglZIRSH1rVXVj8Ii8ihtahvH0O
/57Sy6HmzbTIe4FsRCLqv80lzLIs2KWts39CEQz9tWgggh/mQecoF42+/34mWW17
MTLOudM61sfFAkjlorYOjEVNUJ+0GxIq4vSofNs6J2pX/Ke78OtM0zJw8fD5V1dQ
JusAo0Jq1811GDDoHqhu395Bkpw6/2K8THTMaaswq0rpZTGeraJMxC20wcp1JP/R
U3qKsVS2tOFaRHElJZSiyed1LOjjUhW6zY0o3LDY2QBxBbWjmJzaGoxWK6NAkmfG
1IFZU30gzHjeSu1qfeXP5q0GMKFkfGYFW+bLg65gbQc8Zx1UIHmDfz6086J5roEt
zXRaLz69RkcQBPx5lPzPsouYuA7QOD+VrxVMQEa7Yh27weceGaGGRu5sT+c6jP2Z
T5Q6nXzaYaV1sJ2ov81LeSgjDrmuHCY/FdmDUtb/K18vZCkI5UgcS8gJfCk0IZVa
Vy6z/CFz3h5RNGk7GkZxsxki0rElSTUPzdve0rxD0SOav/0lmri7Hx2+uZt0+kPO
/lnLCKAImzTTwZLUjiZ+MRFASvGC4eYbQrCzVQylAODRqrCCDNETQpjlhHnAROrW
W+VJKE4Sa2Ox/LJHs7futAmFPsXyy0ptT4NI/1Wcc2O3LtPjWIPFttjh+qiS94dY
JapAvk/v/fG3UIhKBzEBMxlSHfUZFTBffAVMZQVJIRm0LS3XpVxRJdew455zTVZQ
FUUkMHgBjg4sS0n6G1rs4iviLM35Uk555muqJ5soKFQiQMubn4WbZs98ePkSFa9D
CJpZacjSwQl+QmFNB6/Ruu32SEW8RhI71EzUa26Dpv3223JDnv3rq3vrw9HR6Mos
cWrZWfKfyumzpFf7lWChc/rLznreTyXaGqEyB6ley3xEgaR/Lc3GfU9jkTZgvwwD
VqI5Ne2So40oOB1oF8udO02560YPG+b5+rYcx9dLOoXbFBNPJK0JX1FbasXs8DgU
rJKkVNUa2J0oC6kgqU6mCaw677x9Q38k7P7k/YontawRs2EQEuv5F+XBMguqWCyv
dRLCfMXuUt4aPgrq4TCCfcdAXCo3FZC8aniXtjIyF3W3guAjlU14pYUgLkpQbV9d
TeGq9qc7ybcz1HiWJLr5ywNe10bfbYKhjr54sVnSLRvHCRBVukYvYolv02DaGnjw
A7mV78vQWbd1XvmWVvUnyyNZSpZdNVRHYeoOJaKAtU+UoSwK0ZMn5fLe00hRv/gh
qeBjNJqT6C8Yb1+mkBjVgm0pTfDYgvnoZWcvRN8xTrTHAV3yzVAnChdD468g4bxI
oL10CyrAloMkXpKROwxfb0fgU04pHUVhbOO4nSaHNDiJTYW0pYfx2DqGLVzv1yFv
lPe90FwCOVNECiFdTLrl3fmF3ovoV1ra9P6ElQtKRCujsK8S1Vg11Oe7/hVvOloH
fGk9qnepZJxFJJP55NgF1OHcD+rZnr+7aFvliwwcBrzFIuLK3BvD03h4jKO7u+iU
Btvezlxh1Ru1MS1fVs3wQfqOQpTR3M52lhYpNzEp18HBCVxsSQAwBx99Z4roQiuB
lCM8pEYm2ilTJsLh6xNhngykQzRDTMGPdnRuFOwRsllL2Lu8h4+tlnHe6WhtL2An
pFE9XFoSmpKQbAV+uzg2ryx2wZf7T4X8BXes+x2iZFE2WHf2HIBmSyW0O/l2P/s5
PgRxGJW5bYleRiMA9c4NVf5G7X+c423zMr6KH9PbS5pmSxNCE2FNRy+gXQdJnST2
xsa5viOot3AO07ZUfiEE5AHIOfkcHsTJrdOJpB/AUeKG8zgS9YYxHtBHLVFd/S83
Rg019YA7qgYbhJ9ucSmHnM73S9z/6KBM6ff77+d/liCnZf7gpq268xsDIytSQP6u
PiJLa+r75JPC3byDBK8rtH5teUrD45axrFVnsEWXtAgGrf+PW2d3nh/rHSYRub7h
70YN7VHYUU4guAm8TrxP1bKDX8NwW/9Fm3LhDBMwwQxuhH/63VktKEiXQLq23hOs
XauCgObA1k5SvYp3zaibVGk8myb5lJ8GiSvj4drKqnrSOSv3hudTaC9KlSbQ2xWp
sHYkFHJ/8R0xMOceGxd2dG3Lvmp59ph5YPDowojNmJ8zUxNnb7aRjpQlO++/P44j
xDKFZfguzd+iFS0MIKWWiUzcc7zE4/Iz7ca5whKwWjc+zwJ9AqHEz7JkWWH1/gl5
t5wrey5+e9yG4M37wVwu8fL+Ou7T+arkmEtMU8Tfb+oieGrNMgmjL41uhVn9i7AO
mwR1CA6ex3bT6di/wFe4DHgJ4yzH8z93VYkzmSx/zsSqGa74aGZo/7U7ADXQJxdW
ERO/TMlJf4gVTH2DSJEy/4eBI+IS5lzT3uuc7qgzDgW9zG0ame+hPMXBQ4lM3ruI
1lvLzl2RqDnaWyxiVamXUNFCRtYZz/r5ceU9l+TvmzTlvUMDSCsJcW9RVC0hLAq9
59U2ADgxkkbjyzjwisKwVZoCDu9XK0YixDQ4WwDK9bAviYXxz/iDr70ox/ez/crt
RRFfYSIK9IDyvUJJHGqBIZK5ACu8HjOx/G3lWWSOkCbivpJr0Fv0VQfNZ2uWiVQC
+Qug4GjHz4KmgtpDWVxCIDdkn7gsSJ94+gV2+UdkcomUO2Y0ZexOMvwHqW13fW+H
apyui9d6Hy+GwnCfR8LchmqoM+dt0QThLbwsa9gPVVnuL5tZSO7SDpmavsjGvcXz
P+NTUdh16waATFvRDR8ttbG0LiBcnCRjv8z02hb5q5KhCM/to0xoIeWDZw4iN5mW
XJXqV4YxzpOJfZRG29nYv77RzM0BUjwuS/aMdUsGEGpTW9ONrBnlXCzJXTaLyko+
1vkb3V8Lat4trRMx7yKKP7hNM5rhxploEY+i5PtvnMU8HkeZQhx1qM4hdK3MXW+g
WphVh0TMm5i6dgOHUAl7IYdkH2UELHo0ePO58MxwJj9nOV5rLp3/ejpctYAPVyx1
9G96URXOUizFpQVI4GjIn5h+7qHTeuAZ9xmrdQWqmhQfDsgCVimR1GJSevmYLheD
fsMCWhvbCBhw1IE/aW1SOTt86uEL2h45mURRaV96WLdyIVoz5cmlM5yotAwk9dhv
B5XYc/y8PwOoM1uaae/JO/JGwT8da1eG91cENQd/hjZ7HkO2+KChp4I7XPLSWw3i
pMWK9EegYgQRHUtDrAi+kqz0Eaj3zYs1hPn+81olg3Th04Zo+6F7kXUMEHIuubGA
xAm2ScjAUUvaeJCST4/8VvoZRgOdVx57MnsmLlNM2mhUmtYAfpOp13I2XUbc4T3U
ZsPc0THe0MeCbv6TbXhjuCQXGDzkKflzYGEMDt7K2GbprtDV4myBzerOUwjlVYxL
61pwmNcDKcN8te0o/sLzg1DYxiXuPsZyU2+rZwbwR7zshjOUVM7b1FNyoJqxJxMS
RdZ7eaJ8NSHv0S4ucSCNduomndReiHUYj7kCH2mKsXqHx+uz3l3ZACtS39X8Aqaq
vRXdFz81PSCyCgT35QoFG5+o5wmI8UJLgY8PawUjeKexfS+xyBlEle6TncJmfn+7
kkq2/hv59wUoyxeGvlm4S9j1a1tGx6p5qY9bvWkzsmTlRcmIcN5Eyh04Xf+Ptd/y
qarnCZkrzoQIq09gJ4z+/KfdDeUtJo3Yu+RfhhqY2yLu1q8zXxMBCuWn09EXdWvr
PJs8lR7abBnz3xuNe/TD6emTivxJJJBxUqP7BUmBVPTltW/U19ZU6UHJodKs3rMy
Q9FYPNFMxVfi8MgVOo3iHW0zmL3HrLedBnoLaLuEmb1pjnaZpRtMBR1srWSJeSp1
9fYZ6e1t5ZC0b9LFnnJToQPWODR9zMggCKAk3RTd/9JrwadszYMI9xrwuX2AM+nJ
736XdImCSP4MLH9TVSWlVxiukqRwKqkWYf10WT89tXd21nomLgGyFSLYW6+9+gRZ
M5coRAjC3ZkhLQYEp93pzksDk74suKP3t7o0QAXHln2iL2dhHOV48Q6UE7rR+cgz
9JtEtBNAdtSWstrpt00/VWZSYmywwyKOuC7xtzbibx9XjsVvLUPSBSlxiMBQ3diB
D0KBoH5qTMEmNmXPgjTbQqOUAyryyPpX9C4zmD7NYbL4c88spI22HuiF5xtG3MQI
ZJCInXPY8NZkq4edMK6Mk3Znlniz9mvalbffyAkSdNU/INEi1Dynrd0gWsNwApl7
W7K7HTV0jVcw8yd2+EtC3Vw9/ktljnPPUvR7NkkU/qdWaNUB4VPA9cSePqj2X0vt
Uo21GUA2daStWzGN5eP11uWL67iGvVpFqh77ZI3m0gZHMyhUzlluZSZFEEu6VS+s
7Mvmh6BO5d6rKKWuZSKxN0TLEIYV1K+hdqC/63O7RPl8MISdob5klFbGNr84r/EY
NdN48VFTrpKAcFsuEDhUycC025mokrN6rduPi/H35EEhTPYEP7NiOhOMrYj2+C3S
lRuXPVDjY97IRof7NslKdhm+u9KG5+m0Xwr4VdZeXd4+tsr7wZsklLkqldJYBjS4
BMg3wDw0ShMiZPcxkwpfznWaai+USHK+quYAJgmqKJe6vPZK27ZN4VzJqLYU3naF
6yW0FCMIel8sC1XaR4rzwLnj9k2nSJxBuU6Vg/fjssiI3Nh7cX/WdcG5swZm8/nr
KL9ZPvNe/4UHNEauGQ/wAhhr+Ehkv8732C4N1c+VOpWDOmOtzEigMIO+o2wu/JMV
RIffhJSX9M14AufEhx+bCvwTA/TdiQz7KEUOVIa/pqZ21xhyQTQolXk0gjOZTgca
5DVENSWCFFfOF6hl5dG2nGc2+1QF1zGrbq9FU0CTiIGAd5/pygx418jP6RJfY5Zg
p/Q5NwiuQgmIWnOKWXPA2M3xOAsoX3pa0vQK1WJOpV54oQfLMSPkIem9csWyznT/
SycKfV4NLZum7FDjC8Mhh5sQoiKrGZTur57i0vGPqDKcOdr2dXDLIus3A4azTZYA
TF48arNq0AZeWHszu6UPHiNspSgkH5F2lYhXMIh1urQHV0cnGwtuAVSd+arkgF3P
k6AKVIVaVHXEtQs+Jb+jLsGz60duf+18M66qCOrryKve32bLhM6RRTRFS/Lc6mkS
klMHMHyOHL7PHEAnwl2tHgGLU3VWExZqSNvPNU65fUkZGd5TFzT+Q8k7/+ui75Fi
RofYU8EZO0zPaSTU42NGwMHLFLKNyOhljDw2t2ysrW9ddAMse+qwGNnNtTzZgYbT
kM27HybteSYQ889tK75GDcYTD5tFXGbt6QiVKskoFXL0WvCEVVaw97nA5B5TQgTP
ZDjfkQ8Qp5OvJ5gombXIk/T+aWzv6iPcl0bCdZzv2fLFFhCrSY684Oo4VvM8E1jo
vvxpbYKLyN+IpKfwgdQNdpZKEGAXg+mgZ41y+Tq8cMYIzG8qjhM2WrgR9NMVF8I6
Quppui91bD8o6MJBfZunvW4YKJgWRPCeKQJWyL9EpwBODV3g+D2bSboO9NlUo8Cv
OoxcPNxYPZnAntF7XkNAv6CA/taQC0mPCB0yacaCCpbwA46h2t/GpDkgfJRn9fbK
56FqA17GTcMkIEkxbIAe66UyxJvDQdzAb8h2goZEg4ofgDOEvgeiZjDUBrTTDPz6
PsJJbIeZhjHy+ylfHWm9gqorFDtAH9yBP6K1vMk3JWHDNHqiU9+TcWnIx7odW6U8
msJAuK6LjIzRD7SnWobpwemtfh6I6OT8vEMQfO4VPpN5QyICiqHBEgdvI7jYzkvT
VBCud2PNYCczNXg4qTmmQV9INg0ifGcQ9pO1FjkeJY0OeDP4JwWP8XPkz6wtHpxH
aau2meEG2ZTxlY64rhOhcHyrj7eN7S3b9GKCZBzD+/FNFGLr/YxBsYRjqmd1506V
kj3kzoxnQylU9zz8pnjgnNUFd09Vlo1wcO1CvpK5nhQ9so1BfySU/epWVwqCcHuY
F/pMnHBKQLVl7wnT1QNoJfIKWYjy6r6pKk+owrZ7ohNnsrTbzjbb+ugtvaTiOGl7
t6t59uSQg8IsK/gFl+dfcoEgUf2hVSqbSQGlSTi8nxJIveg6Hw9c7YMBgRJ6bCAb
Nn4gwNInTKno0hx2B8WgwfTG9osiw7olvrD/+qRXG2ajL38X0bFYD9hBAmvuQxdr
804X4RmUCU/+AxtQXmQhk1mHqER4pmjZ9O/lFb27bg04PgfCni1W/pzH+xZkTBmg
q3vQ+DSDnw286So6U5mqiOLzNNxFoYwRshVAeCcbytCNqfz1ungnvsNes2V2I3dU
j3ypyMKNDHeepuoS7TcFbRKqfkn5OAaXDGOpNG14HPmmmflWekdbKk8O7xMCJiOQ
zug5obOspB9QMXJ4EVyuQRm1zKfgvdhnFcsxD6QAzH6ICbKcPsU3zNF+THJi6b/p
i9LUS44BqNJflhBhUbX+Wf0yHfjHiWnY2ENPt0bCwzjBd5sU0clyO09cD+GMnBHp
fkQLq5FVKs87PP7yrsO847DJHIp3sPaz9uH8FnEhQxVlGpbd4YSPe/5JX2cS1Ir8
Dcoq1m3y5cqsX2C8+N5GWb+cEW5KnZeHvr2pZe8Gyat1eir+h97O6ncWwQuyaqML
I53WurbKsQmBzcSsw+VkyNsiUCNivT7UZKZFtxcgrP6VnJIoV/YKv9l0VeZhIsHX
UU2p7iFYzuMkIbYHEeglgMiLYWeIateUhjhATOP5WYJd/mDlVbZv8vCBbJ01gHub
q6E9/iNmkLyckWBVxz0JIHccfQ8cujY2fF4U5P3YVubSzEuDA7ADYS4vBsKv9daa
Hg//8SCfUVVBI5HJCHUIzRHYyQchl0wNsTXzPa+ODiqXYFYR7E0CAdA/6ZOLD2Oy
FeuHCAxONrP6j4SX8m/lc6fsbyA46Hy9GIAR4PRcbEAwskrAcAgjhcWoB30kApMS
LNJcncc1zyeUojBK4JnIZrqe7FqUv6sSOFT0DN5gH4WMLn7n1KP13HvGkNfQQRDx
R6pTX9EwynVkBWoryJUiEYiZCW8jsFSE9fbJbY3gRqUBW6odDBQwn20+7xkjtrxz
h3oziW1svf76uSCFiGbPUx04zaVsgB7U6dIRH9AJtI/cRhgCndgdssDEGn58mYz+
wQTMvS+lTEjWrutbTi0mMMLkLzkC9NeaJK7EKMD2H+NTT0I0vZ8/hB8Ywb9xnV/3
DT3i5NtxiG8MuF/B5UFpgKhsiecUI1l48wFTuKsTWj8L0I5vjb/cL+IpV4CyjG6d
p0mSUKlOJ2hwdkaSFvarRtRwTTn8x7WNkds7C/hbGF7Z8J0Epla/R3OfeF4PiSRA
KSQsrlzgqQi8fviDGDVDLeSe2fYp6Kgrx0C47J7bmxddqYBJ980OSMsrRZ0p4bmQ
Ma9SsyIPmr2plqtRM1EDeSM15F2x1+Q9o6IuZNLBcVqSRGwDwt7XySjqovIgMm3P
L7L9NoSTraKaRc3BBBmoJnGygBvk07B//7P16b8z2Xp4GF705DF0sXwYC9rze+Lg
cjkx56iGfiPfWLxQ0MGMsVSI7xJZYP/ctME3zn6EjQqKZ5YJPAQNc5phg90OFtdN
qaV3iv5rF0mMqR29cMNq5mg8L4/jYJQrDSUdkwN5pUvdozfXo1pRgExDc/8HXpxl
1eGjeeTX+kRsor6LRUWwi1Csdx9xtkuiSvb8uLZ9GaKfqwELx8+lFK54C2mLXebV
EYglUi0W6ZiiJyOd+vGcXvtjhzMuDygcotPg9/D5wjx7+AanKcIBKAnXI5bZD4gw
XDhP+F0/unQMnC+b/IAfNaEJqHm21g9oB4xyQUqeqUx9jT9Uz7Zkcgk9RasSGFFb
sQ3CsAORuCGm05t2rwcDyqyMVvBfA1/I0mFH1UhJqhpO+Bo3VEEUcXo5ih3udbaj
1L0THbLidwjDFb4ijHcVYfACSmyaLu+xg50cOObh4O6X/qy1UZOe0v5cWFK92ywf
GLQU+fhTWhAh410mcvbsODqobkYkB7lZvgySQ5dG+djWmeihnNZq0bYQ4FXlHEot
isnv64jnCJ48GnibFGTSs7t4NZ8sF+G9l5RL328n10/YwYc28t2IqFmtJVK7YToe
XIjB1wUeZHGb7hRjtM/4wrC2aydJNTA5WK2TDXXZDOiKIYiehZHzGMvxCNtFXZvD
2kIYSIVIpauNwzXqCQhMQf5rVysq0uxd5YrSy7xJDKE3bZMcwY+IzWjwbsZQpHxO
dCn2EuM/EwD9W7B8f81CD2sM1SlycVx5QwBWB1Jiiw4B7BvKeVysa4AiEkaswotD
PzI2gmVWmmeTlVN+5sukWJfJ8lh9XnzYvv3++oRyQ6eXxcfaCkuZL9nqlDue5dSU
/x2OzaADaDOiSRozZeBhW7QlO7NZe/JkPy2d4CFz2GaqushbKTuUVtoydBhZCLCI
++iQbe/jAaYlXWbm1EhOyuv3AYas3KiXmdzhxpRAB8q+iOSMMBwGtJpCAEe2/u+L
yYJ2i1PBdttLTvJRraNnYAR2189wkRthpQCoNuR3aDzE3v2b92yGKuE5RnBgh/E6
M0X3WM+mao1hiVfFSlDvtNOTxqbJko7EYzCiID4SwIYaCjHmtacgbZZZiu53mkiL
OUPFF1jsyPVJIGtceiUNXgGivd8nXBIjdftdAeVPoZJtMNfOeTtlBXb/Y35RGQIZ
V5prB03B0u0EOpJjF2m1xNCKm6HvGQuWBCcpU2ezrJiwged0OtWy/UPgMlWr0v2O
gKn7MTsDsVrPckdvUv/tNpz4RDjU6pOQjxEl0+CTUK7c9O+JlVr3W8HzKLYEfsE/
lNHso8eu1GvVuk8OYtXQQNFvrQ7VClYdil+wtphtWyE/SwpB2AcmyVKY6Wm0OHiu
rP3mZM+xxbK0w9Wl8gX5ngNtUZFlzF/bZj9eFA38KFPjp9Cv8z3vLQYTbvPvQoUz
sXNG2s4GqAcq1so1dtGj3hNdTOAsb/nJFoEqbASXNTmHbvQs91KYo7AxO8734Phm
iGziSODOgx/LjzL9kgPBh+bI6HAT9a4U7EQFY2Crq3nmmwk1PoJFrVFyIDgxZjWC
yKojxCGUkFJD+Qy5DMSopkoXFd+qm3lbKv+7MlDbXeGSJDSwDIscKl/6WylkLyjR
RSVnKr5SaxAOaNvw09jVW69TxJh3JceIvHNdjMROI7nM5RcTLVLGwlmq+PyS79c3
pSZSoXpHZ0VBNwNSW269b2HqdjFOIKxKvAFPbb13fpj9JyjR0QcD3JyIKHDnm1pp
WTJBMQokKsEkUTWNeeXkWQOuFY5m2XmvvbAePIUlEue7QhvzvE8odbWikLS/KgSN
qJTws0+Tp6V/V2bP5zFAKtkqSDuDlgW2hAtVHoGwQ1KPid8CgpRWD/rfLZHm66r/
Cy/OtMmOGF7uQgbpNDW6tEmD0pdHSB5pkMXAWgsixSOusSxoRhdOHLMpmi3NfqLg
PQiWk0HxtXYpyQFpASwTf4vXRWx8z4rRDQLvFYCtfaEJsovLDMhOjnscFx+Rxbxc
w5Y5I0x1CqBWmvU2YVsrGoRNMYkTdiFELWX7cYXFe2mXEjRfC+xAtW8FP4DI318f
rsvHH/gQqOgkdHqTmrEJe4Vb3mO2sKcaL3Hi0DHpo8tCvSC6/gB9gWPWZCsLboKB
PdS1OWA8lg8GfcKDuJ7SbtL3ZlYEzQDXUNaDW7yGkQZeETpOMNi5WPWKW5HN73O/
P/5VRZGxGSJ3wRyqcbmhsHk5kE2ExQ2sxDVND7/hPMRnYfaLg7yFx7nm87pNxenp
KeEAg/FtqxtJT3kFRvtulev7O0XM8knjeA+NAEymmAhJd+WNlHoN8f6x9jNcRVQr
PHxtUk7GifLA/HKOQW07DDh1aWSJk7zUz9rwvv8fjtd99OB2/aDf5bC/T6tbOfT+
eO3OzNH6wI2upz9byKFBxTNXXNAUItqyXKvV0zHR7RxPBBTqVhKpqyWwBT/XcFjA
l9nSfCzv7jMmZQ4Ika1qx8zhRcj43t/iT0cUF9NUG5vQlSG9w4N8Gr9gjML5jgyY
evWHUk02cv+ObopnNOwHtIvIg9dc5glNIN3mSStuIeE3m+7ledYsMci2+uczWnMi
PLD8gCDpEysl7AbOpccru7rIoh0XRTm4ux79Y5odell4qWrKd8hrh2KdRW47Vsgb
e4soyuT5TXk1oCrRQZEKTaYw5220c1X63fL3ehGRiNCCd7EqK6UTBgc8zd0gHA24
X3d3ijHAtCa3OE77RAtiOjd7SfATiGE3bRoTzztU2B8BK3gDuVLOa7h+pXs3lMPK
/s+laEnJwd0ECKEjKIvKtUNqpyTMNyW1r/qvXM448N+GBrfefBB0oiGSNJvsNdZ+
W3SxUOgjYf/E7H7e/JRCTMW4wgeWoKiP+edg3pefdQvXo8iXyw9cax/G5Naynxp6
lmxa1OUwODpPpJQzNkg8SFUCtgOHBmwADxgeU7XRvFWweAatzxOBAEwR8PiwgmW0
+GwOjZZSyw+o4tyDDPOYNzLrb1lWHlQZPApW/JboxZkI0sECVZ4mO1l7gS11dRK9
iBRz7W9qUd/jeNQ5dXH2mDGP3ROzljD5llHDnSGzdA9Z9XBY3HsiARld4K7ffj5o
s3QD0LSVl6hNuC2xKFPg7rnmsFAYBQExcnjc0MGBd3dfsST75h3wpLo1DM5SrFrI
xTQgXaXek2GFLixIb4ZDUcstWJTfispllKGuxh0Tj7yueP92nuIf5NwxxTuAL9+I
Q/4ECnRy6OnbwXcCh4OOqIh8kJAfoyvZEzH/daHUu+gxs5o1NcLnqrXsZcIiFDVj
st0kenhHvix0d78xEkuv32o0tzWjy8AC/yjIreRmgyHn003SKLJ+Q9ktNaZI9ByJ
T2ew5FUbDEaurTM/pHR3egs0PP/uZOFfeRoCy56rkRkshsQ/QqVW1F0BRBjBWqp0
Go9BoDCSJWe63G3hJrUEzBSkNp+eZKE80kDtUo3D3ThdNCBqzakGur2+p1BDT65R
6lPo+i7AWBbX4Ms2tek6ej2l/ntQd8bOqI1XT4wyHNh7Imhkx38ojdcA9jnACd2E
Jq8dTmlJwaW7wjvSjGk9vZR1CC+0DEnEQECxGhy6kicFaIB5/HgDxa2v6nsZs5RU
bcrAi1uAqhUwSYPMjksol2RAciuCqzRBXr/WI0CJ5eLZHoNGV1vtL8/UZ9k6IEIe
x+6q0t75b0PY5+nXRhQ8gJoKMH73zRrV3BmloZG++LAeF1K6/d90bv8jwxccyXE8
LjYZAi5oVGifX99Nci3Pp4hs785SsaPGJPPYlwGP00fW+iyTUcpGVfv/Zk4ydJmA
Vcw2Uy1/xude5qobvpzovw==
`pragma protect end_protected
