// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
WtA6OiYP4fw93Ni8rcODWBW3/1isCH7JSu5D+D45ZBeTs3A+CUHxHNJdz+xhMV40PoXeh3oxJYBD
bDKl3AdRujLKoSXeVxNipIEkOWOxjwojVKL/K4DbyAmGBh0emWb3qI+egB8Hx8uEtrL8OgmkqYKb
QGGslOqROKJSw2Itg9TkZCNs2bOphos8rP6UJz9HL88astURgb1awN+KCR7qVopYFHwWuG1i6Id6
6wsmBjfLHQkRNQF2hoWO7m+kYP9qDQyPSgZ7ddM90Ww/dHq/LLyEqc+B+a5RkZFFPNIyU2h5lmm3
1uzhTTyBE2yzLQCWlmPRP9se2w95kWjPcxjuAw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 37136)
0ZJkoNMepy2Ba4Br7EgmiAiaJjIpQMPWAasOYrxZmAHbsxEPo9scF4XyBnm3qTII7kB8qi3HcGKg
niDybzWGFJKgU9VehesAG3l8cXdw7ugETeBbkAgQuk1MqDOe43yJdImw9tSfmZU/JpYZpHt22/Yl
ZIus00yjNU/FX4j8PKtv7dVP/pHgO2xE/TzvZx/Bvz9DrBk7IZY90/ba/3gzGZkj2wFbcLkBnkSn
zFpUjIJltZbgHOc5ODdzDN8FFs7P6UJFehoIjx/+935Uk/RVBoaYjgraHeE11223ziflkvedYY0a
CfbXbgUgpFUhpFSszORPHu3CBAQsKhNs8Yj2Ymrce6T3tomyehH+fCKA2Q0F1STzgWSH/TXd0CYp
Nor2ZqrgYOa0jgh/sLR+wQB8dQYfEp9ggGDGl9KkI4AjBT6VH9t1d1glLLBkPCNKYsZcravVl5JT
mQFrRe1cg78s8GvydAgyQqvFh8vEBwd9uNcOxk05vq4L7dQEmCI0gIJL2YsbiCX0DZm5uZ8+fuJP
A/j0pQiJeOTAjVm+cud09YbbXNMulN++fBKqXjDq2x/mN/B0fvDHDOEsv7YNVgwQJJP0D17chto1
g+ewQuMTGQNLWe3J54KvBqsv6rTgfYfzhB3gfNLyWsgl1PvTYlsqE/oemV6HKAZd7v1W2TXVk5X/
xzlezSLlPH2YZVbgmaGO5BAi7xVsGNvfoEPvvA2Zc8fGrICZSzH/rXei9xR5l1AyYX3f3Lr44GWL
p8Ek6P3c5LLjEUltl4yHJ47RY+IFubSJR7ZZ5NFjNZayUhotwdHQihXXcbkKG0ruaM3Qbso9CIyu
zXY0h/vmEh0IfcmJEFwMUeH2dayEt3aDQaIEf1Y+Uz4hYaCYUkhERbQVAMJxOE6GhH+s6NOrYqHG
sefhB/vcseM72OI/1luVWDfOKgOPNX2ZpBO3H0fcB1E0g/hqUWtkKUfoHKBMsxM1Dsy3Bv9/LZrh
6GVpbbXAHQG0CJbf/ObcbWHkn6LqiK/BSjZAyAohrpCVm90dgHYy7wAtlIyxOzxTyMrzJXVw/L93
PKp4/W0O5JU5mbzyavVmlvrY66+59jKYsxQ+eR+cSMaeuNIL8LrFFmgjw3D1GiULFd/0V8wbGX9m
N9POMA9Z3lf5RHXkz++h8Bbn6AEUtrLbyb4d1onSixLiZgha/NyL2PDqTncYdCOt7CgpKHdezn64
IEK0CrnqBvAVX/Ed89tmaTq/73BY8DlvK+t9w2J/xIxhDzhJ/O+BwlkhuC/CLXN6Tgi/kDAS4tdo
RTV4vVwqVcgttRk6k/MaU79KmJbK6HGqAsu+LUGs4et9t1fu5JzaSUimxTNI320ZaatGunRlldfn
3F8c5qv19/0+9q1ZWUVREs35mKVf6a71DdsmBJtO9aWxrj8Ktb30GuXtsT5uZyyTazoBQp/3GtC7
2Ae7PF3nWa5iMExEjWRUfOGBtaWFutY6qWJ7tjFTz+N7FnPyls6g9+uOLH1ykW0LA5k/QS+MF/Kh
o3Mp+/3Odq2KCm3/wjepY50QRH86sXemA7VJPAtLHnoLGs5ecGKwrPPkc3+Z31125b0ISlvN4FgU
1JmbwnBq2i5wiIiFsv0zr/V2aDwksO8iiIFqe3dAB/jDWoiyr3JBAWjw+E51DpihfHHw9eZHGzrW
rSLwObjP8We3TWytR3elkqTnYz4b7h34meQdO7c1Y/L6ePQuyFaDuIpMdQ9vL87dKikHls+9H6NU
4Qd4uW1B3NGsCD7r89U+qELOPdqZv2lnL51xbOJIxJuSCJP9fxjSTQQyYVdgJdkUI6nE1NrkMFim
YC+g8xRv93AAH9BLO80NYkR1EpQex7YPzim5c9Nzy8WcXzPH21JQGgVqfIOuzpnZPp/T1SuwYYUs
w1ec5qiHRaVTA028FIG0BNvkosdvLM55bXz8BN4xrfMzC2MWUNUjmJIrPeCOyQ6HuHxeRnuBUEPJ
PqFtXQy017GaTclFCjDd/RRRGsBoBYp03ax1YdFeoCKLJz+3VkuWuQB4/rlRbOpt0NDqilhXEosn
uhBbUmpMHTaeJHPjzcSRi1MTjrjeaeU7W5TlB+gApSAEIJSfP6kPEXaagSnYLTiZvXo/EiD5mA8k
rc2YrFmSF2gBPH94/5HEhH7fEU1yiupZFzw/yzq6tEL1jsX/kj+rERECHvC8H1LA1hCMAXM9Hr14
NQvllK2Z+ffjQnMSje1yIeYBoJ5Sy38ZpQEVW5bkhI6KZMEYuSzpeKypd/9BuMVU7TAqtPLIkI2c
fDAzRj7EUhQ35yddbx5RVuyI9r31fHDLaVF0kGe2exEqMuAc11tcIcH37sVWun3x1IkBtE34pfH6
j0Zqo50vAn/0/LqOCcEZmj++xodyL+kRtz+SgYDsXRaMVTo8TAkg/+mQOqjz3hjOWqvtWLb+MiTZ
72+e6w5neu/G4XfAkVA40LE/SsfAp0fQ0HefNCmx+RvgBWdv0os3BUXQKLcRJZn62UnrxLcWpXHR
x/6jAdaDUuQU2wenxSS8YK/7MHgqT0HhZCAxi7rJlsSdDky9f8Luir97kuRnGYf35RBrHjg3NIfi
Tz+wujfjxblvl0JrTDe62KU3LQE18/QT4c9nWFihFUWhL5lr/Bw+2ImwLiYrkk5Gl/lXJ3Sv4aWF
XhoeqdwkrP4QOjoFrJB0SDBxj6R849alaaRpoZiSYfN/FsxFUYpPBfbqqYH4Y0VMPClyqLy2rVM2
fO3Dnc3Y1MISPxzitfC00mBuAxprWNdvYpeLjhvLrzcLTSZfhMcUNpw1uVkG8uhpY04biCLBawWC
yL3ffeRnpK1iHiDs9D+rr2KfcTS5a9JMyVrVzVUkFad25YCqKZ1GwVcpPgq+IPe3scYkvWaijKnb
zgNlp3sO3opTltufW/0+YXgj9WpNq3zVVey+niH9JUj5boFDERYyj4tKAAQ0udNJMGBi7XgyNSH0
DfemcZ1RODjowbSSMBAjagMeIfQT2r1QTHSfbUERzZIGcRDwXh01RK8QUfpz2aFULyBG71t53RAd
9bE2qWqI4jdntv+bFJuCnTjj5ARbCQUKujnERxr3Bxlznox7Hk41re9XX0z+kNk+dCfyVLNm0YQU
lFeulkaJphcrK9mQcd90t12ekXGk9zR1ud21flCmobKtABbxQe6T9mAIL2cLeR22qU0n0IjZrzjV
GZJo/32vugIdF4C/w28iWZPayy+CmtVtpCR356HWqYmdjtgv1+h6kTOBNdUzKxQSS6gkfPXhwY5I
kltP5FvVif38Ji3PZZiO3sQaT0xPoo7Tcj3LGLiabKWDbBlaU1X9pfnFzMwm1490Axbej9qso2Cg
0c6QjjJ7g3fV6YBjPlwIwN2+fvmoyHl+CkiRaD4IpZtp/+YtqAxocraQaPgExE8OyYViqm7iUWZo
P4cL6PcVZBwUxYq/MZv9amPXkYrCJwickeLdf6fhDprTv7OjOGqjN24RqaBLJOZFzzQ/Ujkrm1DO
XEEmJmch8THPN0e9LQR7VIb762T+IbY4CU6KI8Sh3UmIg67mWh+r+oAgtLdgTB3iE8gsiH/r5M6O
9qvalkJMltdIfFq8Al9zaKuAsAtLtPKREDIO1APAFdgoisd9/vXFHty616CkvY9QlCWdx719sHY3
hOoKigMETxtmxZtv6Jg8Hqm5l/TTVMLJVVmq6/KX2HywbQcyBWMxWioT0eF1eI9dalmffoxWpWVS
aKKHskeTeHYCxNc+tYr4iOeYPKLKn5kXo3PtJHqHNvbgozl2bf79C14z0JCabuFKfU58X7Ha5EN/
fWt/16QHG4NEECDN11XjDf/l+726pbcX22jL/0g5ht7pf1aDpoMtIn5huebVc+Q2HngUZJWhQmSy
PJ2ZsTAOv7AJM19aM5hopIvX2McdoqldLTF9ajLwRpmOFewW2EUBnhklYkwpEB6q73/4F3od67lr
44xdPepgO649H2+ABPvAXzHZCkjMk7RjLxPEXouD6L/9erZKpsyIBz5AjsjKzAJrB3GgoGDJiAD9
o3+X4ex/iHZeEVgDUmUBOJZvHL/cUV306ZWwErakAySjj5KlWb36XP2EpJdTzCqE/zRRUprpSEpV
bga8K7DS/rV4UpXA8LSs5fVC+eDGRbo984ICBSl60LwV/DYW1HlA09fTFNxkePxUKoWYXbjO7J8m
pS+yD67cAzSifZACV0cIiu+QgNVFd2+CnIiiY3Z0cwHI0x+SmBxvkkKmVk3Dq3hrmbyoPZTAHC0F
0i4btWnjVJV7QqCY+QZM1MgVHzZQ32GxWRGd+nKBNB5DhlJxwzLxa+XeNGGs3+kLdWcJu1tBTTle
Nru2UpA5T2tpit48UIYrV1BBLVIZgZA5JPNDek0F6xG+Snx1kIcWZ5x5/mIN+r2Qan9uMNIaB/bT
W/jH27Y5Zu506hdU7k1tAPoQ+gaK4YNZgGvi5PwlFkTcqq6cL/uBxlEdVjUrlbdGLUXdLMZOqSqN
QmZTciWf6GDk4P+33N0uYqYu0HlHRDcbh7N1xTisq1peK7IOkGEgRUmQqkXgONp629z7sKhi7Zlw
EOcypbOfuOSfuDVADb3TlU9agunlFUAjP/zsIvTcgC8hdS385VJZLJEcKAZTasnNos1sb5u3nsJM
Q0IUPib28jaW2xD9qaUN8USL+sqFKlUOJHpcs8Udcai7+p6NfY8G6HqbqW99WO1d9Ct/Hz97MS2A
fS8Cgyq5VIDVkfOsXgbnqQ/+UQijx8HhA4Mvee9TC71xX4EqvXpCjf3mjRPhVvAHPdqNf+e6bBUG
3QoXiOsdLY0Xf+Uau0HuTE5rRjwdEYEIZ/yzmIu+C4co4ArW9NHzZCFeSoWUGgs9h0LZSEZbFtgk
RYm1IsO1ecTcpgnPxK1RQgEGeqkqPQbgTjqUK2XNDwVn2RM9+GQKXvuAuZn7nzt9/fduOgq+RdRY
JghqP3FFbt42bcY+OehRbg41C++I9xeGZzzNisU6YNM1nrgEXghOxUeY6eR3ZsrUojJ69AGhraUM
PMB6EtU3XuKxvM8mrAfJY27vm+6e/UBVAUvde1WsIHizWh/O3Z7bZDGPcmgR0+JQe/Q/fM4tClc4
hpMVMgKMeAtjozJAaPSkFucNVtrJ8nEsEJw4mt03dVY3vK/dLaXwROWbGxRBYya2Slx/DJN0iTsQ
vUh9ujdUw7k9s8chEMw7n0bY0cQlrRbaLt9dVZjJirK5BB29lcCyJFgSxZNI6GfgOvhLEBrtdScj
wuU1nFFMIOOrfGMqQ+dTM73u2Ghk5xsswzmnsLRpitYBXrQNzy0lVLMteHNF7gTQDS7/1wS+gxDF
YXTAI6QFmfT2EhNQoANJh+8wE2ZLOute6SZPRoNE+ApBfXGg9opYbGEVSBfZBlFiISs91MNaALYS
xjXK1B8t7yWrZapYaOtxFUUPeGkDMXJACV+JiKx8MGHOzCh3ChYocSNSnAZDIapjod1Yu2SHJHh/
JUZTrDjjueCn6hmROrCABIvmFRAh0oXtjUA6MElJts5BZKQkjewdNF6WPnnadp7AecLXi4/QObT+
wR+yElYNF2nnKui4KGVHvGKOYxcdzDdRufs4g8igW2/v0dBOFL7vZsh/XQHjmjGkYVpmUX01JzdA
xi2TygmEizg+gwK/ZgokaOuZbuqVSR/H8OnKnLl74284sTwrklgDzef/KJfU0pW6XSx10Sz28CEr
kxxGM09hGFQ/DZm3Jt8m/Pz+HENU2R7hGKwNbPfpsVyw/TBhDTwR/R9rdjrPMpc5skBrfXmQSgIl
JNZw7UP5arQm/6R2s1aocmSbiyzxvVwIyCWdNjhbpAygFKEIwygGmut2jOh0tiQtOurJIRxpseGE
Q2BuOZJ98ZSveEJCAmSZArbukoWRb4X6ipQm37qS/mN2Gx1NmZL9jIteT/LpyG4Q/UVUw5NSHfUZ
Kl03G1L+w0xlcXrKEq16xp/Yx6NIVlya1DKGMNsY9Ibb2phw6kwiCrxBtLrqPrDb9wUwVMYL1q1K
NEWPbSAcgHACOjiDV60on0kHYR29HDLwuSCWIZMFA5XGbDxTkdkzK2WYe47ZyWnTmvvcugCthenf
9NWFV1Anuuj4cW1CKgw8qjA/O1gbsF9QeSe+dFu52VBrXwtYcMUofCNjijjgk9Uzb2DGrXE+tQXR
OpnAyOJ5JCu4VTZLz6SuDkIETG3gGxuD6X7USG/L9cKLwVA3g1H3Dr9gRBjNsNcaFRZp3hLGSRXx
27Yg/v3YRdAbsKOFS0POZ3xQYBoVMGRczIy0kOt9BXRQBa0vI99xtEVuy5DiQXCsSseYVkpdc901
Rkry+VAokFIV2S7pQKQvUWpCN2gRK16Mo8QJmaeoktSc8FmulFny7HIHcSmsfkqPs4VTjXlB5t7t
islM0mtHWei4vAl41jnbPP7d5Aa3KO6rxy3zo8XGOh7amZybIvco/2/5ukgJlBCUKbQ6nAHQ1mVU
3CF+1mKUIUiiM74pVtcvXRj/dfULoRekTvabmIdNUwtYzmV9kbt+0odDXehHWu1ixarkVWQip3dt
RS2ef9v5nNAJqv0Aq7VGo0O1mIIagsNqPjMpf08NKzetnooJLGmoX+vi/CRTwZR2Ih2LtUr2JFV2
JRMj0PmjMI0ambYM7BN/uZ4DHGXMWDibLKg38roGP5VoA+b/3YE2m4irnzuiIKAJqVzwTzK6STHT
8D5JgaOp2AzJtq8pBzfUTR4r7zAFKQLN8L9mmAesVcQ9S7m4Uh1yJnF1mDGKKIozv4o+c6S4QKRw
3I7ZLqA9g+aAD+9gD4dy4qOgmrAjNc7JUbK9ItpDKM6JjvjA2zLgz3buIZu3QCd5cctMcFn8pi2b
T3ONv369E6DjgDkWYyshEOISLTrsKL/FgpZ4sDyqPO7TawGzvl19WfbztvKJrjrwIDBvqgVJxokr
JAdvrzfrIM0QwPxgCZkLB4WuSRnFyBvisf6CX01QT+iv657CwnNT78OHKnnX4wtk4Ek6dGK/Miu7
puYbinD1nuG9Bex3NVFcRIY8DPSkSUC9llMLX35GwigTkmzI7XlWKLB5ogpWNk6C6GnSBOPAP/3t
+sS+aL11Y/d/2B7ecqxzncrICDw+NFnKF7tC7DH3D8O/yiZU4ytecXV4lGGpGhcv4n9qwcDTBYRy
IabHsWPpKDBF6nmtIDmIPom9gL/5s3RWYX4UqYeLDJp1Ugj1PA3q+tEfWxkqATywibJSl5RhtvC0
ai82Mv5BuPwfLIL9y985dvrT+cygx8PYZwtaUVClksk563rTpxl+t8b0Bzdy+MiSLXiApeKF6i53
TQZdMyaWRAcgbTHxuCPa3J7NK+yobuL/gj0ZpVa2g0+1UUF1hqu3DH4MfC1yjOiaHcMy/BBgVpDE
onUkPZKkOLzciQYk7IktD8cP/lOItLI65qaSysKiGUzmKnHjHN+nFO0WE/Mzw6nkggtsL6O1qzDX
hB1y+cJx1fi4u30syONcME9fGVyQvPy++YkM5834yckhVgtFjP08kMsYcu94Q9/4jwXFwjqLiVVl
D5qGKoXH33mM736dIor3BTNY2s5eRLPdusO2OZEALwnBSXCIN1nDOCfIF71J9P1vGasMERw45Aky
diLodwxhfOeRIBuE5a0n4tilrTjT6KnE+Sd2Bb1gp983+lV0himm5xyzqlsjYAsV0shDHbAVGpTf
0NyypKwH0K/cQdlKViEG7pPAPWzc9ZB6xMBNLvODDC3ZXG76BZ907oug6dvOsT9fQQbIBlnGO/VA
mMR9F/ZwUQ1cFwogoOZgHtPGtmPZVfUOlTJHEijrAxkZH9dKrDnD4UWEgHYJsAjB9jyDeXvC3D9o
DF11uiZKaExsDFrx0TuQrFkEObk7bLjisTgRZ/Zo0vFAYKTuhsEKmrBnF49S2b5hMxFk42xwM40a
5040xwAhWrn2fsJhwS1BLa8S9RCHOUhoqphnpt75QAAEqnAGRo4MStrnb+ya8AM5IEAAV/zWl27C
jg9JtAU4QleyeTbvrPA125kmx2ON5iiUf/AqZs3GvPupHxUsbhjPihFu5n6kmYc1LQb8v606xUTB
5JhnL9svsT2hKZ49Gc3J/qG6KpyxJcZHpTylp4kKpHXwGg/51OvUDYcM47dVlYh8kUWZp0y+SoSN
3SrJLjeiCBEZUo7G4jYrp3nBJLoM1nwRBDCXAeEMxkOV1R/Kcmt4nOmzqXlh5eFYEtL/1OCSo4T5
xtpbJLnlK5VqUHUJ2TxAXLF+IJzVBjWBoE1Wp73t8458dwqdfq6sG7OHX0fGlwsOdexZBfZ2X/DM
3HQIdWSFDFJjqMDCznUQHB83bVZWx1xj0LKzS8vu21D7hyN/F5E4Mg8HgffeC+0JxCkKvNUETB5l
TyZm9VQETQQ0qgYajFaSVnLstCsOEyc72fQk+tMw3mur3D0RL8jzfgrECJkIIUrz3+A7duuknu0G
eCFYQVZaifMa4B7pvzd4ZEIqF6fODuAU3Ig8J4UJ4qjHYKuFGchsj2rssraZXIOkS4T8e2EN+q9i
76+RrDpAO3JFDIqmz5UcjCEb5domJ9cOPsPiA6k/UUdt5r3fFjrB3XYKRFEV6HIpcoF2nv01IY1n
WRwQsTotE/W8+znz9m6TpJ421sCGgPpg6FkeNO/iDmSm9xzLM4it+K51lNcemNNdMl6jqw6oJCuP
KvnzR3HdLLQyKMQFzy1RtCNVpuDfjjdQcLhyh3eV2A30BvXjts8P1RqUqhZuY3UIzWEsinarLVhX
Tu+NwEgKL4evo7fHuvjYm5x4cMDEmE3PeOMuxBAnL3HVf4HNGDha40mo+FEP5iIrj1O+E/Kn15b+
r7tHUfEKSW/xbd7P2rVWyNqOePNOQpHDZLaiHiL0fxdWZV8Tf2lpUgFQgzn7ilq4EopKSHllrNTc
6MWSISZ2TJpTozTzGRIPE59fUVDNmg49c8DPAlbiEToIHxC2ADbvfvJCwxwic6zBnQwFfH/rnmco
Roii7IYGArXpWwyeR6xOSaX8QwvyjLdLzzhrWGgjObvxHtNfGnhViA2hhBRusETYHTHvjOmiWssg
6qwUkuLpQRXWBcPK3eQrRs/B0yfy5NiTD4Yw1gsEXDVGIxB2kgoPwh/64G/FEMrT1ero4uvKwrJr
f6+kuCUPNl9FHnm2JL1mu1cV+5TygbV+SRelcIyK0EiTfIF7irkOtqWW78RmYOaCXAGIjnXHdKhS
iHfuh4Kriwgovqn3HEDpKdbZX1z4UuLxoSwER0S0tIxNrGa0pHBAYkpGM7VrgTpLf/IvM8FzEjRo
DccR5YQU9KbJBFiAhZsbByvm36plmz4juH0sslolEWsGjK4weoYu0nC6lcOPo2lIIXV+l7mtjzwv
5kT8eN9uc0fLuHj79LViHQFkII4E1hShgNSaIaYD+hJ1gmkbkplyQlDbArya3+AY4wfm9ul21Fl6
V5MxPa4Ig6vIKTy03m9TilhossfdAlo57718RUH2/et9C88UQEsBX96YMVcReNe2/2Pu+NF01lEr
PvvcQRWADYOybYNMw60ZoJ7Fja/jHWdmFaH88Tgs/rpSXCX6Rx6KOrjvqIec04VCirQDARwrYhZy
SMyQ5kb6VLXiLR2fc+Y7l9BwVjt4STH6TqF0JoRv7JWla4eVsyBdXN/o//3Zl596yWE5t+ykB+YG
FREeczg/dmZ6wc2++sE1Zg/n6YAVGDGnaN4rSfSAAtFosOFhSAd3c/Bvm0DP0FZI5hL7Sys4bVJF
fM8UnNLufwhJeUXgExH7Bg8Q+xe4Kk6f1rHnTHbX7w796HQcb6vAxn8OYAmDU+1OEO+81Fiut+kS
wh8oxqeoiu2u1oU7USj6a/m2Tlpcl4eCs7vH8QfY1NDY8889Nnd96eJbxh4J4C/2uvAeb+e2w2sn
vVVB1d6H3aga9YAzylK84poiR0AJcci/AcyZ+rDot9kyYcbZXupuG4VEiaaRM6JGCt129M0rChZY
BzLULQF0fEdnuPM/ukIqPhI6tUwaane493AvaV43gPx6qLI43owROxY/q95pGrV5LvWSj8+xvOjN
+RB0uiQvkpWMWIzEOWjorixPx28utKxc5FQs8tQV9z0cEvs38UHQeukbE0xqdl+rNaDQ/MDLDdI5
UUim0Qew/ezCTHtUrPPf0Lg0il2bS/qGl82/7z3SI32bJy456ED9I9p9089eAEzBW2QRcTZ7m2pA
TaMQqsyGhXA4kMSbaDa06uUZDNT055aceQB+ATB45rf/BP9/lY61vcP6IjNYs6Y4cEnJSEenp9pq
PPL65f+60KpCT3xT79e2QquNpEgNenZjeigxLfMnzQsZKh/jM46OKsHUX/rMRFApFGShL5QnWoL+
LGDU51FUKLzXDjQjXY4UBCoupWWtr8coHJaj2K5xq+dLFolzfBybyYQ81HJKKUQS5ceabsdzylxS
AdGgRYM5rgX4UFJ3z5SNdf5Vo0SeXONNUsstZ2Sdp/P81d0PsB9VLnB5HICz2PjRVyw/ZNW7kM+L
lULjbTGM8zUIQQcUxbaVLFfJwNCQYGaarz4rGU0olWUx6ppUADVpxyqiVDbCdOiSiwn75CfE38NA
OHcegq/X+T8sfTM1azp82vd0mDI5WqCx3t5Gpiew7iJlboQc42kKNaOSFaQ8WmyxYAX4IOLjaf1Y
IHFC2Js5CypUeBYsyAzvqqI1Gz7PYZos/2VNFU26IBPFgrhAKNuRcvo8+Dp7IOJdsRYe4HmGzCc0
RQl5XeZnvsNBHeJj6YAK1gGnw7HJFmmh6uwCyLKmQxRLsq4JQQe8AwShP71okCKACIyv1xuIr02m
UN98yscM5wPSVkXk/fRLeLFPBBFu1w/NhPmjm4ak5TsugmzJkESqGah/2ImnCV1faCluHIyHsNze
jwFsBhT5YF/MQPRSteYpew1oEn8DohTj44ju5cPVByQViXd4k9csZ5Kl7ZVc44RhoE2Yz9XyBnTJ
eKpAAKaBeSj36HE642xE82/NTGhSuGkvxX0Pi2Ciyyw1Y26V5bXIHTmAM/nJrtprDMllEVA/eioA
frJSquChaypGRquYz7dx6oM/pycAScGZFbuDr56G1Wr6YXClm0pvp2BbxGK2MZqnxhSzN+8uWHv8
9/LnsV29Y/OIvw3Z8mokx3oVyZKis/lDNcsyULySj/kqrDcypy07NHfdgrc+DWDXWSXhQd9EVGMZ
h1y+RGuTWwZW85+U9E+ijP7sNAVxYuzAHB6g5JMruipR460m8TgLC8+DD5CpAXEs6hZMF8tJhH4l
YQY7XRizeq6Qr0vtXNTiCLt4m0VoVdf3rcICzaZjMIZZqQjtSnD0y00ZdwU23Gyhoiq41ztqj+py
TbfpKs40i6VqHPmq5oOqk0MSj8TuIAaREKYfMIj/vOMiTrs4YaNdCUsz301EPI1/rCvn48dyZZln
1HMIkcc7F+xzlKg6WsZyga/7Qx08o7rnME/GTDszNK+6i8jLkefPNQogHeWHedIk2zpdcomH0PTJ
yOwRtirdRVomRYC4wvOs/YKM9NcxSWFtlHSO04A8FQ7jWmBbkbdX3P1PzwZ1J+Dfv8DqYEn3jeUJ
kEU+14licjnWqEMaeEcNW+kM+ocafRy+Sc63wv1FdoUsyiy6FU5z3uAki854wAWm0eCnxJdQJSon
+TP/sM8v2EaBgXUziDYW803qzTBZ6Z/IpqXdVZoP7PCPa8VaQDu1R11URFIHqiI+swKg3djeGVfg
22HQAG1EVSItEt9tjjaMOLQL7AwQg2Em8ddlIKDrHGUQ+/v9EUt2oa8RKryIWmXOPtMiOLSnCXfj
E0t27ePm1we3qaApNUw3ID8kP0i+DIbPF1I6OYjWtUN7F1sF2P28kC/lBzSAROyyaxIkj44N/wqW
OG3/s62yUfAPTzRT6YYIoTSlMQZ4T3FBno0Fr5wNabcCj7eKPkx4r6aEzt01Yo6W9ESFi7hgc+du
6+jhgH+DBqVTDKLuisiRizhbYyK7uiPt6ckyeUts7s4Tf9Txsw5tYB5GLS5THJsDg2NerZnr/8Ol
RUJjtTysIuA/ZMSi9oe7f3zylFGjD/RrCtgELEUBXbnno4NpjhKGdshRkWUtyQzndDyi98SVGXL7
Zsvd7TEKaH1uRLoZGYCMC/i0S3lGOErh/7iQd4GgMSXsWW7LJp0wCGWg5Fjm4nBqQSjzoAGXn07n
Yi+A4U5G3Gcqc+OEI/ci6KP1eDYnjAL9/FeTrhrZROCKyK8w9kESKu/8dtXdJN4wYnfMXZdK7bJm
sGlGWbbGmhQ3sLrK1lR2wlERuo6ehjD8rhiJ+kiy2b7mjOvrJPFuNNgu8+0qHOEhLmdoeDRo4c1t
onEDxdOdJ3cVbE2mEFm7wJ3+uBDuKA7DqTE7vcT8AVnytt+fkDJM94GN5M3slicaA2AHO1h0uJhU
mG7KgPHrA+bpjTpntKzlKXpklAyslPS34pJtsoM4NQ0jp7abqM3vc3T7+IKZxwQMHSQrJv/2Z6E5
GS1XDh99BeMEAeHY9OLiLK9xJPLHsFUYtF3lgnPYyyzNOTDLKiDO/6PVALcMeHXR5P5cYG0ePsO6
fTcdNzBroZ2/I8qrtHsqNu9tVE2S6WpfVjx4DHNbDClOz/fvOXvjUx8IzhpAdN8gSDnE06QFMyzd
STkTTkwUqvaiLINv8T9ziE78+wu2SpwQ1vFaC2/cjew7r+HovNDeTUqVGNyef1jPZiX5Kty5uSt/
c6R8xkJvOAf+R3XMBCgivwATAzcZWAYdt0NFJZbwwEsnBT+f2nSSUsRyDDI1VNdVTbtDVYDP/zN/
zBc+i9QVw0VNSiDw54RNABxisCaTCNGar5JjcYNnyCsrWlvXyApeani7mvc0VjrqHurUNeUEcBza
CmVaDS6OLKm6dc1CnmMJ+yA/QjB/xQ2LU22sOuOpEGHzD7jM0C2Pq2RRPYZt42oWIgEtKqd5c+sI
z2Xg4oZJYBJ1QDiCQOnjhmaIejq+M5Aq8QORMX+JD3sQYaQb6B+bm15B/02ZqVUwyEzCvxHhcuQU
ndBZO/jXRqh5+/fs3K75b+U+GMhm8OGzxkFtJfimERDX/TI8AgR4Hti1WedECk3D6fTbWJSgKxxJ
/Rpd6FwmIwvKq/nNGOg2vFKtoN2+MhtlsxtWTPEEW1jv0gdKxQi9RUHtQmTn+7oDsPsuyJ/LAzE6
pdk6VP9v1BrKel2kTX1hTxIL7RINIPExD9ejDfie2laoIL/Dd1m7s+Q7BTZBWy97Okxv+2pkgrzY
iPI3RrxcjBXw+jt/BdM4FI9UYifWwzePWrq/mZOgburd4IWnTj9POclFiohnN98UOwA2Gy73alT1
/NW0hVF6vz+B/QZwNgb2d7sEVvIkzRk/BvYaKtMmZRix/CvuaKt31cwSs3hwZePvsQtRWpotJatC
UjOsHkbMcwVc4cqaSWaCbnTF9AlimfZrkaxf5q4k6mqQIv68WiU5jMOJeSTYPmoef8HNhS0kUBSy
ZEiYiE/5nyWMZMzS9+y5uTE7YgBDH7Htn7BhsGtHwGctP8NdSdk/r6HfbZ5JUIEcZ8/8FE1vMswQ
HVzuC3oLHckJLKQ3lKo7m+hCQSl4s3QHXsRXrpaD5N36t5BctZpGladeQKxKYKSQeVB+rKWK2x63
cC2bw64RpeXTStABKIvHPNaVbXtBidctBGw4fvyhD55zyJHpEG4A+shkVHoHo3D1r5Av2mvx7wb3
1asL6xb9FddrfPCIYGhspwycQyH4FAR3uBoMJuYh/o44jpsm6ecOpi4MUUwGp6YUCOBK80gaMELv
yIXiB+yIm/3xAkeukOV8f+C8YnnuU/3JqQT1yorkoipuXm/rKSCLFxpSaD85vxUztEMobwHL9/FH
9moB4xlqoim8UIziD36TKgYtM+YRqxiOnhSw5H4qC953mA0q4vxqyflE91dlhbeQUJmIrDuPRFPO
682yzcWJIzzMLZ0TeM6UpESpQKwMPveYMw0Vl5+TmF5pOkuNe7dem3Fv67s58iM32dJs5Bra4bet
qAFOPz6pk47KPLmEK4pJHoQ4tU+Rr+vg7WPY1sPJG56p2GZehZjovr7C4s2F9/RJCQ3fQTPUjE+A
vmFRu5coSKU+aOWr0nfzWJmtvsLHvHNqhWNpGhtt1U6glEESSXtlUnmhb+atl+7Pp+A86Yo/fP5K
KuoGg6ju+NV9vZvOHkdZ0TsCjsDWLvq5JvX0LWz6AlBRmPgXeEwdQrAXA9FmWWrHbgFOis8nlOhD
34vFwrB8+uYNDWstzxyZv5XztsB0Vs8FNqJAuMyoaXq+14YlQwFemmOxQ8VkMoJveoYRhU6BVZuP
2sEpURgLfF49iCn+ZX3TF789Z9YgIo7D2bE8lQiiWkA24QzKM8VOTY/0W1+wxxYn5E5plRJu6rg1
e41iExwXHIR/o5e6GLyweJUwYEqNLAp5mnafOXtKuygRbdJ5i+CdV4EQ9oSY+DOrNzWIRdSe/EJ9
EXfTC+QuEsbtlTtL4oLWzVQHNStrrVpFyORDmaZBy8oCAhe7mZPshSD4pFc7Dya9RyP84QVWweSD
5HQhCix1jIoYr6/FvHfOwxcLfgitLAyw0Lj6edergq1u7i8TlNxrawUYCkx8+P5EkaXxppTawLDv
rmhwg6Z50QdEP8VzV+AtBdBLK+x7QA0t06jbF3IFGJi2kWy10ORdJJCzYQmRGTw+bHI27PpDIqFk
biXOWM1fd9zh1aQcs/Yuq28vZGyd4lU6DyvnUy1saiLfk3VJS/CWLnPbCYBGEznjAk5/Q7VjkGtx
ksuyB63yZtIp4yYpV30Mt2PuuU9dsMbdX2Sy/XqBKfuP0fOutUBRW5nXdhQmQDYMufrO+yOFaACx
TdIO9lFQeXGbUdXFyDZanBEooSULF22zvRs6UWLYnpGDG2eUpLUG8Wj/c5D1FfM0Oy/isEfkRLXB
09DUrW6d0pyrLkn0d4EJoNgEir5eeaWACyC317FpgjzNgGMZaVryZEolDosktGfYCTKBBkRad6TO
37QdAq04hU4I9mDS5nx0lKEM5lS1eRUoOhkTvn7dGwI0QgD4FGO8DachI53q9lNEvLOUo6LulKUv
D/fhEKjAdZf88AOC4GjdhBnI6K90JHWclj7fVvL9vlsTIJ9FHrphYhJxWIt+sYU/q3/kN50NO2R7
BgojtYeJP34Zb+IhFnY8Dsak2kWZq5qU3k+qa7Ad8bBVP4vFi1CV9uoZsWoyNBZys9WNvRy7pbIv
tqTjizhIb5W5HvIvPmkavjzmfkzuCW8Rqm+R/yAzFUH3GU63YLNyWn/DucD6Sa/7jynp38VU1JWd
boP1pdA7TN0FD9is2CheCJvP+8oUbgcHJn4MlVMio7Nngx0ZFtOIqrguxRpxsqq7UDTvS/U/vuIK
NnFNU7SE/rhObWDErRKcRkN8CisBZNKG54I881yLZR4VFbuuI2N0up1S0PumWkIzmTNVe0Kx/nzA
ucjZGrYUzC24ii/ihtR0EDH2A4CHGRL/Z2yktM8HeU5yjRCauuHDDNWo1WNlsTIzuL+izc++9DvR
AleBL0fgHA6/9NO1YswUkjLWatcg9z0Pgy8+ya3StbQmV2Cgr1OxVXISCI9c6RAR+1aI7PDVBg69
uBqhuJJg0GfLVQHV+AGfr+O8Okj4h7MJBAFvaK1tMaE5L9aPETqvzcLiA+ie0Iu/PYiD/rRhtFVU
sdDh8Cd1/6Bl/CSuOfEeS6n6i264v4SRMdK+79VC0UNEGY4fTdRuVsj1A7Po4ew/qZL4BBfPcI7Y
SXRsryu9O7zpSQxtVQSi4h3pXU/+l3VsQrKHij9dkYbHC6cPSAe8dix6MxlFcyLvOI9nrRk7b0KT
NHt7tn38pAuWpfgMAl8IaKTT0IMQPbTrqGqE4ZAZS0rqvpA2Y0/ylXFXX2GbEnh+A3Wq+HfR4Szw
DHPv1lvrrXnR6QCIJufeDdRxrB8saEj92w2gapyeIUZfQZF/0yDi3LIZlDB+2KwrnRNQSFLrtOLh
Dct9VR/BH7bC3PGuHmXVz/AbByrZhrLhoUJyA/w50dElWUi2ubf4V/ZcAWKAwo8M/arXFVvriNUq
LxkGGxOzoWqb53oWEnXao2atrG7RoXz0d0cymVjziTX1tNtnaKuM/yusqElIH0WJyenQcLLu7iJJ
HMZndbD4XCZpVzQ/55xBbyCVW9d9lmdfDhPrHd1qmEfAaq8e2/9buz6YbYGQC+UFe6eDOCRAHmn/
4PRztuTkkCDnOr4PO/YN5oIDbUIbXGcq7D5/4VKaNE9iJQpGnylDwOibelZgyr7vdbxVS/s1IGwz
vjZyvs1qJbMzG4i1tOSLjnzas4RORP7VeYy0ampOUsbl+dOwlnyETu9tRd+wkT6hW6D5x5OCBCsQ
g92Dyv4fM2EK2n0wX5GiZYqK4iQWj4wo0iepcrJl0WVyNO+pLMFZ0x/uBddS8M2+LDtikvDGoHa5
1PEh1XTMIo8GrviNT6RC6pkrBkv6Uaf2eSZjhSPTwR9H/A5kkzVR/E90gsEWPpbfPHEu7AJ5Fq88
GbA/N/ZJNCqaZg+zVKgBRkrHaXb9TRppIoXtnk2QvGBNHm7y8LXT/fTlp3p6YpUO9d8di1FgHR87
p0e6+NIGCkCumZEWTRu6WA3i2VJmnQErSsCCnIzuy8GBe2ZV+XVHaMRvHWPBGV9XkeP1WHsw8Wwk
RceojWUogqwE5xaCl3acg591iMZOfWFA+pAmgPUsBd7lipu3kGsV4YL7W8Me0BO2o2Lk03PMX+6h
/1ucXUEaNwcoGepjonto/Q1/uaBOfZDA77EoIymgLA6Z9ev/v384MpugTgK1qVo4t1+EafH0A9G6
966X96wZ6ZtCo2pSjWXn/JMdQA0jSLqh5s49FpSd/R1i7W8BR0XxfVcmXEPJ/JZ0tPmp7e0hhzAh
gz90QBWNsVhJ1PSn3ggLgyLCTKL2DsQnIYYB12op91oiaEdVSvYKNnIXPPon6bxzISiuPFggUD0z
PTAstxUCT7nVqiM6zMMus9EaPrnJeLr/vmVgsCP8A4zdFysvgmtURka7uwkYNI7cRvPNJ3Ew5bGt
DnXWpIf3ExDgze5/Nky5jHFhkQvRMz4Ul73PY+kFDuMHduwLNrugNtFC6jG4zamyKgtkO4XZNbF+
ZWbb1UZ/Tv+G8aQwga27Unfz0ftUkz3DTgCPNvciv+Cif8a2Lrw22l2YpJZNUsGjcKkpZLy33x1K
T8Ki3KntrLIKk8KfJzsaiYbKtDGVibSu/4N0tDfFNRsoqEAe8kGf9orYbnX2chBS0D1KT37TDBAS
Aaoj0nwaC2Pa5NfetBM4vgHo2UM2EoA9gIFwkFxii2eoiGsCE0ISJrGIQMg8sauijjuZEHbcsT43
nwA21AywbqasO+GE+LgmUs6QTAlQ/FP7kBkgpMbPoTDg86b1a3phn9kHx/ricPhpVrcMzfKxSzAM
+9gqO6yOOo8JZkdvEfAEtarYq2yABS3WlAMCs62WWQ8BtVxA2JUQE17Y7WXjStCh1JNcw2QFaxQi
ik+xSfV6d1HmYmQz3ckFBjrIY2nAy8C+8wGjchL6SOs0ujLSAVwJefUV4bZBVKlmwCWJYR3wIax+
ipNy7EfLvs2Qnl6XLWjkLOHSlIRU3A63v0uQtAU/0Qutn6Gk0jgXCYwbIqLta6BWarhQrFHC0Vw5
1XDNQHFNLX1ZNBR359V0UScO7PgMfPaJXJkoToQmaGIv//i43kElBpc9Fr0Bnq+CtcT9mYphcC6S
9jLOrJbJicmSgjKta2IOqL3uqXEUflY5oxeBmkgmHNNjJvEb+Xkn0U+FodFQz9pqK/7WJLl2njfW
AJ5kSQ3/4261p7q2q6mNDdq35Z7OM5NETabuXkE/ZPWqya7pjoTnhgxsOLlAvfNvklElqjXX/FKS
SWTSrje0BhqPxM0FzWfMK7ryopAjIiaRPSVMBLxLePI+VmkD6NRB/CsT2G9c9lsI2C8omRKWsrTE
IvZsvX96H7BEWYKi6hFzHEALPBesfEnkdMtHkVkzJDrbpyQTAANIwvEw/KoeC25yOZ6n0PY85tZa
Sl7oprGHAPFIsfJSTsmG4vptRHQuVY72/qRAC867Vc4N+GcMSuO/QNGbxwgW540r/nTRdhx0OFY3
hgh3QUPk1wTGRKZrJukK6E/afalYfkMHpCHSUbQboNUk3ml0p5cTKj1aEDOFqWbpIl1TTLVkuYQN
o0lJ/KCLZjlptL74XiS7m2i7arMyfTgg9l+Kz8m2LLTVJ990TvbUlhZVNYVeLDFyLMPcTQkRSYol
KH7JiaeM8JqK98wz7ObmLQyfcnZh44AEDSsMIlDokixepUQXsgOUD7fBRnQCQMlngGC9mTuhI8gi
wucycpCtxl2Zu5KQamvrOjwOqE1/qQIobpQiM9t16x4kmwxoMYDiwjsrEPcAAbsTb6X6v7SFHQ0/
CnBI+S6oRCOVmKCuVknTmT17jtobPg5w734oTV8I39AQ2iG8CqbUjfEGTU6yixm3zonv8yJB+lNC
s7we59SV+pSjiJDPNYajIPLoHNEzb1T3JNGD6kvMiaCb7SmJ+H8lqm5f8vfaO32YD4JYCAg6v/l1
pmFf4LUWeYQt1JqY3nWvwGwFzIE0xTJoWKA0V9obhrPbU7SksD56M7tYW421rrIDLaipP+alAV9r
PaoENIb0SG4J0TuOqQ6R1Zq7LWqRmJ34eyO+eIR5YCa2iDw69Vpa0fRexxaES4OZvMzNoDogZgEZ
binkHLrHwH4hO89/w4PMKyFE3Vw5dX9FU0rjDtl4NSjy6xF8R4RGslsyWtjOMxG2NOi59wfTTjda
tVRyaCrG8dlN0BjPOhTvIlqapxgLhoZ3O9xgLfCCfVdu+hAJtVRi5yOyHXNdGcDr9KbctfVePbf/
VC4J3SHzlGkNbd3bF3Ph81ZeA4k0kHOFsAr6BbobgzyyUjMxfK50PFtS1jUxGUD48nmX5CZifOTp
8YfZJfsbHgZMj1yYJW5LaKSv35SKUXDacpVon7zDc67FnPUvxdev5zz5nWivdt6pfUutmEHrPRe/
WsC4dQQiVHggGQ+sO7Vz4kkCDOsnHbqbBLcsT7h26a0/JgK3oFvzfQueWW2gTSqk71Qdha3joE2c
mmYvQ53EDU/SDYmkpy0fpzzT0Bwt/WyVI7jXbP+nHkQvbB7y2ly6trvzohg+GdBJ/1Jot8Z5WN4T
44AdQ9Q34hBvkHps1+U2MTLau9W5TJ533iP813YvkxluXdKZCZ8aEgzl3k9qe6s0Y2OoiYvHWZTm
jc9UipS46uNHv+7rgeq00pQUWw5MysmDQHnyyHa4I4LN9hdjtMZJVVEXFwZN90lGO5nQHNfvxvZm
9ODkE71/oYaiYXWOtflTYW8lbVG1SepiPZ8H9u1omo3KLghpoDMkrLXw90SY0r858fGtvd5mBI7g
2cqhlH0IBFceSijK5E5NIPxeE/W6OTdBo/rod07+jPDzcPxHNy4QczA41f2bxFkdf9momxZNTm1Q
EUnm2qdcQrTyxmaqfSx4QqJV4hXavBfnAdGmtD0AXlP5TwQisxOhmh8sQ1gDk9Qy6FaLMt/iFM5v
4wXDfecq51HZePdZ5OCeix057Aoy97pHjbge9ffmrAVxlrbHZQ3/fqUiYegHxYnoCFZ4IS4ygnWP
hJQK1EvmZTzdRmBXbeaqlIg+Lv+QuyKubj0dij/dCEOPkYeODxkycOh5pY+w9PjAeSv8I6qKcYPZ
1g3oChN/5/oKyimdAvy6ddKHmaHKCwX2qzBk+0EPeWgYvb7+0HZhYUtZDE21DS7+5F7MnLPNxaeS
6LnVUa8GXATFCOU4bjEHf78dyrM5X5XvK+oo0msXI3XJXB29FD37ISKDSEix+Clmd4eQY8lfb1/j
jGY98Vghuy2ehaxiLL1CAplxlZazJxXqqT2XOcsHsOLrLTD9k0viJVDdLJvun9/i4eIVDYelN9Kq
0onWvllBtQJ1/bg55VMHrsYToYUg19HlEUpku8WkoHrtQDe5mhS81qh6aVOSBhbTw1TRpase7rYa
XBAh9ydMySxQ29TL+oAgFNLsiF1IUm9abbqa0N8lp48iEHfAYJlX4ckxgDcjEur0dr6hJ4kaGlcm
ZUySvMJDpMtZTFIVOuqoSAB82Bg3JVVwboXnhjMiWj7QmD0GVXi0J0JLPIICBjN3rV+oWOAXCeK5
HygXOoYa0LqPLeZQeEe0DWyEENaYn76nYesNKQjZnX++A4YJ7gZRk4PcPA7Ej0DPgc8DoawXGsKz
DrHnkD14WQ9Hz1oy5aCCoUxpxgfCMqCPrXoXEjD1OQdmZJpQr/ID0ylcvMYpt17h3t5et8ondFCy
+0AGhJa2mlyIP1JZxDtVIuTMcz63AI/44oZZ+Xkphtt+zrs4/acbq7FNWRDAAUNOmrDmXmsM3nIo
mKQkurDbur5kyfMTAUpeO1MbQU2xCV2AMlINwEsK1U7td6rnlw7TF6gjw+4FfTHtI9lYr1oDhbht
7auY/dDULijvDMN8eM6kAehSfJmM0X8qUA9rGS8xOOgJjqaBTLhfiuYg59P9ZGPsLob5K1oIEmq5
7BvyQ7zxp78oi9d7i2WHnRz58Mjbh9sYY+qMrvx3d7++wHxudl/epe0Lgo9LK9Qp08xYem4oqbv1
+CeLYI3XfgJEDxTmEoDiksW/li4+ESfnv4oj8+VUCQWNUAfWTeYzocvbimacYH2w5l5ByrmUId6O
pvCtaBPOM4CAUeB/X6nTU4/By/9yx7cmSse9t1toMQ6DVYLVJYWVpq7udEdncHrj0z24WbnYTirr
fY/bL4ftPob/ZVYbLIkXH/LAvqu5ttM9SKIcrBTknJfncFD7CFYhSlXsWKpLwkRT5nyfwUjEhMro
VcvtmjLOo8Z2hasRAANULCf3RqUEfji7zH2ellBhLphTl8kS+MnYJfoL2FlYSPGyZntrYNyny1sl
9G6FlJZHsAgVU6RLOeU6TZvTpbGB42X4bow/YQuZSZt1YXgGlTv9ZyvNXr9IL2CkW3AfUerDjXi4
JAv1aptoFxvGoMN5cpNm1ahXgjEm78WZgQhamLe0Y53M+j55pJcPlvABVM+RXNg1R0YhjzQLfv6t
rE8mN+eYTPv2FyPIidVHV6D0hmURas//OSn7K0QwSs8nwwMPayujUoPZetu2+c4nZATlBPKgNYXa
MmdidC3/JwGLe226Rk/zSEAonqLEq5obYZeT/EuR5Ykz/PO3DPBMXM5VygMa10M4ozSX0R2vr7Z6
SkWjUm6A4z/9v4Exg/uCvp308tHX554irlBslHceqNvcv5nju1bjXdvC6uZsp4jbZOS2R3ev5uRX
E9Q0ugksMimW067/rIE7ugS1W5HHIDpq2cnJqsXhHkzqYWofokQ3AOJ1PpDZma5IIiSktNsocsyR
3ZSOpxaKcQbM7moMY0y+2NqHV8KYI7VmE98MG65AHhA1ke0xrIehMccZgtcYsD/X8RwYf+ld1nbf
0GrDxOMoE/C1brb7WLPTs40cCH9UXvqUBz9B+k/U8XGFalhhnbSGb/3eWO63vZXoHpR3PR0Lciom
CTMi+fCjJkJFTrOtDvLQf4vb1O+ECsOQUX0xadxe07IHjKwNUSvAClABdg6iAckBfi5A6EHR9VLt
IC4w7x3DRfZ+CAmVR4luDPLvYd0DVhTG7e/ptp6LwUvw/dS7m3a7hOxEJ5/LJglcI72enGkz8oJG
jsoJuVx4tuXPrCm2xXj5gaambD7eZBB9jcw2MuamcaCSPGq8XWCqEZa38RngD9UM/Sl/0zMp8wZK
WRIuo93q1iqRCc8OEbSE1ShmBD+XUj00ORpWpXJDh3NzNcRnRTZkxVcVYcdR77N9nkGx6qxpJRx8
CmJJ7HJWMytmb/5t4m6F8J6jMALjOkWs3Uych68JBClnkz+V7tHc9qGhMTiYgU3JqIJ8WFmr5eBe
KAn4t86PXifSC3ewk8Kdn4fNZVa69q7llMRmE0EPFfDfVLk0zjnRhZDeVJxcawoDC708IGCaelT2
TTpciGd0+cUG6oBjKgHYb5HHnh5Yz5Mad7KtcA7UncUZCHGLixMbbqoE/erRAaOhaKKcM8jIriBR
i1hPH1duLK0uZip3TZygUOKu4TSeSK36gZtgtlbMoGy65YLlDwUFvQ9mH3R9OByx9vNUFV6dzzqf
ax2kLNcLYH21jWFk/tJtlVojU/L+Axujpoy1qP+mM8n1AGBVFVm4d/kU0XbOkbPYaByXXZMKH4Km
RzjsPDYsAWq0yuAZ2WumQbmTdWSwcGnYhd4IKPs9zI/s9/o+qLs7FuyZ540Jqg7OgYHHL3kYdwUY
0N4WSPAjcYOZy1z0yGF59yCVVdZEX7tS5Bm7+aVm/frolMF7jb9cFsDZ+5Gdn4Z+y2yKGPh8NAxX
BYlrF+qeoSBwjx5v6lRnidQR4vVyPXAVqX7P4TqAT2mBurr/WzSCkctPQovviiApGvbKQp3xTCv+
Y8JNtDWhzSsybXd3MvbHPM6FWo7hsiCv2T+iBWlEGx89a2EHcUoobBtjzKGN0iKeVNNJ26MDxd+I
o8SWsIn4UWFKVzohnACv7lx5dTmRDapHHZKALdXsuAEl3L2azsDj9w0aUfw3RtzZ6CKAjl0ITJWE
5P4QKm+BBt/ZOloqS7ihqpHOrdJ7RRfaVs+ezEkhx58exZ0uUQ7kR8vQ2bcUbVlyAhKaYCWnL6Np
YlZtlnMn/wfPAeYdcmxrnFhqiCZrGgeAH9Nb2haXC4axlJXfVtJhlhQre0P++JnRm6MLX669lWIt
jaVqirOuH9F4bJnyWdGJuEiOyG07FvO0xWVmTyYLnGnZhiqeuHxCGlW6q4vcH0Y4qIF6EK+XjzwQ
3GTU9q4Nn2+6i6Bu3MJtfv4Ncm2SMCdOURS+iR98F5c3eXzLUk7mDDOLfbA4iNnjBOdY6z6LzxP7
DehS4dJVL5qMF74cykQhNyLYe7i5wICWPqRbhX2Rxl+Ng6DOvFjVu5/9Lm1HywuY6a/fjRX7rFVz
BuUtk9hY5qS5TQ52mlHQzDGEtmqWJflOu76R24uI9T6u6Qut/l62a7EhmAv31Sctg5fkp+cD0fwl
K9fN96usXfBfUR9oR1X19kWVaPvRXudr/746+q9+WjuFGAtkBPUPhxOT+9bmzquUj3dOdSBd+f7x
uE3/5L/HMwhxLuLgazp50F+98MRE/xNK5V5gn753VJh1CvYf3XgXDLPWtUllAvAIvbKSxdLF0PlN
2nE3cNOe5KKpdqwRDisWy3zRT2Ho3wuyZi2QLWIzK+BQ6a5QDXtjCtTepoRALZaphjhyBt8jJiJ6
ycVwcqS+Pr1DqZc4fshQgmzm0w1HhLIxm5LZZZTsel7Do45lF6GRYcCxmrBi2ZmeoDeky6zmxGpn
n7b9GNz+dQlms1dMBiKZsMumQfRo6wYdi8ixWDWNTQD51XGu7Q76EdInB9DhjZDTBpSRE3K3eDya
qTKVMdqg04ddnfx0Ds53qJGLhHL0p89e8N5aZozYXlKr5jvOTrvTMfuPPULLIdMShEa7h8OhXwIX
UhEyZXE1EmqLw9PgyjFXqYkrKBi6OtERUO8K7UeHGxKF/GUFyzMdLvkQbQNXxaza9e+rRcRePf7o
jYuYaZHoM6C/1c2qWOQ3fLkfQq5p8GZunlFJiKXBylB7l6pBW/MEJupvvaFaznAQMMGTxl/nO0U5
+MiyfPvPlGoOSW7XeKM/pZEyhK1me65MYtS/5CISTgLNaX2yD+b5TTc5A3+si2Q0FAPMXP2YdO4J
y8d/OrWamGsZyP7NS2xxAKJyHm6cOJ2F4yfBwn5BHoB7qFrqcc3TdC13uRfmbFwL8JqNZbqM0rny
sudd/UXXYSruL8eb8obq1y6Cp7cVkWcqBkdoLqav9rqZWAMIrFPcHId3b6jEN1rm5WzVNLdjR6M9
Q+SSN5cSdlOTIuHJGEEwzuijtpy6325p8Ks0x5Mjq9e0GkMTGDsMg/IIQtKEr6Vyq21iQrlyZTSS
W1nVcqons8eid9IGe73Ov9QYxACMxA0q44Ev41L0Dq53gcAxrra/wRYnBABH8JB4pD6k16ttUgW9
xJhXNFuIlIa5FUyATTMHFzvjj8N164bZNuhxRT/u+y4/KgWcBuYflDo+uamd0fvTVc7lnmyi3wI6
jXLNpOdameI5cA71VrPwNeQQp1zOrv8TtmcRaGYLQhYwvW4WFhj9yew33d+Du/fjJcZcHGvWKskq
ah9lQya5eWtZNom9IIDorqbamCvcngKghNENtptlAuOqqAhFczOegIS04a7SzDyFSVfNWnP6xTyk
TydvDntdFMo6qS4w8aG4MItOJypr0wR698r6vI85IaMOVoAsL8h4deDM0FXz3uw3X21KHnSUeyou
cEfL6P42LtKR/aUhjx8N6DEr0VNYT+b34deAVs3prf1Nt/S5tgL7i/l1opZdmaEMYakZYyMdtRro
eCVeF6ARFNSwDimK+1UlNNKvt0rnbQb48qXeRWtSb7GQ9rNn9eiERtw1aLpW9IdV6E0mg89sg8Hr
RD7XNaQka/DzXQ9rlBRgcrzG88cvRTePyc2vyQwq0Cpm3/nqgaxmI2i4gdbmbkzeC90uVwfGNcvs
+OgxjyD7VNyBk1Wx8qmPRdrvNqBUtf61nupR9bN+Sdf1ahm2JctFBS8rMMT+fJFn9WutiIcxbP2o
bynGKV4SMwCqPge+Coy4JrJkamIlUVRX7oqeApAjSrjT6H4L2+hCKb8NUaGqcvJM/tYGVJLMZ9MU
YCJI7IoLd1eSx9bnwSKlK7ohn6Jbh2PPXyE7tzChRjsNoVjS5w2p2ESWsQOQfsTZHFhKIR0c9x6q
JH32kMLmLGsv+yN3MI8h0XsE++oSZmu4MUh5nKzFPvBvty/92zmOBRVloGwJVLaNxnakf5olynF1
JK5eTeVf1lCNmdfPhH2r8bwV3oSdHqG2J2aSkrhty9TSe47dMpuNmUNgqTRwivJ85Dzk6/0BZ5/W
RpVACBcc5jijD77hFiXGMw5lNk+MeS/zUuvl1waUjGYU5PuLcdTmEh1xZpRojv0Eqoxg2fgLgd05
rCy0/fC51xY3rd6et2WZYMpuEETCJ1GlGOYkOhS1dGfU6XQdVKMjHuuOabzGNUQTvOD+PUw4Q4sV
URTdgmIhm45VKLOkorv51kabvk5S5vNwD1MkQyZ1fDcN/8SqkqhcU5IiElEQSWqDfaCpmrhm4k0e
LBkJM8G4ZvE9OuDr2SFrHkflQjx6iLUffCRjFoY8UXB2stmRchfzMrRXEQlgNNJVWcpX8EZrOtY4
2bonRdI0puxWz2akhzBX5PEA++kCd5z0iSYGjbxnPlCowaw/DKt0KOJV49nfDrn/uYe2cKJ4lrKj
1m94Fs/cUqx3yy92r6FMW+vDoHsFk7IkrZWaVP8K8XPijvAEd55PR5zenXwtA5YaIGYO7c0lCCOf
5NtqQKLcdHFfjGNl1AO3jILJxDgmoaHXpqeaS/pruUwJU38RTWc7RmCvwGFGx3x8wLHPHCp4ldS1
nZvzc82FAMnl20zheNGu31QtBBzbiEl2FdMdxLunJlORW33nsPUvmYkh47GjXvds5Nm+Ctc7Ue/U
MJftqElUSd1VG+kSmh/kOgjo4AJiXeMg98A5P318zXPB7A1t/Xw1LkS/83VhK3cK99tF6spzsHYg
bSkMiYAb76vDVolCWlC0wi6akrAFlrgJoOlE3B3iNLqN2Vel1llWUWcYu8C6wql3hqBzOQY/aNLJ
zwRVGzZs8QwAvd4vBHQHZI4Wa+WTXvmPgULgiz0+k78hFvQcB77zz+fgRv6eA6PVy8bllBa/cpd+
O+gXmHnNEEE7fMPkSLPkZosNJf8Udbn9JLR5NrVw0dbE9I7YoXQcyPcPE/PrME6mXfiB3wtQsVHy
Okc6jZl7eD6YHt9akl2BkWbxhfFTJGno4tFgpLSe/L7bY09nc0/RQu1EZPEFoCoBU8wlqVLcT4Ef
twAd1IAVyaSvGqQ0/Uo+tQC108VuFXJNlPvKKmuQ0JO2Fj0lE3Ac2h1F2Gc5zDgXKUODThb0vxxo
2pU5gchVuV9EAYdyz7P/QxHtwNQSieEF33CpnPW/NdP2PrRjDAxsMxn2OAHJRQs2ERL8OW44t5NG
EQO1NHpr/Py6//3w0bFw8VXQ2pY+I7WQAVNrDz61K19yD3dzJ7+Oed6TffbjdX9rVpOWxZXwxxhp
i1xYG7GkRXw7ELAVuVyzEqKLYkWt2ZfMKdMW8OLbQdYCIC2Zhud1XjMXLkOUpC/yVhrdMF1pOfdV
cGt1jW2zh1eS4zqW0d17HqbetZgQvMsHwHtLzB62iEO0rUj19LltJCzpQX+eoetpbuuEsYZuCW0A
XjKaAyLq/XFk8DKHlbGAqr2DS+jjDGwCmKx/n+wIoBNRSicM7eJhT0WulLvkeuMWtjAv1lZ4XcJK
1aA7CWvMecpLnOoUjMLFsQGdmi3r/reUHpFOA3mVGnMQL9O2NNpLaTECwZOyqBl4NSX1dn3IaimB
901iC8MSw3fzBWubhY6LQEnP0HhE6Z5JsgIJOzHNz/ysblufrOdjchRdSdaE/Gbz/qFGbs2HN2Rq
pEdDJn7cTXJ4aN2tIX/668P/wLwv292PM2NjAYikqBOEvB9DHxEb2iFfJMCQ6Kd7Ta6YhHJbnSLe
CRIUGzsGl22TWVOz7i830Qs+wf4RqJnKznwYmO+1DDBLM+7nO+Q6G07aeWXT8IXE5WRbfsY2NwRf
CWBpL8qJyL6z+YnZyTDb2ULz2uvMkjH1ZS0OHXswLTcx62getOFihqGUpKBbUPOq5WAe6wsZ/wY3
MnXuZdm8K24tJsW+Ey/LJeiq+RLxU8HBtYI37Cb5I7X2Q9zCgD0kd0lRpU35I19T9EZAHhvZxjDZ
3WqPFNEHvdvfM5SQUJ1LnhSFYginXF5ENnY2thIn7ZseMSs8XhQXc/DtS9Sa/G9T7QKZlbWSowGw
jCMBhBN3mhyiD1C6rwDJSIM1LpsNF0+Oya8So5g0+UXKhC2yqYF29lQGNXECJQ20/nhjnR4QfwVB
XdsfUni2bj8Morgx6o2lp9IfNZI9nUT2n6+VCICO108ZqFjDyKA0+gqhka9UBva2vqkGTmNnmomD
xsUhyi3WnZNJ5gLtXJ+/I0y3n5Tfc33e4D6U9XiEXaAtZpz0W1WnKYLSAE43qyLCEwFVy7ej+p+C
ckVqAfKZKYB4RHN0bJ11QplCaAkWxdg5GwlvLdhF3NGNSQu0dWBsHhYKFko3encFytkBbzfyU26D
SX17yEDeDvyfDV9RXe9kSBJTy5lcft4Uqk/amu8UIC3e3H5X/hVDxndX310I2QbrLA4ZHZJyMmXW
MIVJ/EV4xpSSGRvzZpdU+kUNINhuQeFHSVTt+sT7gAuDNL+ygFHv//7waRT8R4wHKuOnYRz9U/5a
eSCB+ODkFC0x1px3e9uoNEHN8oqaNDOrGkMRmEB+vvhbYOgjb/pxhk6odRhBBG8IYXR5hPfSQvTC
pfi3hfQJ3qNNoqHZ9FfR7183ndp0onxy0XzhTqkBg6pWZo+C0BzebqrPpbORwhDPloo9TIuXHfEn
lNCj7SM77CXzRwd6bgkc3TWgioM7aEKm09t7V01rR0/lnvwUtVRtxvcyOzLGukzLvqPJjokD1e/w
mQXpgIrUrkejNvtNEixMCI7/P/XJye6KA0rH0ZwGXMZH8nbxMK1P1EHLbLXEj/4rQIlj53RjlCME
dQ2IqXjPoVTYWjKPbNQDsVJPx3IAMDvVGWfGSgItClOyDZtO9KH8VQuQBY7GhPm1QCNXsAHLXIDp
EDLNuWdn9iA3WUjxZDrsuXGQPs6U2INHVt4XcNRv9RT1s7c8ypE5bbXLl0FKGNt28lJNezm79erb
F9a9CVavW2AdBHsu6EaxZRj2NZPEO1Lg89+ftqh/ACP1tEpCzi4SyzQH3j5czR5tzesbzZ8JFbHZ
h3Mrw3WC47n8l4bvpdCyIqhtMX9ZcutmrtSOc5Ll9G/lF26W1rwcdoBM7vyM3wW2TvokQ8mcug/J
Xx+8/VocjAUWLN8tWHQRxgM3jY1yjQPka3GNf/Y0xV4rGldSOBAZZmULNbos58Cez+UW8UDr8+gc
k8XAnB2M5WCfIxUCkO3LJtUXRGSQuv++JNuzhTNOK33dQbDY/EoAnap2YGhCH0RZ08QBy7mw8wtf
HBosAGput+Dsew08RV0zVELmhYJfC7C1KmzFYLaDXW7EQYbPC/ZxcSxKwuyvbBVwZac08Xqvx1Zw
DTzWqEC/XL7wiVzCbZiyB2Qli/Ufa5XoMlSKUrSDfazfqTLUVZpapUZFM4GTJ6DyIg8Y63Urm55Z
TytzYlTgJlHSfYkw1+vcJtIaeXD4jDW1gboorSXrgzQ0U/sfSKBbNKyVybpIiD/cvv7rHGjVv6nx
7Ru0UoL+KMZYtFINM1x7OBjC/178uoUG/y1gnLFLl11buQznpQ3PdLgUeKKs2XN/rdJ/FpEqazKb
lXO4EA1EGywvouND2m8WSxFhZi1Q/U8OsQ85NzVEGCryLhTP8RSZ295GOf4EeS86VBWPJw/+VdwQ
5K+MQt6MmzXNaPcoXMSP8QcYwNmhFQfCnx34FyrkqzI/WrsGVjtvLLL3Ibs+r6SPvtpmL6Rhz7p0
NT4U+OrqFlI3Vy8jxXA4v8tM8rTeZXuzpRpNatVVj0zjvdvgeQ2EcibcHc2TscrXPond5V47U2KZ
hpA6rUeVbbLu1ovAMsxna2aoa8riqRPkmyGW1iUD7Ed+0vC51DAsJY49g5eb/FJ7mRDNO6NuuBYu
yTSRH+BRTp5qxVsavIGLOoA3Z6vLRSV6bPTr+tZq6Eey/RLrgF7f3ma8+c/apYxNrUZ0fT7pIaPW
3dD+j0X+QbFZiX3boWTV61VRupahtv9Xife2cYDpbglfkzpHuEsulQX4zvMLJsHjSv80gM5fBmI9
28itjAAH1mmzeK6Bb7e6EblLM4Oi8FtURrzjApcfSQe1gEGgcRrJX5hbk2Ih6ENVljZfLNDNW5Ue
mLOmGh0kyBtlzoGDCFFNUT14TC/eEBe3tyhEnIfe2avS9eE9Qd2Eb6IjnOdQnxe2uNfHo5DCOiHc
kxaGFaPGQ60x0IywRnorRtB9xVAjUDElBOXvoT1tRwFN96qEYBtAZwZPM3CgO8X/QKzHHjLqbHU0
XBSdsoHRW1i/U5HV0VMcSATHyw+Zm9UXsYyUDCsd/u5+tRu97iYi+r/Rjr1jWgqwYkZREjXkyhPm
XlYFGfh2UcMDt9ReQmbR5PGBf8/aUdkIyRolyi2/XdNiAg6/5cXkkO1b/NMY4wgx4/I4hNWVuddk
SXbAPiDHgA7RbpfkdOKaMReJli8jzSftaJiVaMeQ5JislA+PYSGnchqE2TfP4tJQdeg2VFYaLvTP
5aX6PRUlIWdPy9pwgXHtNHDInTykb0aDKmEZUJ5ELprij0RSLOr7Chp6dFPQG/yURG9bv5/eGb9U
LtshKAM5l0ZjGhk5pyKqfOVss+iOaQn6rp2IqjWLHMdfm3ApVTojoV12Qh3wV49O1XjuMlPJrvEj
4g2NretSy3rOo+kv0fgMnqQTFWkOiYUySqbGj+UkBSuCE6CGUB7fAYtegPEkYN9t8pkKNWKBlzpj
Fyke4YlD3xf4hbQGQWCMQHL0+GpDX63qOy+ueclCnC2edxpPNNL6aY95birJ5+nQKD5LmlbVPQjw
+aJk4YR7I7OTP3+Syann979BmDdsME56tcK9/0K4KADDqud4twLGn+N9iOFSFhYNlUxoQV9oSWSU
jC1BfB/Tre1m2aYsTREv0Gjh6B7h/L+9GkgY9pIS/4Xx5Ud6AxofYSJ2O6Pi9L0drnbmYNAKCXqL
yUnfPEhVXkntOy5hdgTPECo4iXLe1l99GW4lOkrxa41Rc8gSkjCmC+1JCFCVrJ0UqCm2fKNLv1ef
du1Om4Vg9jirDjQJ31GSHiPktupZZsQLFDianUgFz0ugD9JykzbjEeQE2yP/c4Xk+ihAc7gPxhA2
Qzd8RESVbg+P6NR+hb6dv3TrdOqiVqXLjq/TPf3GrfrOrWs+8M1iJs3QEkQfdIzC8KcmRjg+dtKC
2bKWiZOhT/TAx9xDJx1UkcNZwKNxB150elG/NiXYN5faNPAdg5oHOt1LVPRruSKUlPIhKg4KfnvW
yzy9DFXCipxCLj8e+kmewpGwk8n1eI9opERpXDsGZMogaec3C24fVV3ZUki2IYPm8wpdgpe0s4e6
B4B905pchJqrlu/o370iLO5raO271yCooXnOkcE5bSKFfjwtAvf9/SoM9SgUrCZkSydKkRGPRE/y
2Pwu+yQbD4VyLbDU9v7n5+IpyxJVP6dIVcMbByU56eI7XqRvleLToTTFj1suHmQJ8WnoYEa0Klta
6QWwBRcYsV1Cts9Qrfhc7uaZDe9hxqgr22BvwDShJ+YWDTfrC8LWESFkM0OjWjs9Mnwnmr6Xq940
U49lG0ijAsHUZZVp9eloTexz70k5tr0rjfEnofiyraY4bFVh/hNJMDhwr7tXcK2nlT/gX14JaC7O
BaRj0Um1U/PMjbZsHsFgfhvoRHDE9CGQpqh5JRxqvnlHOR3AVSsCDdKXrhmrrsSvOYiufwX8Vbnh
btZUYQOi2hix+IeeoF3MHgtjhjDaDWxaiLSKfj5QThyRPiIorA6BkedBvD4KY/Bx3RbfO9nFOPfo
CxE4CYuS9M69wTixoLd4fi3nr/TGwFaoiWBK2SqZWxfBKk0z7uxd8wqGoMb+erhv7v4dB7NfNSps
0jiDXrXogtuYa4lismuUSB0BTH8idF+oldx+ClvEjh6PoAQq3MzwM43xxzDUjBgawkWEhU6ZY/gD
tl5F4VISNbJCirmKM3nknIYvx0g1WPlFETr87FXe+vcYxEcj9bYX51gpL8Tek8VxeK9ZrhOBYSiQ
G6NUtDR3vy5p3Ye76rWPRYjib9ugmKyrEiv+HOl/9oOOArtLG61PCGHH7PD2fLU+zCQzux8xWdNV
O4YQFTB1HUv0ej8F7PMxbOKYC4ty6xbDd+MUwb9/aaP5ZFPXRJSsfCmo7FP45/30hdM4TBrFA2TB
dWBN+7VkK9VVDHuvtPVbAXI9RSL5xBoLtXOwnHC9Lzob8FDefbZWfzZmIN1XcFLqQeOxpFhjvlWR
Qg5u7pRtHrfxDBHqGZaZ2Qdf/2tpPsWJ6yn7xVqkMcxCYCGQZjBOUtV66Pa1jw1AsjUELBH7ggk8
MYviLDMUQMxjYX/6/dW13a1ujTfLV4NqOtSdmVgN3rzUriIcZ6C+BysmtmEPi/rjjiA7mmf/m0Ax
fuiLU8KAjBje2OW1EPUWqn3nGvfiUGEgyPiaKQ2P097BHbT23TCJpDOa7QYX0L30GIhyhs9VCxVK
bs/2iK/Y+e5sGJ3i/+wzVkKvF5YSDWrBWph+etQW6G437xm1JtWj9a+hdLrzu7exFjsFV5fGnm6n
+3Oy52e/tO/uANirT4t3TYt/M3j4P4GMwCpilrMJ8ssnjYBYEbUGGsqtJqJaN1iSBT8m8ZJd4C4f
QuZBl0c3jeTcyveEzMw/0gwS8BHWclxamrujl8bKQirYgYfeVlk5Dcs52WdUblGnNFiQLjQ10TYE
JwrbpyOP7bwF6coZagN/PDj5QvBjlh5XH1HW5yFn8X2IeEp00Xj4w0PXWESsB9UKvvmj1AP+IZc1
cmd9cgiISROtZrVXl5sDWAPnplV0eCyio+dy3qUfogHpMhPVSjPge00yjE9moLEbQj/FmFbzfcj0
6DI5GRSeHOJUNuWjNAvMXissp1mcdS2nvXhsreok9NAxFI8EfIPNS42L750SO/0buUQar2S732l8
pRNiPYtacDqzb9Ns9INhDdPU7ptTZVy4uSfsbJX+VboOtWEv9wOiwqZWYr97L5N9Cvz64s+td5uh
2qoqF7PHr5aofbWJVBf5NUbUhaOubsaTH9s/r9zXGimJBzyfEX8DTmnSyLPh8cX1yl0NIPTmBrUa
fTWBdRxvJrtciJMopgvUlKshXtVnObPFuYcUWkleBGj2koElennn8qciQItCqLYwRAA4xELNu+G2
zwmLHpSkGBZFSAT5Uu1UE08T1R8IxODIWLmWsYTpSCel6LOkM0yQUEYlj8NCG5aAqfl86Hw2V0zv
FqUhB41bFgHo3Ls0w5D7iVxBhBY1KmF15eWMFL5gHst3iNqFX3F1YdCeHfPonMqn1y81h0trr1SY
tXk4uOmaEIKS39/DIQqMlT/8XWkExJN3I1v20DEVSdU/VfYKk6GNoIGJ3KaPTjHMEayTTtCBz+fz
TuYEMdeayNKQElmNfG5/Lx4Gc6CV3oKkgniapBgLnm1/qrUltBppYuDFtGk2RH5K3IMDGTma1e3k
QR/iYD2A7DBYpnEqYHZLOiMXNABe99XS4WmRv7mvmcK5PUW5ZnJ+WsxHCrQcrTxxzAYg4kgqRVqZ
jb35xpV4jOel7iPg9jaYWjTBxarh7kcy5AZSjN16oRchjkrGceb57LTdwN+6QbJCPfL87P4HKYSK
CGg/BrTKqO50bqXS0UngZBHRECQ4TJFBMBDhJH9xdh9ZVbQFsUyQcHjo+gRn3tuNHdk+QS/h3TEC
xgQ+DNQTdK7bBtxelBbNbmoyIwZ5de9/JQ8mY0sBfZPUVARerIvWN1YFxUV/eD4pM0uIuMUTDam6
yulBWpXm31dkDAqOfMqaNovRFpja3H+vrea3iGpign6Rx2bE9CCNTkL3DJp5szY9vSwiGMV7iEhu
SwRNUYZHoVl1bSrzAyfntKhYzN3ARsViq1WNnUBHHPAGQJ2CbNB766yb9oFh8WbEvOUaEeS76aja
LXqYKYgxukcQGHaOXV4TJR6N5m91LcpyKZkOFdP2ieDPGWqlGYv9MflOUtYAW0u3KTeVB3coMsUP
HBvKdJ9Ci7hPbcPVAzMl/8sNNaf+5ZOooZkcXLIWg/SISh+KGPz7lrWxeiT64vLW3KQorMSkbZcH
Bez4zSkAduBuOix52Xgyue76inu+8ljcNDGOjonday4hfRaJMJ3q1kuA0nnO/i2OO/M/MbkjHIw/
kXsx5AaXJMeTNkaMPj1iLVftVDPSeayCodtWH/5Xmzdg38hEJO/LC3aSTeTle+enHzwzbR+HuP1R
glsNcgFrDJDg7FPVHRRBBGTJ3VVnPbuyOZgzp06PXt2f5xg/XYWVvzTk7MW6DTmTjyaLEkxrUgeb
Glaf0eeu0yKItlAZcl8OghUpcUDqiS1u5MrkmlcrasVQwIZNopU0mbR20KE7AFbT38PYahd0DvPM
VYmcLHHiK2Nz7tmDbO91lZAeIHPDYhEbZXPxyVNGSMk9E5hH1OZ+91V1Gth4wrS7SozHveEu945G
n4hpCsHCHC+BD5RhgmGL24CT9BOFZs/EO0R6fJeJNhxQdDBkxKN08b3MfrXgS11wBuWwdD9kee62
s8d8LiRmX/F+Waf3R23aPlS5w+JxFa3BlNVkG96lt1XFwFHh70TiRXUdLpwKXM7JtnBjPwcmSGKo
eVMUPRq5nX85OvVnLi5IWe+NIHkfde7rU+R3QMVtnh8EloUJWUP8czjmBvS2jkQV2lqurXkdoU60
svWBvCYKxdJb2kmuXYtdkkYTJmH9S9U5oR9afz8LH2wCUKmJRK5hBbSmSoCCQwr5TuDj0uqp13ID
lKBF4Jt4HAnMKi9L3j51+Q0PIuq5pSkM5nd3Svgrx/Si8JqtWJYMxSlCC9aczVeg+4iIKxcAyVbJ
t8rSKuM5Uo3/jN0sMHediZ/MkmCfEWpz8eBy56kUb69EMxrH1MDOgX4pn4E66eZMohWGLWSIunW7
6ecGAgvqPPVnHfU/nKPPTkUEw1DtLSN4fAoX+fHhy0fG5yB2QC0skCVuyF8OB9BW1sTSX212aKOm
Kj+S3/g/twm8vz2BRHNl4NQgwvpywCSUs43+g7ryzm6LCr6rZmvexfNnXOkecxJax4kCl3G8kkrY
fycgRuijr3RYrKiBjzStsKo4RJjhrzomp2JZvst5Fq1XDc+T7TRaQMLOQSlzGG9OtlpA9uMjpWCu
2NX451xmz5VzqtW/BB+rK5p91sv0YE1DWWBZuVHKYFPJexffI2oZZrRLQkiSrplkULLMhoqzbZOg
nX4TRO4+4WNxhJf8LhgoSkUDeyPUx67vWPPxqi/9qlEXrwcu/L2s4ujJVZxC36e6drINHq+4dlR1
5XaGDtpkfmAJtNRVhWRj4TmbKxgSBav59hqQkuJ7agbm5j7II8KokE2cvbP0GPaRkQP/59rPn2Md
ZynnuM+qJ4Vg+rYKRe5FaX1/zLWgg9YCy2/ExYFF+v2gMDz5tRXJ8DPOKyxOjseXnNEDRzpMdl7p
cXjkBnyTIMYCSBg44Ug6k5bSMq0g5ikIa7O9Ox2hsd/EXp1WUT414YUEERqFYR+eivN3+qU25Exk
NB6+3euIHxu1lE4WCleWynIJuxaYVdfKR6mn2klvm1k9+OE3kMZ+9ga0vkq0GRc8eg5Wj9UBe15q
PIepU0NtdieirigFA+0zohM/2o/XMIm7vO+PZhQttj2H+t+2e45EW9QZcT2WUdoyGv+e/2mc73hC
niBP6pLXzUS2c4+gQOCszjdNKo40l08NkZS5LparW4P7kcRbq8CKF3Rxj2AS1ggzqyx/E6VqriFH
EqOgEI4Vr6JWBEXYLdAvN6jmRHN3foKb3DTjYqImDQ+SNNp3qZfDunJKFXVK2wWqVqmAAagdPSUc
JoHcsN4Ub+O7ax2pXIiNq18GlvAS5lkVxWtZEvIn7erFqfW6fkhpSLTlnaYkBJRrsp/pfqwwQa/T
nBa2VomJylYrVAZVCAJfh2C4XW1l3yAwBhAtoiRyJPWB5HrW01+Pibhkz90Em7i/fumtkKFMw+lL
ABEV7m9VmZ5b5CJsI3LVlOl6FHkePU01zNPQbWOgMaunxjteki0do8PQl4HJOE+kYL7udRGJ9kug
/5AbiwJqlJx7MTMeWlEZmh2sJlO7KJSD/CQJCGUaetqVVXbSqiMqO3G4rXvx8hFRBjDuzyYsOoY6
vBzhT2ylNsZK6U0LukRQ2bAsuiOeBX7tc7IindBEWHCyoN6J0ptMID2tTJ0keHib84Y4j7F5hZbc
Q/L4iANxjZg9hfiiKERmNTbZmBzxDiMQnUQgkfSBrm5WIBYtSHCuMwo8KItOKw5iMgYYFikWAHcQ
rHFAl8thvIm5z1VJcdILSXjQIfNysBkFVO+3F3cRMu5iaOQcfHlnJi+cjGgpv1yVlxmhrZqo3tg7
FL4Zu++FPT+HiQRHs5AlF1o3v/P2Nc+THNZjkwEJxIY5GwdUDuQwtbhs3hlr1r/kRQ1+G2zEBb4m
oN8Fw4V4zrCyi3ppzdaEgiYVHkfjFLpL0DgRGuFN+x6e1CrxivLtIF7X8EzmGqAaVKcNeAsS9Ddk
5RD+ysCDVdlS6PNmqxvIM9iRisRldbf7nKGPTiy9hJL/pVaxs7asY8N9+Hu3MzULQLsgCtBkgMG0
ZzQ35ZaoK+nku4vFZPm7hOjHr3mPWiXPaKeVAgzvLY8KMHWZc+w0WxylcfwEFVfQLjzvlZnwVkGx
sOLvWPjN/bFFcvEWObhhoUQpUl8r6K6e0jNYdwlkhHOL28cqYobxswu1tGYkCegD1J311PzjBNLR
iZo/MLrTHHED+MejIdnt7Zgpy9FRxHCtu8GTBlsbUZXYe4enDWRiuH2UUn0qDWsJkPVcHNXjWXu3
+nNFGdaonBTyzGRPFCbTPFHRu0ffCZZr29uG7qqJXMSU2zzlZnHythZzr9Ku2t0n3kXPolvCPRtE
g+s+cpQBoqkn3cCS7Hig+ZkktlzMBxbt3s+L8SHGI19eSJZTwALHxFymjig02PdKjpMWqTNojKMp
WXnvAlC7mg602Rl1aOC2LTaDFpAnyhOpXdNLiqCEAjbf2UTQLMsYBpZZt5zqTMyhwwN7J3z2A9xG
Us+RYHNRjLv8JTFda1LaSHEurrLfpswRj60TvIjGZ9FBMvfSaGv74nxFwReWzU3lXRmjyhHFyX+P
UFji2/awdOqauZfo10I+ed6mjR8+Nkacxwv+js1JKzZOsrNFOEJ6NeH7t0z2ffDcNVudW+GtJqU4
QR1w79cxacS4d3buYPMFKX2yDU+1LV9rRcLqmqPl3xG8sokqmTkpFlrkd+wabcB6TFU1eRnMBZPi
5Vm2T/mG2qrM6I1aAkuiXCpluotkMIsdREqVwk3ZpzuT1L/K4OrSgW43pxhu+IwS66B03RcCU0d/
Fm+KChWJdlNX9KChrueirt7JkyHk6SNZ/4Upv669dfL4jq33+ghByKnbSEKkvXxO9O1ZCEOWjOPg
Tztx6LZjtvaR1aLrD1rNJ1kjL8gUc79LNfFIlsapio7i/nww71N2Z1LP/rKGK0pbspOojRp4wPPA
tg+6up/dcPNZOMtHyjphbe9LXbSOA7MpeNsjM9VpOd4fWN6Jrz0lnew0fJ55OiUFEKjhJXY6ID3P
ht6DXAI0SxObaqXKWFeGdDiAAzSKgERVW0TJGGXlyha/Y3BZQEQpBHs38AnwEn3q60upjK2phAar
pYlCaD0sw0m87L005QB24V3R1XXDkDeIVAlKMOjxZ6LVUvysxwXMqJWvfDREdacxgiSyq7zCVCts
tfA/yHVraWkwzoarywpqP7AcSxbRQGQQIjBM1CvUriAqJNE6yQiekXi1eh4+niWOcMhVxO0sJ9UM
SCAQCcBWYHcw6uVzJBPpajQpa5BRwiBshJ1Mj/PNNUp25du+88TOpGnag0xjgIQJ54ZTfrfX7Rbh
sf/MGE7UgWwQy1k+QI0LxPrhrLln+GX1MYWwtyfCodGUl6/LJvS2J2fMsdPCpV0t8SyRiUgigfQQ
vzUqgNAxW5LXiDSL/TeuGmI8GkMsofyud6EkoDDS1ZoKoduDDWjpbrhlJ6+bbqKAwa3MfWhu53db
qlX9jLZ0FrQBpkUqcyXQh5Aqr6M2fvUsYMSjpZ5tP2wgOjLKflHCaAWAjeausUOEfhIajNvLiKHh
r0SpGYbqpBE19g86pEVKjlt4YGjIMC0duX8O2GSssu/KzCvKHyU87hnU8Ia7U6ureK0yJSFpeMdm
oUeDsUid6F+GR30LZ8yOVA+27q7Rxl295XjAprCJSoEEIC88qq1KceJ9Jr7t8P61Qudw5TlR88Ai
zc4KRS1FH2HzuehmDs9HqvRsFCotAvhBJCudWTuKXSwkb1sDA9gttJ4lj5Dz4KJxgNI4Y5r3m7XG
qExy2wsO0ZiQyvuaJIfHDnflyXJ17QHruAT2z7hdjAMlbhRez2qxHMGbJlbjo7JLnFfr5p0uX5si
3JpI8htXW4JuY7EUsTVIUGisLOYVBF7vWbNLQljPaKTYejR6ogoepF2sJR6RQgQzt/9xFJHGh2S5
mLuwOdQi0kG5SvmLjJT+GQwTdc3esArgVYPKUlzynqcHFEPbIXAl6+rf38/Uw9Wo6rTJi6zHIV1d
Pve8Y28UO3YknsCMaES8m1NkcCW+3fWTswoe0cZUuTcFl6ZqNxgFzYIwi1pI4Kns7ckLlSxGF5MT
8ZDX/sBN4qzIDkZt1FOYqCiJX66btYWb7tew5OiJFNuVaYSRxogrKxQOcy4POvdEZkVrxRRV6ONc
tPgkcfjejurRaOIkbtc9XkgBoTbJlAiPL4MR+wZmgoEMZ+Lu8OtS148+b1CJ/80NuQ9F+5chDUf5
PrTZfPSPjR2Y9LF7KrmVbxabU04Xv79DOs+/aThJZuvZTdRRrpyo1XxvofySR7+JEoXd4Cyf4ZLG
2wkq9B0WYy5SOPsSoR8CJT3rSO6BGRJZrSILGw5R0e33KXe4LgbJbr9A0QWE5ATZGZYcUG5kk3Fn
Pjl57wehdke/Twu/qJYYUxJlq037UAlTuGVc65JQ9usirdFEbnd/YhS5dC+TOX/xw/fr66aE9ytG
8oV/yJe5cNgcObVywHjy8BUAW5H/NH2YWME+f6gv5aDh+2d0n3Ja4i0xrq9IOamVOz8cgUW2fBO7
LZrcPhad86Xjd3SMcXFHkUZGAnF5Pidb3hhf6DjcHhcBfxgeDApCnRIY6bnptvjrPYtWmr3znkdY
Wsmam57UwQLH5F84coTkmqhXPwxLR6+RLMlJ0tXXxeYXoVjRIobso7qvzciU34s5MKLxBtH9ycS3
8EZ4JFyOwVg+YgJREU6FRKVjiS4dL4JHYxQd30Fw26s72OIwwHNpczd0gSFonMsl10r4VKD1Y7Tj
+O8e+EEnTo/jXK7zyAxSnMgn9ylmRicjvFnwDTlw0IswjWyM7Ze9EKiGVHY1f322ePu4/wQrHZyh
nFQBw6411EXdCkSDQxYP5/RYitZ/hWZtpkEovCFWqOsbyUTbSn06b7MEFPpUua5ehfN+eszcbuM2
uf+fei9fKj/nnDMXk45ORwg3Bwqfbtahj2nH82YpQy2JyWzpR538Hd59Urwaazpceqdz1zieUMqP
kyH6W/nXu07dI/MIAFvP9aA+iAw+oi2dk1QpyQq+oi9+SXqmcSDBQLzUmZ/AazrO8nw/Ze8qJeRV
dLRQqaiyagsa46pHhRPb4wZFkjo4ujqls+8k+EL8hPQnZ/9nZ3MSWx5fS0JrRwnWSjnDuaFOo0Yh
3HqATa9nNck+YhT939f+TqRZfnRmddV4KKgubtCzAjwGyvBTpyELt0pMEV1V70BTKKeHrdorqTP7
du9vncmrsTK7O1SIY01vpvbyZE9QhbPgcuuM2JBEfoa5GcIgAALykmnU+7GTt+UExwxCcEBUggjy
P626KpzrgLnfnKogs3in9uwSs4MvEb7oeAzyEf0nLlEt0zZvttcutoE5EyFPpZBQmCCeNgea+dIs
JMyDYonvl06cmbQbIQjWCt6pKbREvUK18ZEVnhd7MUWEjwefgkzoph3Rz5vD213JMw7bC/PtMIVT
Fwa44tMkb0lXYRH1QmGRfP7k+v+hbi5FOASf1hnMn2YbfJ5fPEQE4c/e9mlpBr6FZI1+yvOsB5F2
SP/b6ps+F5hEZ1J4kIhniKcoIPh2K/mP/ELRDv2b1NBDQhqadok+o7iPpyf9s1POHbjyoTnM48v8
eJRAyVAIdn6xsCnQOGay8Stsn41MnSr4yWBcQ5UEKseAidIeqQB6HyvO1Fb95CCTGO0Opagf+r55
9izQ6OBvPR0Oc9P5c4gipCkz9kMWrz1OwKnfBTqzvjX0k5Zbtn00YMBV8wci8bUCaACj/lbsXHAv
Hh59LLFmb4JyZnDQAZJS+/YO0r3uUxLhjP/HKlXCVjbWihsS7FLgtpN3Fnk42Vj8kXar0x1hH/EX
MQ7HHKlvhOr9G0ZZgDUyuCLzs0EoUSVBV4OantgMvdQkXnGJWNlQGkxs6x0IWrhp1oId8YBS0fA+
Z2iihdiIhM0qZ0E/bE8OdBHKu/EJWr+/n02kOx4WQFba4GsqPg6zz901CDRvvs6eYsbHhiWnxqD0
XjoCPgXB++aHzu9KXm4Zni05ewHunMMDS/HPeGVsTYauRMkxobHAN8J1tGyfd3G1isNQM6WH91zB
WQkQ6cVO9QsKWVrr4rovWr1TyOFULL8zivLj03OAI+qH8O/3rltszESbyIbO8V1BE3HnPvXylv+B
QgZf9jl5rkRpiLO3JaGL4HZ/rSky1r/nyshxLCziH0oRtua5Fb8m21Ra7dCwHGEZNmb73eJk1Fcu
w/SOv2OoX5d6IhthQPlBibCgiHfQpHq9QAXKdPlylNduavJ3CVvqOXd46b+ukWng43xB+kL7fvEG
u9TSIchca/lF5ydvzlN6ADATeNcX6h+VH5+LG8yJMrqUNcqVMJXyp+YzC2QGhLcW6SpyYmfxQH1t
u3UajLLHal1ZVy8VJUzbFivvTGlsTqPb5emD06o2WHsD/8jFrIHoZ3yASoPm20GWnqIffUEbFmdS
j7GKwasRs/+N1pC8HFs7HjVDWlVgzr9l98pMfDD0M5fiWV6v8XCK/ty4t7tb+UmIwocpfQ+lnGPH
FM3rEIX6H2lcw1LnE7xcY6iy9P4CiN+8YKHNvXN1Ru4NwEixe/Okotz3zLggcRUsrlA3BcPwsE6h
g1u3hSAW4yYnd2UkUq26VJb44lGUhnVkfBMV7DqDuqV/x5fQwRXtoeNXai6dzP/pZ95J2QidK7Q7
p3ocsbboxbcNjoJRd9Eg/XoJmOxgzU/aEgcZ1rHkZ+/wy827rrAlt5EpKI6+DHK/d3yrMZRj+gV7
7j0LJr/ntm01zoseChYjF231eKXY4KeFmHAUtLqD0VLK+JS2SaekcMzggzipLp7HU61mc+iY4L66
qHK6ji5sSoWhM0sUTH9+pTi5K9shFg6/Z1RtjQ32n6FnPXOA0ZqQfzrzeHdLsYCsx7HFOmbtsSpp
ONztwLL+0xEPgCuImu+VlRMI4Wl1pHWDNLnB3BKJz+FJdBICoBNUTJVep2LoO7xrcQOltRCJM5HK
AlZtbxDTsUKG+03voBIHFrTODRjPbeK3EmQt3XgGIbzbjmTyU41o5vjwEjgIOaMbry0rTXD0uGWg
hsumkyB/qzPR7tNhexr4JqzArkcpnCKpWwRGkCtiw82W/TQIbuquWbsO14c64+t5Odg9bZ00gNXp
l3LpXKGen/XudXve1PbQoOxdWQFFUEgINQFIpxOfjOUVqEA52/3Zyura8FUBfMmQyyVZTd1VsvUF
EHbFq8DqrCahutnzw3jLpFBI/ees/1Tv3cCfb3+7FiXq17ErX5Fiq9oNOzx54lpaSc1H5BtvzzY8
09seot1+QLIcZ8H4cT34633mb2LmZdTjeDd6bVj7Lmq5oQaQ0Zzsp0QLFUot9AeF1gE/XSQzGnpN
sMItDI7oAvSpyVo0KLK0i8qfw62Tw/qL2AteJV6+knk0F0VA+rOudgzYjNbiVy/mMe/K9XYTCBpP
fgQDAlOdj/6b24RDMX3R9zA5RasvgAgVdCzXsYFLEgpb36+ELpP+RJr9x17EtnZ0i+ZZqXcVrcW8
GPNvnzge++pHTud8/5W672MN3Wy/bOfNf9/Ay8ToPB+mghGOGlAEUZATiHkImnqHRt9gUKiINq+5
+LOo8fXKGL70bDwlEWH72CEZEkp21nPY5xfsFvVwERc8ITAtrTC4LbQXK4yYYSs+s2JfUinVWUIE
edpL6+CarENk+WdaMoHRvUpH/luIMrXYdP4n9q0aBSP5uuaNPTdyq/KPf2ZAutZ02MajnSieIBCr
SXy72bZcdsaw9m0VzQOjPyRfVq+41+nDiYTyCkV2axli29KVv88zwCr0EqfNsUeGw+kNAOhr72N5
Jkp1CWj9rXZEQFMoT19KPQhY7BcbDQSi/4fs8k+20soOL9vSH29P/WGdzV5VF2Hqq97qnX8SJ//m
J2rGzH/EwGQYCSEM7kyhTeKRMm4sEc7v4yEwjKVdoMrKGZ8DUFuBvsHtRfOj8Xz1+VM9zAnOTYIB
okqCzK4clIfnWUtL0WZleTonirf1hVtdP2RN8Fob4vN7aCSLzuUvoWSxTul6qliXYtnsUrdCGpuY
ibbDC50N0tv6nTfhhYxUpzZCNbA3Q0Qpq1n7IH8YcSVDKye55bz3YuFNClSfxjZrZCOSaeDcOE6O
c7uePgt3xno4Ncn10XxBiG1M5hR9Uyd5gjIUzLvddEQ4HwmjLw14FTieXAMs2kO7VozkiNqMwdwA
pcETjS1Nchbd4UTJeTXMmRwbsjxWm/CztlQgIwpVkLcWKBAboDE9bfI+P3T7zXo00Mvsr7ER8Emj
K5N0JFRcX5BC2LFkhXbL8K3r5SEh9qtetwfyUO9ui3xqQUw1pkgbf8HqVtKtB6Hak9OgnqYmeFyr
WG6yacEGRasIbx4Br01JOi75qoFYK2pYTawtK8IUA6BC75sA/0lxi+8VKUg2wqUuCnpf8Jb4cnYI
cpiBF6baPtIXqpMG0hYvdLes0qVn8DfrIeRtdh/Gv09O6rltLYU9WDHYy1pI+atitrShM9GQULdx
UdQDueKJ3F6ynMGrZYCYyOB53VePNW5zRgWjgImYuA46c40vmxehOZ3yeTwJuLKmRw6jLLdImCH7
O2TZ+/ya74hEUWUoL9rt9dwn0DzUzssxniCcmCefywu0Xwgud3tM0lqhGxAVBN0dBeaHr78V+QYo
EH2gniR7EVbcxJUnooxodXT76TnkTKPlOGpnltKes8jmDQBOajnAejfEJRyRN9hrUWhGmseUQxqY
EN3nT2nadG/en29kKAWgvpSMgcAznUdtZ1HbeC/of80JXztVRgo2TO5dNMhjGA86mWCCgKVeCw89
RIRlE1FOLxgGwMAEzqHtut7FYx6FpJavXXFslWhT6RcuJagz5Ju17iit1KFSvpnzobZ0ZamCSZGL
VBzJclPZqmYmlmLpUocY4xHFmPTae2LMch3XXQznJzhA0FjTQ0LzRXfK08cIU+hF4IkNh0ka5tu3
JSG06bhQ0atyk4YXc87FluQFghXbJaEdmnwmC9IxKm0Esubok7Y5Es7v9TPE8/RXdNWm48C2XV1Z
dJinvgvOVJEqe65pRBqeGHov0iQGJ8rKO6TyKy5iVpwwXWrGu2CUs43a8SmqDAVi1G37H1Prb7sh
r5mNB5jVRJSOHGtywD2PoNwN+FaMo4iMIkj5+3dJcm2NTfZ0TP13OO7cTBsCPOjFaAp6XcusyQZ5
ZjCIaPSTprMcka8md08hgFR2GXBbzb9ZaoM2hiOJQkHaMwDkagKuHqFpQ2oUJomH45pmkScpVTJ0
+mRRVs3+2K0KC4tqIgEFjAbm2fuGv5m8tpTMscXoRN2O1bFg59niIRdxrosbPlontJAHx/n4NS0N
rVDvf6ri5rckG0BMAbFU6+wGCq9dWOGbkZJzmmcdCsDnMOUKKI21z9AoabYArVRH9+voqzdFaooN
XUUAbq3/BsABYZ9s+NdTO/AHa1ex44HHltEynoeiYFxSOyDOULMDyV+4I4BYWjMlCdfu+q+Nj21G
/y/+J5LE390Alv49buh5RdMgi9HBhYXxhNq+G8ST7tf/KHdX54YQ+FhlUSQr8dd6ShpfF0meDVaQ
aM35fTAMQx9UyZwrrX3vEmCFUd+4gndiz+zaIosYT1OX1T7ZHOiNJD5+i9iVaKCHJ/QefjuLkaMk
xD4SroKUxqC+pT/rQELFohNPchT4qbUUmhVfmAMFfG8tvXRyvak5US3EkgbMhr8vBttNna/R8ZdM
C+k9rxh1SbhrpY0fe7/YferAJwWVrGYIvKGlAvm1PXMFGjZnpbRN+LvH+xsFToAK3siNrgXwmdl+
272o/Uw1sC3btbaPe81ASL50AKrwh+znIWhsnom1+BV7kniaEvXYHV1cySPRAsFgoPYIPgDf6DU3
U3mR11e/gToa9L44gfVPYc7e/oKPcqAXkfQmZhPAM8JJf8LBGtVt359+9Cx5Ood+5WZ8cut0OORw
t2zpTeajYA+8a5C6BftVROfe3U29Owsol58e+3uiVGuP+uuJ8UMNnL9kL7EwRU/lzIoiHzdTxGf8
32GCMMjIbf5D4YOkR25dQCHepC0GxnglBOjy4/kkETKeLK/sLkYvNf4Fqr1tve0UoeB+biUs++iz
cIoidLONe15jcEJJncs0JuyCRCSKASFRCWkHnKYRAynA38AihT8fWIKV4BgzKJ3T61XC578MhXF6
keYF4L7qT1PCbYqPhvT0gSgEKmpN2Z5xTr9rELwwHVCFbmO0bjGqFYFqFvJbOrW3ksaCok0kzD3o
OBOEs+XQcLtxBL1AiBhR1cHDWLJvM5jk7IFHH37Fp3uVppVuteEpt8Afhwod+gcsHiK8Ct7nLZMy
ig7rRRLE8ZSxRnTBkYo6ij5+oZtugDiIblwhsHuh/99KSXy7LMEmGYdkDAc1iekj1tAxAiFE0G4E
2aSBoDkglat5KqyNTlxV947N6GDwJvklLtSLgxfm+FoZYwghA0WQS44QgYRIimeOg65W4Pk6W4hK
kcJASHLVL/VHJL5U5+p0yaf3W5fnFGXvO1Xht28FsnUHR4HMZFXMXTVsEdMftV2Q6e9tsFXPNO/v
/xL5N75JBiO4xhwEU0l0kKOEykfHIiASxxTRgPgQ5ZInWVC39ERYPe0xPl/7zvt+xkwvUR/1na+D
9RzJiGNk8DrgA+/6l8swjIRqsHB17qdWyP4skoBlaNR7VOs4Yx6NCcnoZIjij/4hKNcJBjUh+w4H
zC9Wk5vBbOj8tsPfo4HNJz2IM5WYHkE/juSLmmaFmF1CUw99WZ4SijSsPsYb7j1x/uCkDPd1qC7H
8xffKSEdXs+f74cLU5dDL0hp+R4J1wrzyFL4UpVheliX1XQl01+4dIFvOaABjcUb2quWLf1WEgqK
jIQQAZVo4PkXsBGl0BAB5Y6IlPCrviCKhd42UTX1OOEZfGV8ahL50AQICoRgIA0RS65HI93a27Qe
35HywkqnhO1KuQXA2eaMKhYupnDLUgD6icU29QZYtbUltqnpZMrx/7u7peHu+szBrQCmpT+mSZsG
EmSCPurdp7oJsO09pQIMf7DBGLAwzJECEd2JyR5BBeRqoM4Yt5LmwGdtrtGbcfRcYgxAmdA0l+ku
EA2UUmbPV6XZzha+N6DOW+llTl4UrOOsBNVP8IwAroQXI2UZk62lf/wqGGY23A4wpJx8TxvRcGuq
Fxi57tu0tLoR7lkhtyeiv3hN2rAkmKwSCUxadBuD9Sbu0aanlV1kk/qLPSoK2fd9YPLF/K+X34S+
sORvfE4EBO+3dHhzetYXCM+yYVwOwl36W0aGOTCw6SFjrveleTSePJUUgOhNmTYs7OAOfpiEVNDP
z0lPxmlNEcxbySt8m/57jLTOswyV51QsdckKxnDLVW0UAy8NQsIiuoRzSavWCPogd86Gz4VH8emF
e3zxNXYCSH26CfyjgXe2iEJBzaoGjB6n59Ty0S8p58hYhoiNP4zVRlxjEuIfZ3+7OdW5bb+9GRX6
NA/uTzVdIcR6bIh54Klsr2pvUxTjV1TLvZtIQrjD831mTap4yRjnz65JHamkHzbYi/UuEsRwfhpS
n30XcIqgAH0K+b+9bD2A3SOngmz3f3m7pXiincSeHo9mnquc8zMob3vBJKkHWzt3GeS/G8/1kQaE
YGsMYWyMuMBvDUHZiZS7ZNtoYByb8WEwGNbj29fDQKNPRoNpx0spT7TYK11yAny5RP4GKBDvKFZ8
dMOuhv1Q96ttF5ScS4N6+OKHrxqjJADhn6yGdnbRCnD3wOly8hooY0j2/4WwOdhijIb58XmZA9N1
ZRuQeYOaRTyGc3VH9u65PXMnieuckTpXo8dcxf7JahnAzl5/OqoqjOAtk6gvOs9Ku2x0XWCc+86h
weKmsnxPl/nKFKDBUIDF31tz/NAQHesLDbXHXpUTHXBeYXHSpCbpuhRnOyAXlXiug+7Ougnj1MSU
2a0BDFwl6LMYT2CqTvlVs8zXlMe6OB3knfjBbg7HrgOjwSXO4vakQbVWyFkQXAFQZVZi92RkIw2v
1ujLVXbBHJgsQQ0k59iKAgIemZeltduoz9vdpL0/yJnhlyNU5xFOMddoBvz+u6iNEP16oFARvdWy
479O0117m6upmfmEln0MbCXG+4/rxM2ntQgr2yWy7ttsw/3lCYrQWE0fYeXcZBBSKFwjPFdN4r2T
2APZ6QfUKUSspaCECw/zDasEXuqeRAhUzha837NmB7aixcNM9RHjle+zjCUpuktCz7EnhlArAtV5
mJxbAPQKufA1FlQI29mZ6VbGvs2UE4u+4T/MdAF47qyFC3ffGIqd4Dahx6B+jVzoyIkc6/6Z1Mba
kWo8vifjPlPcM7pzP9yhLm3GAhe15Ez14J9+TpWN34+7Mm6mlIepz0cq18gRFPA6SqVfIdrYKAHm
/ynzjUGE3pQ/9EuQtRz7LIIfxQFZbv7v4kgL3CK1Lj/IOMJHVNAeUiEFcKc9AUbOdlq7u4jXiivx
5ZTzAFcmyxIa031xF6T4+fFjH5gSL/i3OsYz6uZCHs62AKG3WCPbpqwviTsBt0GqruhkcfGFGbLJ
vsMmqC7voqX1h28qDjk54YvqHy9j06cf1d5cGDG2c3CYaK3kySaR3b8eeQf8TQLkuU++NX3OkR8e
z8zoP0rjlnyj/SGEAJDyjQOK4HRp6wGTCi8hfaH+ulPx6r4SvZHD/FhenX3zcMNKEoWsoxZmHDBG
mLzkqw/mlBYMA7BXSQiV39Q4d5jUTjpC2EZHo5FimZgEIe1JBsR54AS41GK/8q75PCDBlRZcJpKL
taPbd05wG8gqB2W6ZicNxz0IOM9TvkuAAejidE5eGY2mvBpV2SragfkKXKanpjQkD4FGRluTLGDh
S7kMxTIdDwo6AtnLCnzoqpta1zkwuPYykMJknSH2tVWabCjoyvQSaq17jh1cRzgnrsBANBbefZFl
I7UIhH1O7+dzSzhFH68yYesEQve91jrqwtbg8FiOSd1g+aaSxjEHDwMJaW9ZPsHzlmQkCJKKmqUy
c1bxy4+aUNaxDM2GfGVqbY9UM0isirHUBcqLixXP7YmWNu3b63eCXe4Ilxa8WKs6PYhiiXQo48+5
PZLvhzh42hBq339HudtkWBrSE67tgMPAOJbaDwAQ25nhBVX8Kj5p3QcHoEyDsjBI5ABcspYHAzW9
nimZ7Ht/1ykYCCe5ll+jt1os0y/JUweQEz8f/Y/EhUCMvEv5vnvC0EyB3c/mGfSAMaUxpR28RFd3
k9ald6eV6jS13V1NzvrPqVKPbtO+OQq5E5YgJNvgUfnzvr2T88P6Cdc2QY6z/2PkHd1P+ljfPpHT
1noPoseBaTxiEL7CINmnCQGhcnJlh8bD4U5YkZDhZ2hnIFsdWVkQ+lqJCFm71LOEoPFuDuDHFMT3
qtS4KqTyKtKSdN3y2pNfrS2Q7hKoBk5Kt32jBMppgidQMsPl5THGbWcN0NX6NmGcs0RdLPH05Nce
lalP4HrLublludaW6y0j8kYaQReoKu7BGnQWsyHeZ5W923dIUvnGhJEGqdUv1e81PGI3n8HaGS31
zbS/6Ogc6qSxEt/+vTJh/y39YQdgFbU1F6l9UxIkJCj/Iyy3vKtFhKsTfP/7i7RiM5+Ke8B11zQl
4ZHNgEundidv9V81ZqlZgmHiRlIJki0RCK9nTfj1McSUv4byPVcgxmWjNEdDlkMJb7SXIdQMfH1p
h6Tu6/PIkzzQt2Z3Dl+1TjGspZgaLamAPQFj5+Qct5vGFMzM9ST7NTHUaTgWMOKPGIQHChxR31bv
WRsxtlnEDHsiMls1xns+bX1qTREP8nQg5i7W4p93+llcLXMNUJZdPN7A43nKatiHbO6NWR+yXZZR
CAfNMA6RPvQEeR0YxYZ6DJSFhtnKP5PcUHRBqpQ+XaOTC/jbH5/OwjF1FREQE2PjCHfGfHti5Jnj
+2oodcHOXFbLQnO3JyZx/L2IX96VSyWeG1+dY7VDQC94dy6gvgAG2Hzx8OlB9y3wnHpsXu86TrB7
6WZAwTAGaiEMDh+JVBp239HBNMDD6w04jRa/Q1rJS/ON/26NKnoebWUeTFFSLv68HWch+1uVR77O
mrkFWhmDcUFEPvj4w24HK/zUsJ3esHBn83cCNa7RdPvqIOipMp6Ri1egjL+tjYISUghXrBG+Cc0O
wEP9+A1+JLMWkDZORhGONTMKOM0htNudoPBSTmW0DERGrUfqfg4kDwrZbBKmZta2iMzhuQNwI5qD
qpxRYekKJJTcrznJqiOqNA7AH1wTBPm2Fth81N64x3nUTRsenbQTz606e9+BgfHDkq93eCMddbDt
dirL6UthCB7YXsn/p/rxZKCzMavJYQxCYT7/BVGYVozaK1fG3FtxgnO+GNgEAnnsNF+3W96Mliak
BppXk7gnMEstjaR/dKYbrvF/BJ1a3UNkGpgcqMY6IHqDE8ghWkT3wGEm2Q9p7MxrLarTRIb7TM+b
PXRsCq+WsXzqeXlQy5U2LvoeJKaXVWA8GNjb+0cdqf0iYMPP0EJBgx6CD+9P3OTFILFBOLiCr9vg
XSmw++7nWlRr6qzLP4l2di4rFcVzTTX6j0oknK5ZJawYzYVvVSbiNBCUsk8oJaGfYGQ4FJMuvwwx
scl3mDu48hfMSIxRj/BWbbYSJ0X+DQwTHYwDRgkGtDkuzJVUEr+0jvoFh7HxOsTZkMMvmij+Rx9T
9GasibJ+66lLDnD1yDbqfDXyJtMTv0Ub0QMm2gluQlvRBionBuiYF4elEdqfteAMG8BTxkj4OZ5R
6s/QkRojJY93tvqD3n9dXKx9yeHvqU1MNAnv93vzTv54geomdwfLmqXE3E/dbo2Ni0cmVgrRh4eD
expA5p/Af9b2vaIDimHbihrV5IZ5k2wxmdGVKADyDszgeRSKkCYjxOchlEpjICneANxQjhipKvFu
odOUyCPEyPzmGVo41ZSDi0FqSVgju7WDU7JW/DmW+XPvVk+ujBod36W/aKb4OjNFEZolX43WZ7M0
mnIiTKZ13qbR8prObr+LQJW1vFnVMEZKi8mH71DxT3APNuehMqxKftwSbP2Q0MntsHq4Pq/YYdOi
lCLrYUOhcOGwhWJKc6HVzHZon9tJ3u0toTFFmB0qyhlZGDa1jzs6brBGnd4v3PMYdpzWU7XLQ7F3
afqU4IgnNElcX4tKZHaWj4hHeb9EU0of2yQeLFn7YM3W6tUOSlhRrgj5q2Suu5QQO4kSkPafS3uw
yxkB188xm/Yqakkv1qclKIRAxBiNZWfMtRaGTFzd3D0K13aYtJBYc5Ey/P2XvQ3vz6ZN0qh6/45R
scFeHHLkgL0Sg7TAt/EAXjkFMSqQZOCfpKVDOYyLFaIU3QQPBxfEp1wXuaxcHqgvPkhtI9IQ3ynY
nhpjyqPY4hlPPlX9AkhoHV7/4JJn/VRZqRUsTo/8d2LUV7SrjwPtS/TINruH2/WnYYvcQOtisxHk
NrdPKeJWw7ccdiIDxWliwXTX6yL2JwXDR6bJYhNr9WAmhdGzJCjTFg+rAVuEDk7nKnibJFnGYPMl
hrzdJHadDju+CV4yrosGLHBXgza7tla0CCCTrtrbNfYLqdRC3nQLKxeFMa3AdoCnQWAMsQOM14DY
CWeGib4+xvG7pkuSF4ksrwH37/tb3CwnULVs48ovNoC0wetC1jZtk+vjqnkOLDUNsJfbzTBUNFVa
0KCwts8E2IOxc0Xr+I9f5+IOWn+rLr/dN7DdXSJ20jJlc80SaxiZogufBOdxxhqxZcYxcqTqb7rn
0kc7fo2DNvaRn7GMofUZp/CBlOxlqIMRXIS1DuZy23J3ylJHvrvlEDmXCzLt77vQ6xWkxUOUG5vh
5tRwB3JnyQ1UBxGGjV/Sxji6iwIR90YjbEenSmN/b+DrxEpZpJ4Z11XQHPfCGToK8ifVIwSOO4nU
23vTdeScnbHgaVSyBkSKWIUpEGHVVlXsPuELmPOj/nWi/2QzLsJmqo3FyeCsTTMi0kInxtw2Nz4V
d3whT7R1e2Q5LyHczw+DqrVnzc5Bvgf4JoioBjnitfRaIXGRN44BtCiNvsZFJUUX/dU4sAJ3uZku
axlnqWzxqB5KEdtmHJzxhi5tWEi55AmutFEPDJ4ZSF8fYBIEg1uNvy+2ltoQ5p0GJnCSVo3erLVX
iRDWqnMUvOSu3xqjOHcKtartt3xXwQCvOC5+vW4=
`pragma protect end_protected
