// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
eNMhMhTTIMpR9HF6+wG+3nXePCqBg8qEwyIKhXfx1TX28nJxNN4qCFnS9zlX9gSN
7EDpdiNxp83L9+8qILQ2FfGoCGgI3eQEqtPdbm97uQjlQ1szYZmxBeR9ONY1KJvK
CK20Y11w+VlIcZgoi4NvMVijp6b4klQjT8/cMmiZImk=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17456)
wQBRHL6UZ72zDcujmS2hcIJCtskDKGsIbmCLTGs1YzctE8oWDoF5OTGFh7dtavDJ
NxUcYaLVv4wDzMaLgN2hcU9KpCZqBzeYQSZgIl1GFgDXRakBgaQ5K9coxb/rzVDi
zGKmPGpYchGS37Egxr2/MpwXOs2NjfFX7r3Kdh1jwFj4Oay2AG6INeOc3+UUzrdS
2KnqaPC4rfjsCLjviCiGroepeHkzng0qHyith3z0NNo9lH9/8R/Y3dAKaBT7Nd8u
g11kjmI9s3HQqw38glB99Sfd2YLGy+L/mlfVE6D6A8enj24aupkyNkhESNIbr2U6
9QyodKnvwE1yI8Qk8thZBRwaCieERLW63yDtck8d/maLY0L4Spmji97Ahy1w7Qkf
8LPATILyUqmgvM/gvr+ogK8h0Hb6YQedlWdqJkM6pd7mTTwECpXaCJoEZuUNEGSk
MnEVSF90AIP+hGmsKv2quzgTqRiUVAaLmY8ftq7c5IPKKnpGCKNQS3Og5rRlvXPX
m+pA57zMVtUZ6FcB7ZeBtCU+Gg9goqm+OmXBHgYvfSOzbKcVGfzFzQswYngJ1XLL
bRjh07GhmwuJs5tHRHgUcSdW0NaN8rUvdyCh5u8JK349yNJ6PGupI3J9xb1neaxJ
rfueIbHGiYnGNYgk8qw6TixpjiNFE6Q2vwg7H3LG+uw+ASoTvdAzav1sGo2hfScf
9ibHixqL2Z7wXMGplG+3VA8SkkfqvT9RsOJsWkmtB5WLbTauZcbyQVSeRxQcgXvo
AyZtk46wEARZcVy+KShBVTT0Goe+ipCEoct++zacZs3BTAheFqMngeaV7VQ7yQsb
mXPix1cWKm2Oyu0YPKFnG/bOWb8xMdkVa2fjkHqrJlE5HTmRLujmCJsqQpKiEL+V
BhKHXKZX9RhBP+VJkfx/iZvu/m8LiH+zO3ZDk6d/be3EnYhNeug+ORiNRXWCSW+s
EejShenXKawteVd56tIkWOOA52gkrtEcEWqrrCJ9LntJx4kD3YAUmy7wgTvN1mmF
znS5+VxMPTCtUNx43+dY2RMm3Ecf4TwhSd2nSkrIcAGwulCgN3lZbkpvW1AD358W
AVa+nl9Vtcp2UPhamLhF3xWi1cjtNdDUxTA5Pvl4e79UD8waP3e5UW1gRb1q2FKL
T5H2rigG6hK84LQ2RGkrZDW5ciQH+yGZIYDSxlEZ9fRKBK76aJ8fb/cccLeEsF6G
COuD6Pw/PTvHJZBAw5SgYjGJ9tKAz++7ceKNb8P+cpp8uGUNkJxkfiJ01wfV7PFS
zOg68QLAnUf0W01eKpV9tkMl/mXGVkaD/I89aL4pVE2G6BtY2oCs8pjg6x27r34T
D1XSzg6PwZOQDTqMqonq38ACffbTe1LJ1xjHR2SBMLoHrhCANH6PK+XFf+VkU+mN
2lAPOUGwA95RR69WsUHId/sVrgYesKiiCbjd/PIv5l9hUuiGV1gaDy0GzWqEIlob
yYvXBCuMYKZ7BTbciDGV/wCLiGthrs3+INJLuexqYgiF3macWxCLwymo52uNu5aH
wDXwe2iFbYUJ4CZGzGfZJwTJRp0CPfXCDq+pkw/USGcVKaCBPHFoUHKmhDHTMWwI
8DhaMB0RSTgBkbEjx2+LbZIb80CMUsEWRH9dki45xLBjN3K1MS/YXChslvSVsxId
lFB6zlfxR4SxiiZscd+xgL9ds6GkQiyHOsUBQqhWTjPOLYOqHcFsVDssEvnLIY09
hOyev64zk/FFUL/efbYZOuznGQYqfVK4UWNgspM1+DlBUo7W2n6Hj3gKGklG3xsN
N1NOZQU7YFt1dXJLvFM4Ypaohw9AqyT7zi05ABoGsUhcTZqGH2w/vIy7OcDC79GT
7v7+QVawP7oPYAyWGsKPVvfTb3nH33/+40LIyFeOUF728q1Ixu3UwxIB0rcliT4j
ypcIW/pOZk53cLla3GmGIpwMfQoTEj8ShsnAn5Jn++5rt49WFXJVnqMNUpAXPvj0
Db7BOpUAfqvRQuxWEJcEh6YHQ7SwVMGbYv4SBtX6uaDww124uvPi5ZF3Q8lLLGq8
SBPjBO0xDoZJJFxBAcdPtb1y6aX2Tra6R2EOaNRon6+LYrzs8Wv/+7Dvph6J6nio
zNvnd36I0GF6Rh6YD6g72P3aOfYZ7Tc2b5yjsRAEYZS6LfIvEn9+MiLs3keUuL3O
QL710YjEf1o4wBzrfpsNI6XMbLwafCIx/xjUw+MuuAt8xBg2HNq6qzB/Ks+lmNDZ
13dV0A39q1pqurmKJ0amnlJDxfx1CYZL9ldKxY5LLVfxk/QQFjC9LL6BK4Ge/7Fm
fUJBQQ4mIHOOeKAfpA7vb6t1INURKD+cM/jP/hsVYLmhKd/TX6itmSfAKu1fhmSH
4Gb3is5OzJEsy+Qdv81Qts1oU3mbZkrRVt91vOk4JsOqOZvT3+vM/qZ7hLYabiyG
oalM1zbg3z7e3jerVTGCYR8Tt1g2W31p/GYJ1W8BvhoUkH9rF+MwFHIe7SKw1Kb1
GZfdsUMDiAMg+qWuoU4u/fBRkCMs2bMQp5bNSV1h63LB2E4eE6lQ0ivT/VvnbgvP
cREIyEbvFSQejfvEs0EwDprZqEkoAo0/t8Hf9c8Q1IRO++fM+mm/0zSAJqqWY0DA
TOcfmeu7Kiz9OK4sRB9koz2AnLG5DHMjTFIizD7SLdoNUP8Zzhh8QaOqSei5GVNT
YhIyWgBVbc2CsDQhdnq9RrGnOvdChpFDaQubvafRlUUMBVtOxAfr2YZnltbPijHS
4rKIPP4PRp07PbJKGlpYXEfaqtFpFuA8BG8JxocgnrmfkuXW0dQ92YddyM2VT2m2
KlbQ46AdShkveXj8BUXVBJhpSqrvwRLXctjfAV+kgVz1fM9wlkp7Vf+0TX4VCfjn
WjShpds11bXRqT3o342iT1YJVx1FrzNSsI0euG5Lde6n82p8rWBOAoScGCYuQj5i
hruLefOUhs+/PlBQiG74p/kT2Np3595SGsOiwVheZg5/geHk507IjklFA/VtYtF9
Xgyq5LAM5DyNbFcCwOFQ1iSH4Dv/Q4iRXnk9cgNQAbnTqS3FoaMhrMPXncA4dwlt
6Rxm7qHxciEobTFvj0N5IoBQtpIdlbunsLXroKO+eljX6Uy5Kj1VWCnbGIx66XBE
Cp9yaSXlMRjJXatfhJ/eiT8FDChlAsVJLPYArQYwN9LbfsQ0EoUpiitytxjOkhYk
vVM2JHDt+s9DTvQFrvvxeYr183c1sO6ijY2Hkh3XZlrQV5CZnLxwC8qqaJxfM4b9
Jp2RaqF4bXuvL9xq4tm3H927V0SAfzAVk8EftIcZ7qimBI2Pn0ENuPylt1YsB6CH
KO7YhUb52UyS6onsRGOsILRndQzCqpUZKJQQKCZ/c966SUhWRMpu/pVprcn1Xj+w
Sj2aLadgMWNjv/iNk6IzuQ/bqXsOrKe9BfCAeegn2w9rdHqp1yMAvJaucsUDpsmr
1JTlDDpZYUAmv5w7DtdGWIEmVgZfpPxcW+sfEUWnkndm2Mf9DTFIkXSRFLDKbP7C
sLgESjpdpEMtMtK7aspvfp1wSEthtx575QF8llcYr1hEjs2I08ZVAkjtCXcp0bKx
quXMHx8PWcuiHRzXvfFrPAgiGUZjH0pTMIJO782jw6fWg7QAMXmMgsphAX6fdzMb
zvZBR/d4p2Ui+CPE5XeCjF/HCi2fBhNEVSAjOF1LreQwzfR9zJYP1x4cCNxbBb8D
E3lQhmJwY52y7bNmyrVYrMaGX3sVCsOFUnpwnda8XoAM8zvqeQrAfxvAketg6Vgy
cER41g7xZyKt6ob/9xE9MZjH3+XQTh5DDR0QS0eJzx2hV59Xtqf50UAxyduhvyDe
ksUYFVPn6k0oaTqKknvIpr/CsLybhB08EvUAiu19w7sZeATX8gLfwzjb5iJ0bfrk
VEmaMUimMew4nehtMJuWv6HphvTAr6lAdKtf8CtNfLO0pW6b7bBSaHW+zjIQqg0F
GKbb2wZLLQ4Hh84QoqWfQrGgulBv7D3o4OPfaEqw+3U2JDEudODFapz+E59iSrXt
mwfFcQyu04vQONMr6uVILYLU6d1zWSJPJ4p3L20XPANz6JsDlosABmQ7D73EDXKu
uBS6hkR67gk0i4w5SsYXqjIKfy6HhxG/m6EnaPoZHHHuPCqXGN3zyxDdN1H8CLsY
lbo1SX3VulmghaB5CsUEuIvhjsdNFcQDCrYYhxvsXS/lhRapc1Of44EiVHDQcQ/I
q7WpFaS7h3ZmMcsHMk2pC9WlXaUGoQ5xOFL8sUMJKMTQuNui8xO3MWuiZzNHIQPA
rOW02lbBlPd/rdmeYjsrTSnFsiSrOlmDyJU8vXBCeDBu2no/iwpvStBRrrfkdPQa
ex1oYGz79wWjdpD0kzjh0IW2iZ1s9MsPNW9UZOLGw0k70ap0SRfq3jTlGubCIdep
YOFcvw3nbdUznp8OmgbH0THOGt8uc5UIVGgTDxQFe+9rwYzGIYb2RqJQ/iMUTZ7s
qijUKnQZ+ZN5CV8ny1Q2UCFjbaw6NcAO+CmXgE5jYP2chp8dqAAAoW99044TB9tn
ll3nJaidcUKc52EYpN5767stABJqF/9+mChmTN2c1LWx53MeHqQKasvHkKR2wwNw
Pj0OtHyFvbuU7aRXCMNyXdUxquLfRQ1V585oVueE/GQ5769MsOu7WpgeXZJMmg4K
jb/aot0Srh58GKWD6pkt953Q8Bzt/m9vmqgC2y3gw+9HeCuYlm67kdh/1+BEM3hG
S9jXMjQrGyMruEKMV2j1wnk5z2qUvwFPSa6VHRVGNFwwf06WL++nXyZk1TfjFcqo
nQ2fZ6DNE3BUBzV/jpdVgu/4117s3K8NLc4Jr4S4JmApMvZU3p9e0hRKhQ1o7GhG
Y8vm4gHbf6EWSE3KF1OwyUZpszESnNkeRewrzSMxtLah7RW+eRnFW4ZCvuGuuNSQ
C05P6FKB/fjyGnO7GTi7ewIXpXm0WBpkuSBZI3xthv1/nPAJGt7K0EOJjJSS0CaU
DzODb+XC0qqK5DAMjL2UkX/c6vTYi+RdaCyOkRVQGB4lfDWTNGBFISzT3T2QTY77
J0+jQ1KEcKyQDs1XggIRxVAdZpsZQnAqqWhmmqxMhyGlRsNapetka3hil7O/qI4C
DXow6gdFUOJruaw1CjvGldEwVMCtZWApiagMlJ51UXKT3Hj2rfRfc5pO2QO5ZarT
+87fC6tK/r8dFyLR8iuSYGyRr/GOtd69oOR8G898o3mDBCfTEJ9Nc4Jyn2oWh5cw
6SL7krgYEUel+t/CW0oKfTiabHeRU4zJWM0ZH3iQDFwl8MlBP2917HgOePTbTQhG
3NJxVhFAKOmIlrijGP6ncrdBoNV4ub7G+3+dfl174zogKX93lGmYfNV7NNBwMz7V
CDfuicnUM0GyluPSbuCoInmbI6TqZdBV8BSbjJBAXoXatKILixCr7PXn51TRRWUz
oZ/D4DAjKfC2Kqno9GdjKRiknjhsnL7P56dVT30b0MeDfiwqbSyUro3CEDKUFARb
uwbVJoQdMqkzRb11b46S+LOme/nb79XyhN2h+dskUtWjUAb8XIyGWqc1HA6KMD89
EVKeNIhWcyCKITe2Ki8hr9R14S6UZ9LeZ7QAil8U+YH3qkjVOhs1gYMYPpBMK9Ur
TBulPDjYfg/j44VNAKgGoDFVrWAQik2/jPRlby/0Jixex5KNs/I7T5AaEHyV8GNw
Tqsab4GvwbhE2swjDQ62MgtwYlr5Z1nnPCxEvalLFIitrqniP5BAOQVfOuq5/E+C
MxcRk3akOUmyc4v0TTgnn6Q3J8JQXiue4ZPkidvQUVVYgr6dMrdjoe9i1SyU/xCU
6jTJnAo9Yenn1gR93oat0qj8OuX5XftUNQGmqbnAtYmx+3VB/y2ot/W6jBgIaWvA
IGwtPkX1Z10wb4Iiemo2I53iD+a4kwY9qCe+JdeITQ00QAbsaJhs9JLejL1J7N1m
1apumohNceTlCSfYYDO+l8PWeqrY/nlXMbqydOgjcAoFOZJrQktRIoRQV7AvfjN/
RrJkVjtrj4fN+5vYApTmWVeGmQvqFPu/TzoOQY8+Eg2kNMyu4f1cFn6Zd14nla6j
F1TC209u70S1gE+6coeRCcYUJbRbiGBYhCszdOm3aloA90//+bgal79VTMYbiYrQ
KT/lmimQYKBbMLcWYWZqjDUzIYAH/v+JQXw4x7nsDfyivcMX6IqLC2jTiTgZVmqa
OZiv95q1Y72o4ZQ3tcG8cBANoGijLNyKtww91NbcpEt7MTzjszppRUgHFg3pFsS/
7p20pt3/8SGJ1/TuJUqXznXLAjtv2dcyxalXAKFHuRF2j0oQBGlwKn/1qlHzNcAG
5iLUMq4gRnRQmOjIxFvIaJ/FUxAJy0MtiCQrakiG4uly1B/b2xYWn1Yi52CvbfTL
afuDgNRlbJ4QBrG36I5gwSrr4Ev1/0xcT7GDYEFS/iKUayvBCKGT5a69XW0PHPqR
aJQ+zykq9A/b7S3/wzMVJegopYp3Y0qQ++OXyxZpCCjGIQEDppzHdZ4EG+s5Krdk
D12cs3KOIXo0gfGaZhKp2JTgUmdlB6ouuLpKKQ1mxtEFFAAP0/LtPgJxJnUXlhNs
F4cOTqfx/GFK26wz2EzWYwyJCIkK673q3F3++gCLuSAtlFAB9um5waw729bsOd5x
ZTwp2y589ODWKzLRG0MUhQlpAX9tnuvWyOKh89oEdAdqVncmfBoep2L/juzlgv/Q
UmIXMv536eAhzmk1ggyBRqba2IaNgWFNtBx7dGpiY0LVMNXWabqzxVjFJqAhpb07
3aPDiRF4OsYCAW0mYXC3o+AigleYe/E3lQvr//8Itz6CWg/PoYFhmXWiH1AB2FVt
FJNSHwPk0ETJ6g/SOMgSLCv0vaXSLg8dW3kZxKjLIv+zXPhdu4akM/CDau8XHCbA
C2oMYwRON8+2H+uilJ7wXJwjV3yr82oG6V5Spdj4Mv0IyLvO+QdMZJImMhbCsSh3
dShYbtQ4TbSVwdfqYqhvKSWUDavqTTVHwBMqTDX+qx7aN2w08ZJzVoBfUaUvfywb
fwunlzc8CfKAsk7Zh2pYidyyBhx2ynsDHjed3KUEOVhSk9Fe1QSkB9LMGa+P0WNr
cXIQBiglqR+QEyEUf2U7nb/O2WomidleuPOOp1Cd3/NNxbGA4K3gbQANGeud2dc7
cTV6YcXSjZ54vqAdPvWuallwRoEsCtpLoiQI7Em20md/cpFSkrq86URBRnlXqJUB
07qTmA2k+mrKy7K4WMwJiX+/aZXQs9P9JP/nABHS1aeElArWircrI5YHWhcEbs7a
KgRjRrhUJIapGX4wyogJObJCiH8ARDeaSorTjE9DxGjoHH2SgwgECKE/sE0mSFqJ
wgGuSTSlzCxIPRkcs8QZg5s5Qd/WsFFazq7s+xchAlE9BwEM8uHgrGcbbZXBzcDu
38FIlTXMAYBkjf4USY67I920KTFBAEs4aLt1lgQvv+aQMm+acSQa8YelCytIHWgf
s0AzRE5OaodRZFRmM0FC2W/bcBE9TKU7kp2nQmsIALPOGvja+P/041BKREGij7Uh
GVE2syRD0Pm+qKUvSCnj/lbFELQgjmatLep6jdc8jH3eujcuL+K/NCTiYiiNLg52
1cstcdb+xkTNpGxxYY5MFiaefIJfbL/JXzIcdjkNt9etUjjR1bzC1ZAIYrxLt7W+
eipYG5ioACmTSWnR24zD8o1ctWJO0q8LllVzTsV0s5nesiwG6M9x3p1EYS7cwuvU
F6qQwdQujKbD5HE8Z4MUOI4eTG9pYsgy+57nGR58/PCDhrWfgw2drbqgkydmDeZm
Qj9ZMB/dZT15xjFxJ1moi76W95GXrNd2OpSwNpy1OzljJv8TX94j+Zv79WdeA13e
KMGtICKaPkBmqskeMpgvo1KTu/DW9b8XzZBh+opw3I6vcNozIW9kybmFdKz+FcvR
v69pZcluFxwSpcAjzPe0SqK8aNSLfbl7nl8pYmZ7Y3nudbwaRNiRhTWaKT0LaYQd
r/4s9rD+a93gjfvlC+/ae0JWDGld6QohCBj7S+ElOhhM2yCpW3Dv1FPIfbk245Kj
etmN2Mgmj0MohZJjfkpzTc0z4XtTMz84oxqmz76np4BwFdTdA23BTeDM7JIbtFRw
8zU/NSpEDfGj/a3lSoxpDdg7A6VI2XhAoh/MpXO+fJX9eQfoCpGzGpQNsJSwZL44
nJAIhsgLayGB0VNF4m9mleog5b7gr8T6Hvm0um21JpmDLShYd9rxzSnXyHUUc5gQ
xFYQG5IknceVeEMNwmiw6v7duMVYEOhZSbZM2ZDKKqQCbUxcJ+sKfyqkq0L+Fkdo
/rBLpMRrmG7vlpwU6qfpyw8WKHgUbjcUq+9GWRGfB9XsbHjFXp586+eUIY++NPBd
yStiyYyUZ5uoKcKcl+JXV656gJO1y0DxFf/eSfCu4lAgbKBztVjrNCLhDNcla+vt
TaGv9fVwJVISqcEPXdFIld0tEML+gvh051YsJyRERIPlT84hdsvYZjGyKrM1Kp62
Jw9scKP8MTx9Gbf0W3sW5+lg6GFp3cOXE5cJFTr+LFqGaTOm/BUrwx8+8dOWidvq
V6jWors374m75pvRJA9NDkOS+lIr3ioYVn55qIuzqEJR4KoQMslWlgOrEuBJNHya
3YQBXiBlabe7kkxZf264ese2Y1R+NlHqkfPkPtae6Y73tfCxI3uAVPoGR0Jw2hog
xELblO9JgeIdaYtt7vGCC7X2a5KXIfyobNN1K8JnrBTDh5CGsjrPTiNknAiGoyOm
tLGliU6Yh/68ulGkfoZyPTLb3YO+Aod28EGwT8Tdz7ZoLT8HpY+8II8lA99bWPC9
6fhJvnpvQdFfGH7ATCrffbJ4BVYPG0VtpXuELve6AKEDY0SvcnuPtdgbGeEDpKp6
8ZsbZh8xOo1VN/t6RnTAVmTnPwjkiyWc6pM9uty48GjXL4JMnACqu0XMpF/L16Ud
2tfykizgTcjnOVrSIyWNpJOGYXFWn8LMNNiikGD1dhNfTncPQgGQkH6M0iaX5UYv
oJrlVeemLrx3iKlDit06XVjTSoA6hJh0TJFS6+2pgYOUQQVf9ATmrCO1t60WYOcI
bJtuAgkx3UumaQoAMYBcxYGfEQr0yu1cwVIl3PWnh/3qUZIiBFmhIJaxsnAd0gX0
UxquA4GGWwyT7i5eUqII52aPlt+oQfusicHz25mKUnDfeyk8DPHVya4+qYTBRFKd
dl79uN//1IjVuiY3FNm7O+lF+MR9VUAHc1qlcA5ILnEYUbNsCuIWGaS/JqmnRDrU
0tB3os+yCDnWfy/xWQWjvAID+pwkYmhhlYWOOY14H+5EsIDXGzgHdw93r6x7JZuf
V6pyGZ99TTFqLX9G08l1yBu5dTlYz14PNFu6hCDfBLAcQIJQNAczNJv9YCgdp81y
1Fxv2CrAiNjHfpTrHqF33pUvs/Kd+sCjPYnhKaev+7bDK2oBW+MK2ftwJGdKhiiR
0O9EOq2AquTlFIckW5VzwdL9L2XQ6uUCphVn8d4NiL0mE5VJH92ZGp4MGv/Ojurm
qcqZwhWdANQ6o4Z854TwUnK7VWIzEybfJmtCh9LMjpo3nsiz6dwSyTCdNkInguWq
BCk1/rz8bBijusuIgPPD6GNea3Jeqblt+iRZYw0kJGF6BKBho0BMO9w2/wfsvXGd
lxNtxf01emLV2O4kGrKY8ncgk8uWLQ/osXTC+LvCmw2mtWe71/wmakWGV7+2QxZq
WT5zWFB9g6vbnn7/52xx1g/dz2tmvjR87Y7iJ7ukyalprHDXWm53PHym75QF7oD5
WlH5JyNlDlVM0QJntcTkjBx5RKBjAiSNKH0vGoO7L8+mA/4dLTEBF0ME85B+X/z3
ZpzYrlixLuwGpMI4xMBX6RBf8dHpndzQRFPSqTwDT93NFUlgM+F2yJpxLxIfgHgZ
JWgfQk4B6Ed+p5TOQQw6h6HRGlWyDzRMJESXPg+kpeY0ewbkhDBfBZqm3mx2TZPb
+pNAZTcsVBA3USbtw72qqo3F0LtCO//VTJ8WqX6PXT/BwkOEyavE+UoseP0Wx3R0
HdkCWRjSRfqck84ZIbLC/tsUw1hHN8sQ4xXHwqsjooEO4iAzgqPeB+gQOLJO/RCm
BxaFfoZ8DtnQu/0+RtuFcl4K5JNaA3Tsb1Z0timXtFK0hv2VyH53qmBE+1hudttW
pAqVZungjwkPXeBlrwH2f49QKPItlUgsmXZjH6PjchbgvavSUO9tj/yGJn3y9V/Q
FsiXW9GQN9OGPBbKdt1SNhhwlKE4MyEkn3nMg4YZs/pGFuNHQUdLCzA6PoIbd1iA
QWRDggM309/f6i0FckykCCukM9UetdzzNlSEeVwXSjGqEjx1ZirUM3R6CesLU+09
oUIAQgz8D6SCif4AK/otAMzZtNFE1oC3KsuWkrTZ+EP/IYLAcKuLRv9C4t0HX7w+
T/aI35PNHBQpA3IlgGWhRIHBTuZaOrvCWCnh43FsogsgvhDorMPRhSHacsOZBB0T
tKG+L7DEzBLGUP6WitBMDBaH/veCqFt9peDxaVytIAM4oywTQW+blXgiuH5DxwMm
SA4soOhq70P2yEAu4t4yVuaJSFCfSOYsz+aPdwkK9CZ2KnGbPQD4wzQKfxSb07vB
g2LkAn7+SymKVJh7Q41uU+Q+qUXtSRL2Da7cjNTYFZzLSEk9CahpkWVT8QHkY7L+
u/SBfOTF7O/KOL+ygf5R6CknUBVFasVDAOxWWxHMMPuvR5fBsnjcEYPTQzfO45tN
TyxD3UGGDA46ZxQK1Bm2/ektIXzUkT4UPnABgQec19iThhuCq7Qy5Z7GQEq94wi8
hsPa8nKXmj+rDYaKLIPMGKmsAe3w7McKtb9TMYucXluHBHdR7fhZO11F3BoE+GB7
kSQLKwluu3NlXxSH4QpaX6D/ZmI1jJEw0QKUIbk+T7a8RVR+RJqGheToxYet4kpq
yzD6Gh9befQGxXLpRjU26NVh4epV/Uw+onGYhdwHS9Y3FDjjHqX81yZxjTk4F6HX
AqZuDUSjW8xYsZjjcH0Z7syJvh2EzpsURRr8+lrJMb5/2b3qPM8MDHmB9kzrfRW7
d+ZnOj/e6fnHvISX8yfyIQj4imaaouUYMNFaBUVplZu4PHrv7JJBa8WnyfCUdM51
7D29tMUZXa9mVZolTWQHalbshdyKfYI60C+hP2DYgX2KXrXE0WtgEIXmUU1koe9f
6E+FZSjlNkSJQV+VXGmRUyJdCvgOKhu/qaL87IWleR6YcP4nByvouzD8dLcjULnX
qnDniq8kCTFsRhnfUY5Gzkz52Mq1cHbdX4UaNbdi7qaHZX+ULTFP1b2sSdbARcm9
n/9k7DiOiyE+lkhzGKtfAZ/j6ah61Z3Is41RHhDF8Vf37Isk6jo4mnqLiXPt+aD8
5v8pZB3SwNdogOnLBThyOn3b4iUmkBaqioLcZqo14cs4d+NjKyqKOl1OKkyU5d8i
d7scvgL4q6PSPdw9Uwj+EVaqY+x//HDeJL5J1Likrc/xOp1fKOer+boXWQts90Wr
xFK0AuzU2VaI7PvNgxJimWv0dqYVzsnDgT5QXMJ17MEUKolhYjkX555/wm3qoDad
wa4yMAOGjK9VwDOW1xpR5K4jNAKmlJl6hQ5VyivQG4sQUndnGKRMY0gui1Es7TE4
MMCKpXwr+/Z4ifakRBruiBa12Ag5uCs1kgtWPZmtM97NpRcRb9xfs9E9iUOE3lEL
X5CMrtWPUKOiXEXbAvqEx1HS+ebEbiZFDk6NitlPK7EfuBbElEa4JXwN6noox1KO
e3Ql0DljkbkE0FtnqbNRZsZ+oLGaqnK4ze5uFIK202yq5aW8XWzfSC6hN8sxxO4Y
sJ+IobRkBOXWVgSjym9FPOyaJY/1YvPgDGnsJB0dRK8046RoMG2vyCkZcisCGXI4
4LwEhGs+pxw7X7RIVogf1H7Ptt5vrxNt7+fNwWegU8SVrMtzljomZQ53GjQ0p7Zb
ZdOU6LtJntkyWTs9y+wgId3DDhidS5GL+SEVMQw0DiP+9G6dyhAymvhECzTLyXy7
6ATC47i3s0/qq59QJ0XB3q6czxo0vkM1eifbLMgh5MAcX+6fA8+5TEu7QpNVfjTK
Mr9ldfBc6biA5oe2FmiVUd++Wv3aGDlekqhoaAyXUTChmvSKCeojzYLn3J/QreAO
JWTaR1KYWFjzKwOupaS+Uonn1YBTpEkITwmWExJ5/+aKVMJYmiPr+wKlILYrZkpH
IF6lQ+RmI0JkGp0V4cMkYZkyKVKIPrGBG2X5VNvBf3Gwj5qMPQWhXxr84oKmNWbC
bD/XtmCiX86Efs5kJXYR2DxFnl8T8X97T9PaMNCuzyyuWr8xIzAg+U2r8l2Bfawv
NnNDB5ZoZGPfIOqm48mu7oz5uApO7q/PTOLspiMoFpr5am2nmk33z1kd6Pnfl1V5
L0J/C5SgK1MKY8e2m92p4JIpBQjaZ4tMXGLG5C3pHbXYkUdxAwsNdXF1TcsGPTy5
GTrXC5S+n3Xa/jR9sLwWF6Q1kcRiTueLpsZJrDmyFjRKjzu9i0dXvG05tsh5DDRJ
D4B9NRxQsToWMZG8OgNvTCcQMQJQyCmF4uJ1Z0V5y2WLZoi2Ecv9mKFG+evqToIi
x1VQfGVhghGktLKKIIMSGGBPEAprXirzIG/VIcbTs45lIkj8akA/hBcH/SR5TFV1
oq08L8cdrO0HbxkqiIlhwmXkEejLFS/OzPyrsFeRuse1F27WuHOfjOt6I8CKjWeE
vBu8pngXBtWsDpy3eKRZlJaRS3UqnSPO1qUsNWDi1EwpseDcfBuRdL0hJqlM4lir
i7pcIMQ26YYS4osLNs6Qi1NU/KdiFzA1LDSgIT9wAyebOmddSIVqqFN2sVcdCXJQ
gUCuDTHW/WJiWSssDcf0EDiMm6ZtwPNdWmcnQJfQ2oUlrqgp+eSAvBQkYOWbx+fX
N12Iqm5RQmCTsJ8Ae2vnJdIZ+TlRCmCTa6MLCh9NJwXPrgEuzLvCyLVzt40iX8wV
DJlytIXCsELCCcQ2tv2koUAfkbQlssYtdRImJPYc4AVE5Oiv06yw9D7ydZ/UjjxT
MQrfBKeG5npWRfRAy25IafLiPLaPJjRS9AleOGdu7+VUbl3uX8zlFVTUj58T31Bo
Itb6DlVBFqLZ3LFxXLHtpzf6h/MMTE6UelXFdSJ7oEP1OJn8T2q5z+N2g33ZlvOz
pbEHK0zSDFje7tXur0waW4Fam4SOdETqRmBE/PEBBsiXd8kbz80sk+W9DOoev3xt
48Ds/gYG4tyf13+IMZBAKViXsvULvg6CPnFOkC4bKaxozP6Ts/DT+u/sq34gch8b
D89xZxhIIeex8QeWkgKF2tCFyVeAXVmi8zcv0EAvclrQoARA6pOuNoWKG+54jx2E
G6cMHBktnMRZI12XkJ50vvVJfiv1BCnpodlbro8gjZKqAF2aB/fFqob9IBiVqnSn
OXRDfiKSEF8Vcw66iLd4CgtXjDfPlG95XskdjOZwCTUILB1EYKfsXvXkWz8giwDQ
NiVmjig1eLoq9++o7f0ak9EDn7K/HXQqZ3mEqmtTUGnwdAe53/w+ke8J0XItgJbD
mQL0mCU1s9xWZwmtg20uv1y37NV+ilVMtZ3NuFCNWBVUcK0bamdWZwSj+80PS3HD
OUBnEbHie59/9TUTZ3DIWxIv3QCpLp4Vldxl3Z+vmBWTJCXHdrrgpcKMELU9ydRD
DUDu8oBzyQH1ANwRjCWKVye2AZp2bVBox41vqp0H2Boopww+Sdmgd421Kpsf3KR/
1tEH5umzpktw6fXoJmsCbLdE0Yvfr/8t+gXHeM3s3bGJoctVgGAZgyqKGhCbu60V
1mqPfR0o0dYc1FVVSv4xKd76QFq92Y5nl4vhDeWCyaSDa+rzDZNxmB5alZnm8W3q
WS84zMWLjG+yXIBg6a6zhPQO7ygmaU+fjREw1xu53Xac0exMr7zvy4RBZ0k11AzJ
ozt+6aFPS3H+AmlDoEELPIRszvT31qslFYtejQ1NLcR3j6aiO88dOfJAiffYCxu2
Gj4pjVTjCpdPYzz8rjTwvw8JPcWcSyXhEb/v7hntbzhdlTM5sslLiBKZ734H6M3u
LNnW5AvdGxMUlFfRoT/NxvXxAz3eJOuNmnkn2fxy6W8m2aOD3jLj7Jm+QucoMYf6
U6mFZ2YnvyptsMf/p2TwjQJKMUV37iYp4rJJu9XDm0zKwnSuWbflb9NM2nI6CB7F
HlE1NYbdt0DLJFR1t/H7T3THGMkQf7DfSDVWtqpoKDvE8O8ylzXR1wqnU6/aLshb
DFnGaHb8bk5mc6zXJDqTpxTUvOf4W1vMhgJdDqlPFug1Ojewk14MGqB7gtOcPkvH
58lxJHL69E5yOT4Ug9/WMPhnxZn/99K3Iw18Md5lIoYKtfjweytY8CkNdN4loRkb
FBVJeuvOzERyK/0eAJ2ZhLlhlXHpUDGshB8V0I+J+NxeV1DejMLomqDvA/X//ahe
I7kK+XCdvsEmD9+KQU9jzLfLsVAnk0XN9/8Y9d+K6QVT+WbDzL0rQhZJWKotX4Yh
gYU+20rqVRW2F4Nur5GqOlZl1YdZyijhXNW8O2MdGpUdXl6tzN0Tqnk1YXahOpv8
eudNq9Jr7+fICDX6MtnXVAtJcndx+rEnlAXe1PyfnuahtKcPIFzoHGeaePdMBqzq
uBRtE+ylmkasmXZzCtOTxaoXfAwYAxwE5MSlNftIiCODD4gQ09rGr4tPUE/smUMq
ltZ/S3Bb29Oae1ctjH0NXYbgX04NNOBQUQYuWQp7QmZ/qzCDyfZiv8MRhw/vAxbQ
6x52CMOQbTCWUKmMSrRLyCc6r9kYZ6eF0W93aPxFX03JJgIJEWYYNvBcte5WQLTt
1JAESO1bsnfADymSPLXHBO4OELJsXSATo+JvTVFI2jXbMoG9fmByax8NawO6Ya79
7a2xY2BuTUoulySnV74maObSJl6mqZf/J2i+oSUZZXXjvpLi6r05eIjvoHvgeHz5
Rh/VE/T+2zUjWFxNmTkV1oq+7tfkU+us1MXbeNMvueQliODTHIgBqLTyunfeoUCQ
SUanLMW9yOioIvV8ZUo+QElSDtYUxxWvHW9d50Gu9UnUNFar6uGNelTECV3EI/w6
f10E7YnJSUwd3jG88+0eEEwqoxaa/35VaES1H9LAuKf9O/mhtRo1BpSP/0LVA5UR
5FKfbxor72hCyr/MVKwpL8waO1USnz7RFO29IW2nx9zh7MIvDqpPQ3TNOzqIEBCe
jGRuTbDDJQPsa0suH38ZGWk60h4Dpaol0yHJolZAsYSCJdt17880933I2tqgpd3D
1r9KeEMtcxDciKznDulodjAqKFJEGLBiVvXFFqDtarJvraIdr/qJH1bnbByNveBB
CAaJBQODl0QIbpdhm9p+sVbqypU3Hnd3DwsBph5kKtXf+rn6kZKrQziZbahYVXL1
fD2DhVRb45LgIBtlUdsT5TKaw6KaRI0akRY9191wEy+I3meArtP38vQRHXU62RqX
zzDuKvGk6EhSq5FX3Q6R5kboOMFTAHmjBzDmOl+JVRW8F3xsW1VBXWEKY/AyHG3k
Ppe57+OExhp0iy0iXhJpx1Q+CDHzV3dMnfbMX2ITVro2vYjXjzEevWX9k2S5TTPH
pKXBJwE5b02ZJI4z0WV3ofNCtRhHBEmDtNfBN9NJqyWuZbnS4y1x8FcB4T16zht3
W/NQhYDaBDN6tqxdj9qxOs+l4kIzdObUQfN82xYGcKtk6Zq8lrCXwx1u3UiEyIzz
SbDcGZFBXUV+e1nl6+JbYQ41xsKisNpSDdEZxAc2xYKdQ07wj0v/+0q09Uib35xK
qx50A204mfCnpwsH4MdFqwtyXPSgdykJs8jm9XDbZw3iY1RCMH9GJamR3MLG/lhO
iH8chDjTKdh5f9xbfwmjR/zox86uZWtwdQJ0897a2N057WI7JnTdYtj2lSVfHdTJ
neWpMJmYKStatX9MV02XYjaY5iq9nVikwHBzKiHo0l4O+PXVQRrFGNTO1BuQTD/p
7nBMI4zI7mZ6VBI7MmktcVk/ln+MrcF9FHRpeZNc/16xsYBxhmLmeoaraa2u9VF/
Brxuo77KOv/It7QSDOtdV6c0JQGWuy2xvciWc3LGItFq+lRaY+coU1JtezcGg14i
261kENxXlGoUKXFyHOAoUAQhSZsn4NA3fRa0FpnY34TKDTB4nE4ebi9ms84vBLX8
j+MkoPoTIBxXbKWBzTtWEgjhb7ef05XCZTLpkllx5pLauxXaajmMOxgjdWqJ76Us
jWaMg19cjEqckOkPHh2vqHaU3yJHQJ5NAPgM6e+6eHCj9H+1AlSCSRMed0bVSEvf
lSMM3xQBYLX5uUse0UbXuu4qzT9FOrRCN58vnyAEB3Gv5Hvcq9p3RFxzUkHfwnVg
8bhUHEkvpk+EvsS39kfXvZmdKd0gyqhSHG7hJRPISVn4/HB8hU0DlegWL4+FdCBC
Oh+zcb60OgA1YBePyofOWOrBTZ7VOf1cPF7yIsMi9KI13nCyNLwTImJAYlmu7K0U
566XRF13l1gnhL2Bz3Ma0hqyDfkvX23nP2/2JSNwoGb0gUZEFY590zJkmGsTWEO0
QMyU9o5xSCxqputm0lQHg2viqYjV/GUZVA4EFusiK/a4BBYlu5QvfQQYsRG6B1Wd
sQuECvYPtOimaMifJfk6Zu42OlqkPMHtd72eD3T1X1yHSi1hfqrfQYluxARr9ERy
d8OaACiKWdI9YOck8iEQcBxw8J9HFS9IqFixFNz7O4wBeRfygvHU6EgoDxYWmQdX
4/CzJaf5o9Sb5BoTSZAgn88YrOJMuo9E2FGYfI/G7LiOCCbx9viz3EcaFRWPjm5B
ZG3JNf+NE/1AFlPaM7jTALLhRwsXYFfD1XCCvbsANFYmLcmBQXcsmi9sELJOgopE
YJrnkzo2p7b0/QhkKrm56v3dEmI+ab9c4v2meywZlPWk1PQkU2TeYmfJgkh0zzrC
S0yOH30jC/a/CCImXtRmQx8AWuXYwq5nbAg8CwkmyuRgeXUgW4Ng+5ViHFRIZXeI
mcQIN58GThBDdXcQo5A8n7K9FnI03YG6tPnuxXZREGVLwKjiSU0ncKNtFOEK2KOf
m48CgG255uxHq2B7FWT8ORsO8z2bB0beImtsASt1n+4DlhDYIV47UepkQOimUNCF
AIhElmuKvHSG6Qzk3CVyVFMCrvLzMt49r2iscZPh7SC+53JCW3qqQecDi8u9IBpB
yykE6dltjX+j+RyP4TyObkDxNGq1W1rxxg2vhMwcByxh1nEPP+CS6ijHMVfBOXvK
xjSk7q/vjnIsxERlX2wLNeCgH1AsgYIACDKTCIa8SF5ePmu2L4Xc3gmOwAZRRdfM
pCi6WM+WWM43OW7X++kJsK8ks4jQgId5mgvG/qxsxMAx31fPjHg5tfxVTNY7YImc
/83ZDixJDIPQsf5rVzeyANv8fwNQ6p4v2tOgexC9KieC0YPFQEfJTuDDa3EhjdYy
VGwcOmdIBb3HNLFGK3+GiToU7D6BKULb9gUIeT31ZG/tx77OORXIGfA2QHEA/KOm
XnIj26hljx1S4iu7SmTBk2ZTk/tP2nu1cokIItAJXWyGUZVAkf4k1vNVQG6X6yXV
aRTLGvyeTbj1bukOnnr3oI+w0CnjbYRr+D3ApS8LslFbxxnNfo5KgMFVPsN7PHyk
ocsYYO2vwiEoJW7SnvZjPYG8gVTpw8Xu+vtXM/qBT964ig7fvRl3kpF0rAWeX1vH
gMLTGTITGJ27Wo1PoqeSjv/YUuJyKMR4CoqIwHFdWVbL0AsPc6uTwt2s0Pogdop5
43y3YiWVLmUrtKbgkfuz3YYePFEe+EhV+AmUH6R8lJ8sYMebOlKxpf/Cz3NCTbIr
Z+qk1E0/qcDqQBvjrOd3XY1mVS+ZJ37QiFoaBfGyS66v5LtFFyFRaWTKkVV9PU2b
RlbfaXoL7Huq/SNXOGeWixZDMHRd9sgQ2Z8mRDUlofoa6PJB7QZgzzDiXasn59AI
Ud35/P1UuCVNGWfrxzb5l6W/aJg7ejGxC5Iz+kY8jYne/jZfKDt9b4G0C5EZCUDm
iYQw2eRWl6TYaBa6PwAcLmXpee/8cW29bG7xrXra3RU0mJ2XjzESkaKJ+5bz2UUF
DtOjVpsE1HtuRFlaGWuGvL6eNYhwNt1NhANkUU4MVP6xg6RqyDEZ8T1zsl38VKPR
UmjR2wGwpzm9aiveMrYlURIhx2pwwg/M/be/9qnbjdfTiJpGHrz5IhJ5WMXTcor9
I6wpH27kZMcnDLvNQwgbs7dt3I/3MH00hN1GPTj20cp/GPUYCCU37nbcGu85E6PP
lEnoFnjkK4N2BCsO8fNBkxmyeFtnbcpj3LQMtvM9Z2+p8A1v3ZE3j4LomG/O26kp
xCb0JVvzvgUk3LmOcx2Ag2bRA6iL3z8UJq6MmsAbD2OPRLzEjH5eILiFR8QNgcy9
F8CZdYGlxVvONYCkHkh7D7dVVXdVM9kLmUjRQ0S4wcV3uPLRUMJhlZrUX3Edsakn
dfVKbXOXTKlev9vhj0ofOCU2aJ3i7olFyK+AzibNuMBUAmdVHAEkGPgmtYBGPBc/
FsVobWtuugbIRv0pRi4bzJt009Mo+/a/wvkQtqq7qkoP0HejGc9TBBSmsVvqrHzb
E8axEHro3rziHZf4JnPC2LxWD7ZLegqSQyXLJaDMZcQBpNKL0SxhI2XMguanonU9
jz/S+lMpqSt28QuPLmKeNwy8shWCdjFvKcR1NERBVp1OicI+Sj9xDYQZz+EClOtH
Id73QKWkp0V4qwzVklfQwHv7D80NP9P85J3AwpJEApHlnWo1bLDfGEfilG+P+HSS
KFNuD+R9sW+NSJOAL08Z/JuLEEU34kfMsI5ADRH9KEG/zdlrE6anAj8iFBfydJEA
n9IGj7uDoaXI0M62tc5LBBkyvfpTw1IGR7FYVA0HCBDR7y7LsMeMOj3iGPQc77dS
yy7Ca+utJ8U5JJsXFuYK+rcW/S93ofkd0XZXnYUfy9YtmogbQn0dA61J+v+n09Hg
32gqZa6UZjZWm9fw8Rcl7tFyyXsBeVL4UJ8XjbwKdoJWeLm+oj0rCF6u7nz1d4i4
fIUjavxrY6wneB32MZPR1g1GLQw1KPfqhOU1eCmlVNvhrJVwEMuJo3Hge8adTDx/
lwMlHXxYM6xhSKfZwuIumdrXxK26HtXE5YTwoO09Rx2P4+yBjj6rJPP26eD8ZRF9
iURBj/HcSjnz+ivTrrxFuk9bb5y17fra5VHIpST6mhhBxg7j9Z3lnZbf/eR71TC1
5l/8SzCABGM2Dp4hS+8q7ifvhxsppEihRYhEBJYeaFWOTf7gTzCp4smHQ6XOqrpX
ptXAOPSSGy+A+jiCg2WeH0C3XC7tTNu9ftnSNCFcSRvN5hxubURzv8ypBOPWgNAB
DEgE8dcIuqXJAnHhUQzW0U65gc+98M+s+09zC1tlFlxIflSbIoGQVOPgTOGVWMFL
ytN272APZBYGiypUPj9Cxb/KEeS0fl8XEd4bszWfpFOG2VLfdS/4sY4iUcUkzeOr
1fcRbVDh7AYT57/9WM5JSVdrk3rrVefsijs6bU63XVazLsGmyZukod4OOjlBXL91
DA6Z5fHjbcHtVSlAusvhctXPUzdYMUVmBj3sgqvJRQ4Stu5uXhIrMOX5uptXXTdB
CIzJXdtGdfJT+uYcyKnNRSDulPMhqOYgwTWVkrCEpLH9zQLvwCuigjh6LepaXkgf
mHCJxgO4m+uwnmIM3emaD8Sv/PJ5NISbqKcN7kp94tUfZiaGi+WgsuDaqUAjRerz
Qq76AkK89JAFNhuOAGix68eKrF6/noF7Hu/HjZiPQbTxDiSV8Eih4QMLEzKX1p2U
B2Ng5Y94cycycqE9IvDwQIgBT5klfTYVkftJ07SlvFI4lwrIPUZl6vCe/yxiVSfD
QPy5ge/qUIYdJwGN5IGM7WUOyPq4DYnF7jY7JVjt2SfOxgFCACTgKYm+dfv2kPaC
DlOf3lezkU1NU7YU7GlhJ+v90g7wUwrA5NYDvDo11fUePtSGghzhJrmhGQfaGMFz
ma9j2FBDxcDkdIQ+f4Y8PAzg076rHhX7yht1yk9n+aGZ6hb2Vk4d/GWEm/LNxDR6
KowujDPeDQ1BdfzroSmsBBUaJjuUMco6Xbm4xC0c0yCG5jlSOAqMC6ZIlD/2a14U
6CH2pwhgdYFv78ULi90k/b/znO3M74bSppnQVvti5Li8xzVt63k5k+POAH7+jRrO
pwNvRu3g+msLxDXvgxNQYd6hzB2daTPcAoMAF6nuIhuRSapHH7Obze9PyAb8b9ul
3JaW026uuUIVD7EAM5kvYr87uLjIfzl60sF/90sR7v5DN8im3zCZhsujIBzDnMy0
QuPDr2Tk47lwHViXt9S8U+p69kcKengf3CGx8ounjU0VfDwgy7Tm6krvhLAtld9B
4LzFWZ88t48sqUFdwzK/OJkE/Mgf6Jocq50y795v2WV3HgUtdt8ggka3Y3j95kLZ
v4atLFtBpMDSFBsYaGhGnoUjuBQGUeUTi4ezCrFprXvz+/E3Lvto8Y0Jgy1iIK30
yaOo7FXHEAWxr6b5cdkF3cXstRLksZwrPyWxEkvxxDAXx5GkEla/LjcqkPB+5cxk
MMzWCRE9N7qnoBCeRJNx5/PpmqaDsbqkdK29g9O9nOZ6uTQ2BWfo1shgrVMIMcpG
tZFVRClI3ZP+Q0HkVCJuZfiUvK30lOnJkp+Tr9lSERPs6R4anmr54YRiyCMDCXQx
1wNlUECTiDPq7d+KR42F81R9DBT/NIGoMpoZyCdE7vABqJPZb+3ETfCLvi3ewh3K
A2yDg3ZaHRvXfW4jkS3ZKQDsYIjgoTcRN17QxEMpZYxqwRm+IN67AdP+l07FRJf/
TZUn1g4jKPI+FV56VUNkv6uyvQunD2oMjDoODeyMumww8v/w0DAAMR6BQzn3VONx
Wza5VosOjY99wMi2+dU+u2hf8Y/iQOoP07mqHoIK2WBzxYL811dpS7+R8H6uOnJn
4Uflt1k2FpOgPLwSo0cbf94tx2UAgAHFGHAuSB+B/pX5+M4LQA9OuX7JrjpCPHXi
W3ZM810pktR7KnldxbCCf0qtKBdhOXL9mvv83d5OqVpLFowHLd8XCqqOy7gWc5o+
mBrVmjA1IFotYVS5f5IFCLXncpXhW8V1Q7g1S2Jvb8Z2hiPBkuyPDic051JCXwes
FWJz1PWHhT6/G78z4UULmSxsaFuHq87bUJ5Ygkbn9k90ASMAp9MnfVZKZ3ub5/ol
ZYsTmC4ieJKR+1AH8LbWjR9GyXdEdst2Hzrjph8/8/wJtM3tHdD6zHtCo1oc3svj
rs0nxufaQJVqsHuBTRegDwYmEl7u7lXAKsSrQq8xETluneH7jexuy/fIT5gglP/v
GNCWtqliMlq+TznAEJ4aiJDI8s2U1p1tJJkCNPLhcZIuth9evtVz95Bd18LZUt4o
MxBTCICe1dKQFL4rQhqS8pVwwHEpjFc/FLV4OemsDgNf7FlrsuyyHvvWO8iBslxK
P20vF3Ttkcwn6m7v9ZT7+y+y9B0FX2jEkakSUuJ85vlWiAk1f3LHcLWtpOBYHsAc
BHamKPWCh8WOf3AQv/fEYXPt8aX1sKS+1ONBVFy3pSf3UrSpAbMI61HNzMrlfYu3
dpwwuCbSdavEM5vAMw9KkOj64XMIvw2q6/nVUW56Kzxj6LaqcV5dAxMrx2BC+FoW
YnaIO3JxhgiVHUqAFNKYLSwgkoTLQSZVas79JDlRaIw+SD6aVGG1kPCjSCObyjXI
0WkOuJfxtAFrZE416cWK7U0RuPAbKZ4Xh91W/7k5VlgoDT1GREHKdtdP6afxTV0F
nNIH1Z+d6Uwyj+n6DIrSAeaA0Zese33biG/9C/0w9HOOsyqu0Awhdn7cM9pd6RAh
43KoYtufLP61//nm6bRxBABIfYifZNk2hluU7eye3HcXrY7T+owAcoBmkrjYTpj4
b8MWzPAc/hAZnrzrtYEmlMGWkq8HuIzJ17HL0XXdUn/g6f6EdG+xRsZDNVTyYIzY
LPpmPfv8XcxP/eTe+debYFXpfSq9HoB3miP4KpLUL25ozYSfFFRBrf30Z0TQWIVa
+S3vPzo01PV6uIIXcpQigaKk2q6DjGoGieQgRWbheXtbehfMygp5ebdHk8s9wiUq
+52Rd/22qmtHcNsYFQPdKhuK2M5twcfmcGvsKcwf7mdpwTBEediAh/koW2Kf6nw5
EMBL7CAe/52pYK45No3vh3dr6DGROEuNlCzb1uFOKGzWJ/4KKJmWexSM3nab8m4m
7YEHVdoPFd18AR/FUoWM6bqO/UnrsdD2/VH9cLB5UrjtdWmugJEE1qt9r6QQfZLn
vzuw8/SH+D3iPPDRnIvT023oUCcD3PlwSkl4979oGr9u+UAVyvSfM/eUAL/HsCQ9
2i3WuiwluKNZZcIvuLWxgHm9tQPy78TDtVJrrrwI+F8RbL3FxVQU0JBzmnxYuv9S
COHUH4cCzgwEVWUXlHDP9KtRLwCyxpB7vx49WBws4hk2+a5qHeIT1DvVTrz+QHKL
HUJ9Dnw7cLrk4JJiR48dJIKxXSH3mIu/KRXYiM5Zea8LsuNsXFbObTwe6p6RidJD
zYe7syLhOLioGaVMTRGDBLwR4NPUyek939oU+7ISSDvDsTVOrk9Pp3b2HobtqRLE
PvAize2we014ebgOk8JjbIgbyC4U6YZecl9T4ofcvbuJLW3DVqRrkfTWuYfdKHSB
//i4loH665tlKkuyomR17Zv6GssHTSTusZYwIr1dKb11z66x4KCbv9lmw/gMQ/3e
Cg29SdvEAvPpwKwsmQLtnhEzACUrLjqU4rwreS3w+Ps6h7ojZGn52NFy4aXUestQ
LSR3iWb/JE/+snyNlWTYVTtEktzNxzDKMOw6VfWox2eu36o1jnclSEMx5OzxRMCa
7C2rcjo65torVmX+XxjSEg4zAR1UpzEs0R57k31X1BzLJzx5nwG00jwhmTu6tlAq
m12SFR6EooPtKNbW/H0Jr/5BkMMX0ym5m8wTktsC57ZhjqrBQSGS4qqJxfdqP7hd
wWa1A9pBKp8eeJaGssaEYsjyiDZV0gD2BrHhfiH7WQNcKYNZOQBHRMx7sXUGnVOq
lu94nhXT57FceWAqisrCDD7lcee2DjbqgEQMOOLq4f9D+Y8Ne4Un2sZ7rgvXJUFb
L+vdmaLBUp+DA9LCJeEy5Wj7wyen77gplEfnTBgM06tBnwolgR8wtY86CY0Zgbmg
o1hIMpSwdfjWbG89dEfs005XfZFl2SOB8neTPuzFNVI=
`pragma protect end_protected
