
module ALTCLK (
	inclk,
	outclk);	

	input		inclk;
	output		outclk;
endmodule
