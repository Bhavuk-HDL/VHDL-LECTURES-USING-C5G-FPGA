// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:43:28 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
Ck0bdgxHpvJgKX+hEUBsV5T1wtD/fVLPTwy54yqCx5YyC6K1NQQ9qFI0ilFz8D6z
w/kiKXRQ8LpobPY28blUejxkPbdrVKAzIEJn3CTklRe4ksYFB8akeNEZcqgTzdWp
NgFr5OibAxR2O91OhmuGBGy+ecubszG+WHNieEyVJpg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 30112)
Ueyk7rDPMrQdQgaMwdN/eBC+P8a30c0sGd3ELfjvik+V5Zj/Dv2kKpC7oRBc0pGS
nTlY2pOGqLCxXCov/VZDSkgNS/2lTfdY3GGPWowAreDgAQ+qLm7jupwj1GVA/5rg
NIdPURH8HQk2H5LAx1TmzO023I7lH+8KUh0LBhEKXaI3N4HIi614znc85VmQuwGN
Y+TO0skbuZwHC2pAGhA/1uQp9nRAclCdmDsS8apYNTHnMOgFn1Eyn4LfDszT1sno
p9SNKqNO5bol0+xncG49JFeKANTp7ZtLh14YOiCuvnKrOTTvT+rsZxighEwHxs2K
NRMiMl2tVtp70HhNTa+jbAEknjvH+JvIb6bUphLLU9jDx9qPegk5Ns1U2wmgdqIT
9iz35yW5Al67D4hwBgbUqPXLQWo7rY5EGa3GG87fHr480xtI0o3dpLzhnEsfZDnW
GELwbBDdNlUyTpGxaOdJOqCnRzPeIwwYmjYTgWt0oQYzMzR8BcIunnJ+8mjQ91VC
SlibQ3Oz6PK1lp4B+RMtWdqK1dADp043Zq6Ig/qzb8DnpnoObSVHs8syWsgOO30m
o3R0Biw7aX9IQ1BqvX0AoDdTF0fHgF/VRmPWz++t9UHfhFlU8M5xzxnRSydJDsJm
xCCTJQdCm8oVmQJstU/TSBA6/dP0/n0r4hxTCKOzyNjD/LyVrlVj22Sjm891qPMN
KK0suOAl2JIIbD0ae66BqlqMbtyQoL1ri1Hhb1uEisMM/J/+RIJq1l9orig7wZAA
p8kZ4ZeX2tNwwlXnRXdLPK7wFp7BZVwlkjD6B5rpUcbgIhVpUaGS1+EHHYvmzcDF
zqz/FjalMOd97I7Q/GYblYuWBjhiw2JDgfToR8dSXjaGxLdg12ZWp7LGdy2HGkNx
ShJqPcwDUm3RE6256bxTVzbFzTNjpy6pOHO25r99/pqQ4tP0SS+gQ7mAZcmNty9D
EjUUjfmyRJ7jssh55M6VxNq07jFdMDeOxBhjAW7Frjsjp1Tl6vXEf8icWyh+V5X5
OCdj5pXrtTmQR/wl+Q0xyNDm0g2kBlrPY2OO5uJEjlpQcGWPSSOmNlHb2p24Bimm
qDzm8jq8n0Jt4GOxfZYfH9jlYeult5Nsxt06sTG7MLfbLLwSEYgT8Pmnh+nv5jMU
7WwwIGYEkai8ts8yIHd7HA5E6ED86PWyTNp0je7SKUDfIF/HecPoEzD/Ijprrmkm
HxgdUxilyDYSoN7vjblHaRV4zalgzMrqjPZNJA2LGeRJJIH/MMiht2JaOdbSk5BK
6AnpFO0Xr7lLApPmfQmRxIg34oZNRh0TgBHVg4xEJ75wGvG3fY3SL8wFm7mt0FXk
3eO5nr2oaKIta05WyHQ3EZfcww+eeZYsw3NP4Jmutx/nulRqHAWI+Xsa9H4fHiCC
oGhMapqysIt+iRAWzv45c+kGXhBRZf9Yd3NZdn2jSvWbxlAc0AGi+YmtvrSukhuq
wEZX7L7z9OzTXRCr67sjBLAj1/pwzhJk/Sashkpjz9AYCKgMG4adwvQ1CI6ckqZb
kzQOKUTNE+veDaZ/4EpBlkMYmHGSWWIBMkfJThbAxhuYSSTs9v4KL4Ef2+sNW2cv
kCj6lK90TOM3bux7Ta62/k6TUriqmsB4t/Gie40AFpACc5/jy1pmG/vGhhCFwzVV
RXoSCM8dU4TmkQLCkBBCwmwzH5i3snZFJaoCmKPkAf5DV3BSfPlz4z0OFeXH8muk
ZC1lzbL9ePIQE5S8aU5EWExTcCI7iykr7rtEc7EbeKDzeegPUn1YfbEGXYU8RCBu
b1EAJZYIIllnVOXjsqNcRFb0Ae3mPB6UpQcV6cMOQ+jpomEUiurQyun0Sq0Dai0+
gDE/oYWCwViyVLp4wf/SHy8r9nCsNDYQWB+ArDoc7bw8zJ06G0Rxy2Z6DjBOQnZj
Ei/Xoej2jS2mOlr3HQJG5UHX5/oqDJ7dbAWX7gO07G1T6jR3ZIvq6LTxsa4FkK3j
V6Q8snaF8UudopLC0Rgwx8o2qp+yuaA6qq8niYbTLcOOCEy7/xfnW28D96Yh/EBN
eZsZQv5sxcnHSM66VbcI7Ip5uQCN19hqF1h/h4ST+SJ3UHa/Y+Rws6bjY2ZFk9DX
cTOeg33mGhd1rq1zPtulIDJhmNzHOAB8O3yADL5p9xhuYWqVhYycBe27bfpsi2TU
Yady3BsxdLOztylg5uSOfRK2YF3ivWT5FCNWbMznYMsQ98IO43N14ur0bKkoRw+h
UB/SpYxgSs4YB8tUdbDZAxdMUPRZ68yKwrypHQ1CO3DV9q4YyGcoYT4pXVDKQXpr
khcc3sUEAh5EsM4Qf1fbP6vrcK3NIDd64lKfveFNgufhgvIsd50fLaz5DUtqh31Q
4cbU4wvyoyBI3GUk2aVKtlg9WckADjwiULH8mNukZsZ6V+LY27VK6us+9JrVnzL+
u5DAWHB/g3ceRKCoZSpjVuWFAk0kSoM5U26ewrCBTrRkmErvWeJIMAEPu+C5F1s6
TKOz+qFme8xynck+OsEMQ9Bv/g6NPaniQoZ6PSdgIs3YBO7R4zUOPVJgoKaZhI81
fhjIrnwYbRdqr6dkEKio06fVQpu8yK8t5YYd4Fl6jNYqXatDzY0BdgHzXb0D3CkR
j/x8HnJbMW8My7IXB34l14RFNY4gtKoV5en1KtoGiI3ogzUDBCWvSkvQWNsm6m1h
N+4ptZyiDcV2+Bsuq36awwGAvZZiN5kT+FwkFTymUxEVlboj2+IjmbBdnRu6R8JX
ZJmyv4VuuqBE0klBBhWiW7dXtDcIs6iVhMq7Fd5dQwlX53+n+cfWiQ5unE1Y5Y8J
kHtkrDuX+BQoiBAYS1EbadtUYVxwhI4igVD5jbsWF6ALkQBM+dpKhEDhw3xRcl9V
gOlaleCyMJFoaI507x8MEpio32wTeJ5VCI+xl42bzUBCJ3w/xio6+3N6taJ0PsOo
pulE9hcwbDpXDkYJZLYvanRDzgH4aSPp6pUuBZiC3Zup6EcqTFB+UaJ7q1bTHvos
6RZDiEBjmrZLnIi/JoiCGqMZCvX2wx/7cQVtpiXpNYarmLX5Sx7fyOJhk7T46d6e
/AB+W2zOWV5SEZ6oebSa9SX9gF9wXCZFYRW/wrWVdDUXNQ5LzunUx2wNhes8tTqJ
06wNbS6drwe93XSTGGUKrXvoufZLQJjlVCRwGa+4FNLVblkqTbob8IXjKTsx+32T
BhZcqIKN9BDzgy2rj4HkilHpbxpMpe5P1nwuaCGgTHuEXVFOP/vpe25dWKn9iq5b
KI9VzElmKH0VbIPz2c4T5vHDlPFip0szyAUu1HjHsBv70QxWFcxxVDeeeQTaCLls
i+t35uBlzly4Uhc8ZIj1WNOiB5CmGhandRORCKQYxn4KmxpAYWim+tymYLcmx/PH
CnXHGgLl0ztOgIdXTdGlDADWH+7dGHRph/qRHLRJOSMvlnxWQmuPkLzS3uwJZ4hH
SFl5Kwn2FNj5n2N5ix9WcWOpbxcNhypnvL6NSH+cVsL+nJVMJraDEoHM0RiJzL1f
MOBaxDZh7LKd/LYOUuqFM8MlXb0A0IWCDlhtawEtGC33+VOxybjx34Yoq9OSCne1
vpmEqwcUoHTTOaMKp8viAlaS4X4wxFyzUlKpvywmEQgf5ipC7mkEqaGUw+h/+cys
fWrh0gZ+FJb04OOIE39SUcmVmb3ow+KVbQG9De3KlS8JdycertMDpoBrwhFt6WsN
vvVvbsX6jQppEnSt1FxNzQjcRXdjltoPMVYx2M5qw6Fyw0oQ/JE7d8ahBjGAKprY
xrMZwUrOLTn57SGhi2CnC4Cu6R4Kk3xqGgEiN9klt4Rf4M5jp+MnnaPr2fewn5MY
jcXd2qwTexsUDgSxTAL3krz/l/U3OTJVllSs3qkA5GCaeeQAcLc3Cdu6hXJb4Uq7
HSR3eQSR1ypKkx37cchss3k0vmeynpZiItfVoolfnLyjfUPhHTxMDxoc/bnXqvov
bcsMIty/NENMDAfgAqQ06gUFeAl0YyVU0QxbuZVjofRCCs44H6TCbESHDPIelvOj
LDUujKv37pT+eUvAWvkVFeLDChzIXSBKHBHMFhGiTLEIiJDB2ZzCzscO+t47tXzY
w9Zd7/Ch9xQRDtrp88w03AsRxOUbgQLX8LDIm9cmD/f6837qyaf0zAjbCuuXafGZ
t8BH0CpKO+Mr5F07IAzsIVWNWH7ls1tZb+04n05Qdfb2td8dJuz32gjFv0NdG4ds
6zMUKQ9uMPckCxr2pWsfbSyX0wsE5783QiXkqjoVOb+NWnIIcXY0FoQrN2BkMoa9
htp0bheAlgLWE1rPoki1fRYBoptFGyA4Q44gO06JiTjfKO+Io3J9TdHdrlE3KnlB
kgPYYOoL4ytowm/6MClfSDl+4XrwKvSHPxO0vsxBrw7twHgq9ovkVIoBlHegzHoY
dz45/vycSzFzR9yEBHaLylhKqzlHvI3h4+QXBMF6+Ccsaklw7uDN41+0Js1C+DHf
u1VFx/u6dW+mAiVRFgVxeeJEAVZ7L5F6U0SSXPrGpiCguFNQ1TmKMe7R8CklfJgc
8Y8ntKTBZ2EUHwFLcFgqD/Y+yahsq2PrVxZ0NzEDFSf7/sVCm/7jpk4cYGQar6fN
GVDrhRZkRw86SCtRPZuXFDH91K2OQex8XUlFbER8nc2siuJpi5BkNbkcccZuCWI+
0dqzMKHV2GYDG6smufE50N2U6UWJLr9eHiBLVgrmKoqyfaw1Cuym1Zx2h3hI3CMT
NwE5qFciBgGJn/mXpl0DjVnqqu2DBKetVUUAAupgUiYl6lcsj7EpY4y9kUfL95bk
mROxoBqgHVrLsR4wRKQf+sg8whkCDFTihh8aEpEPYXMfyYBcoTuUlgFsYv/kmfth
/lTz9pt9CCI23GpVnnExW3lH1RFJwN+V0OxPkNW8+0wWfwOcJKOhsebNDTcbLxwW
+9XmKQ1SxmzNJQO4d1nirbrritD9be4nls8BkmoSxe1ISVA54hiZY8Dbxa+pNG/9
e/szzWp3A46Zl8gt7atmQ7ogEE08Te4wt7QqzM1woZhnuLupGDUzwpJBKlwhW2Wg
CcA+CNUjUrl6VNnd/BLE3SDfGLJoJcDMlbKTDm3FX6pM3zwqTmYhDPIR+b0AeHi/
SevROIJnRL6tzJsQSQB6MMAYfarRcFtgEzlVfn40UdxZOplvi4SoOnxrtIN8vLsn
9nFYf2O+xGFBhCwhwRltLOXsUQrPmiKtKspayUMkf1WSCH51SHzpgYJyevSsp0K4
V142kuyBgKu/b0+GqKF87eIZoru7b0ptHTmMyQa/EYIxlrtu0qhSDNvjZ+AHfSxk
w2B32tmnF6ncwJMZVog4MHGezDWuyR1YE95vi83xIe4dHjCkSkjAtdrnwybETNu6
1BTRLu5/NsKzMj2lzOKlLkXf/w0itkek0Pj9OELPtRoqmJl3/nk/b25J07yHCVeq
cQMxEchlPYE04/WbAVObi5nxBRwxt1IrWwIGE3CTTiA7lPiN8CL31wgoeGpuioht
FBlzZ4P2wQYXrleT06k8A8MyKgbDErTxMU/w92flbC2NuAsS3xRenhZfMDndJhuR
kF8ROqjjSRkZNPlb3hz9XBpUj+SDzUWOrjqBmk31zgJ8V+L3pdtdN+hA0JaujJHk
QdxgxJx4iAJX/yspIWaL+FZ3uCs8mUisAe0VwIjj8VpM+efpfQ0l6jZwRxIUT3mF
4AoRezQt4Gal5iCsqxlon0VvFw58LwkXKllawzdCdUj59s3cagP/bp8EHj5Jsyul
OH6g+Z/QtNvzLr+pYTplOv3SBbd2tah0K8q+3ZIaALspAPpx/5k9GG5fC+LJRZqu
gyVV5fnUW+LA+2UpCP2PaKHYJEEK7Uf3zQSOpi3xS+K5ulWMcz3yGVKWMcJiO1SE
nCThFIWb0V6As2y2m3Z7EqfxnM1o/LyBJNfni0LRES1eLonGPl0DHMhURYpejJO8
TLkKJQUxyxf3+xF4f2G6Mk9x/MnAJQZBXof6vY3QQNc1nkNegfrpr7IbrOHEU5Qr
clxuOmwXgrT2SAMWrMj854qJ4NtwHWMbsmlaaSnMiRfCS45hpFOMHuvfjMsyoslh
NkzGiqR7WfxwmAPcgfPbcArrOk5z/7eWNjR4rfNzdUW2MjkU+AD6s6x5bePFDVeG
dAXbdoTiNcSXUpBID46RZp6fkLb0mePwNxxGe+SSpvTdoSvJXIxS1fDwTJ3y7jPP
6dJOtAor6/NVnUS9Vju3xRot9Gas2hqlOgvGcm45MOFtwJN3EuNoyldz09OthEC6
fq8+g5aOdk3/tkbc0FqDI+yHV0r1f/YXtVciNaGfMcQoIfSs3T+/C7i/+UIjeDtC
oDTFcmv7zuIafWbMlybHRsSuKtxsPjmn6U/axRszy/Zq9j6r57qkMNmWSzvS+71a
kgJczNBQQSgJ3YujiX9SboJLSyx7SOwruloZT2++oZIcQvxRZE1s982DFuQSqkP/
XGTKTMa+UcZAJI9F+5ew8DJYkp5MEgsh4MMN41VxeIdOceJ61c1xaMT8RqsTgCc/
7Rr55QBOah5F54FPK3b1RFLyu69xB9KJj4/ELxK8FQdlNaDAI+723ULmAub9E9Jx
0d2MitCeB38jwB4EDcQYbA+jK6VSBNB2tlT0qaCdrqScfstMxV+ftQLIx80rVKZW
gilAbRxdI0Qn9jBqdrpT6eQ6DPhgY5OFRL+GezMBXwgTUyddpnF1ojLs1wk3Ywn8
1zYL5xHMp9f2dt15hn9DkcSAn0Mmka0X/o3z0sDVatG5TYkKZOKwolUQp5sBe+En
zSFY5+QLC0mOgPC51LWPsJO47KuV2NLfrv/BUpLL/BApj15dHK7hCfODmYiINcxS
fqyAjvaTCFvV1/wG5yf6DJRKUsyWhXfhcVfIUUvyDzL4zqvz4/eOBI8Amk8ZJFMW
RuyjGPpUEddW5BVeVddQ4vTLpemqmJi+UIGgDLQUYfdxT5iBGVoPAmXGsMtDVS45
suwGKgckNgrQ91FYNqsvk0WBQY1s/e1piCruVZDQ7letrvOdhvN/ajCvM+ih0xHC
Za7taEXYilcq7i0n2EraLWdgdrI0QfREhVh0s+2EdlbAg/1IM7zx/TnG2x9I2/83
NHoXkf8JpVTBs2bdkNpLuxRQy6k+q5mVihYsoNOhGsP7lCiR/UxedWRibkmawEdC
kKGZC5pxc7XB0sEQTVw1aV9WRTdXb9grj/fKHTqnyBa1gP/4QAlsallbc2oUauOq
fYsj0GBtuidQ0/cz9gNpko+LPS6PaRCCJ7fC+8LbNFYLQTvKZnrZKANc8tfqEWFP
51sTgE7FFOJ14MUwn02miRA4WZ07LNnJbnRj4in+G1zEeZYpafIYwGZxkHK2MzoX
58KIVzkNiL3cg49IYNKeDp4JWUazJIY0J3Q0OJPo5SnET22f8sX/1h7crJDqDQh+
N06d5OVe9wAHWaSCEkHkYIkGuGgIXIsG3erYhaQYpzCNs0WhFNxzfrY4HH9veKge
wnsVrBEUpg24pgM6RwX0cTj9M/XeDDUaYCyd2z1UPuZ3W5I67STLhLSLh17TlH3S
z+UiXLGFSq+qjE+G10NJZrA9qYYPAdbBWgLg2/1SlCEauyc2LnYaS57F0RW2lw5l
0vsZZR9zCH51nAmu+g9yc94fTsOwVsDlibOvqCgDQkG0C8dcdGlDhN/z5l28ci63
sdKxr+4mJ6d2MmMeYiZF0LNkDyK8z3tLTNyhrThtmQrbk89fx0k2MsUDwC7bDNZL
ifdh76QTcT5hau6jnwtmdIaJcKi3JOH6LmRjzvD6wWXlYI9NCdJYF07uZ7jP1d+S
SXEXoI+dtUx6Q6zul9Zfa5bWLlMx7KExGJ641SJYZk7fCzGATs5IIipN0Evj82OA
575vOzLb+wJAb6TcDMqUYoVyWpJB6dKZBL6zBRlXcx31EM5+IvNVgC9UoAevTOpB
WEykKfplIk5x/7xm6B6zUtPfnZsCjQ//saxeLagCR5BY7ZlJAsyQDT3MmpoHh3lh
zOMKTiLB/2ViAe6dl0xkXXMTLEQm/IRJj9jMK6Dd546YKCyJ0u4IWidRdo4MhcIQ
bPtDeXeh037wcaCDj3FQuseyP52bbtK3qdOVws85n9slsQWb2d5XnLVNQDKhNynL
wS08x+eQ6UHiy2uHW+bHzMvE2N2T+5hqHgd1Ol6/5fK7q7na5pylZRUQaDT/var+
kA1LFNoSWuMXDHHcrkFlm6JXt3/NI2JucEGltLYrURlN7EpSF/WGM9cy0t6FVUPR
nDbcWUrnDCchqkQSy4xgEZ45bWiVQRfyqvGVrESDMXUvyNlWi3r1RoqNZp+uclBg
n/lVUmjulEghOPYAANc5LLTrTzdogOGrxQ9TJ833czFRfnaYp3mSqkJ4rF5Wcf0H
2VjzJ3tU0/1HDE6QY9Iwyw/imyE3hc0rO8r45ys+k5UuJbG6iPNJKCCJ1UQXY8QX
Ukcb1NC7D5zog5spXA/LpZ6VBrxGiiPFUKXqf8OfRuwVOasBwg8kPBvHg8+hRSjr
3AdMqGxgHRY9P+qqHbcmz/QeDOGM8NdQ6dfpEarwdmqBhWQzMMgmVz0psaSnWJBl
fPrhsIuzo39Au5rVMNjv6HWUZOHBLjyCPhQaRrkaptouUKc7gsLh/fds7o1LL3fq
Vgcj14i0fWVYkgZditSZsEKXz9HHKqUz9GnbLMnk0iePw+ivheYTb0uOpVQfghSA
fdhtunr6Cmq44edPGR/HISL76cGZoV7XTSn2sHx/nOIEH+3mVtpyL8UknKA9LW7d
uQ8ILPOUP+8zeUBmTIQtpHo6Glniv1j6UNLyw+g+k17DWwVeMtTjg+4ghwLMpKXZ
vwYrNyFi3/f6ziwUkILbZAQNN1K7js/FQshha2gf6oxrWbiHMOkxLf/R1rVUp0yt
jSdwvCEOA5nmWstM2J9nZf43TtKQ0IC/AVjFEHtI2BNmX/obIWfmOdk3ztWUOoSj
gkI7E0SLDa7u0YPjUxdyqr2dzinH3QcjCiB+ZIpVNf1HitSfH2jJCEPoRFon83Z7
MqVuU6pP9HO2IpaTmES2+b1dtONU3DSObkpGTuuVsu5g/3NE/oGIZ65dRY0udr7J
lVflY8TFRpQBuVXQgVD+m0BukXOQMIfx+enZ81ditVCk9AB6EHbMKZUMXgoZpzFb
u6JiR1uq8WfSNd+I7F+gywTJtTVXhVOEoB/WAG94TNbEtmnOVStqJjT6nFM1Wieq
UYptuMIx/rxTKOM/g7tm6eQOK532nPcgDfyPrqPXuH0BJSM7oJR5PQBPlLG6eGQ4
sbm24F//OsLZdqFYPRfh1nn4LqFdGfUdgBHaRbSS9OhiEvV3Ej14irAplMTIu5Vg
eh82SBguvxGKBfKuj2W6DJCCJGttAzjUK1F+7y95DuIuYKDywjdoBM2s8Kt2OoLZ
WRuobJGvdp5lGf5zOxJVIFHfs9UrzpwIq0wYec99bbw+RsCo/UpLXcec99z4jfem
kI/Ul9kQcR6w4z6MHJ3O8NOBiOInzecotgeaC2igOHQgnzsUXq4Q6RJkwYVm5Z0y
nJlOSeh/qZfmjsyGFlbJjI4VMOH6qvp1cXbV2ytHpFkYLVw/KvZ1oldxbjutNDnm
Uq0bfO/cUTeF8Kwsco+VKiOvqUtllGgiJEUcUkzJqx1JSOu0tolonxEdjZltQSMd
c9l2eWdtJ1j3TOOE8AiRlyGVMJ1h9o/VRlXdymX0Dccemjp5vEpZUuwkYFP1IvQm
5usDy2ysPCFrJnsZMpgJ0hefCpnhkVqx2f52yNFGx+bGzRdSXuCc2rA27tzpjKbJ
ntjcR9ZNsGfqi1ffqR9Ro5b9r43zJkQJWeuHybF341OonUtguvYEteKoDr8xFUQN
ZwewdfRy1uwhvpTNrLFBmyvJGXUuVX/k7fLDDYvKPjW5xFLC4vlHafbVpMV8Voat
+R5bLAKB3hblItxy7dz0EdViLcXocKAdfp8RLET+BX/ADdQk90y+X/jSlRxZocOI
0Bpni4vXgsdfGE2F2xu/iGEEvitPP5zhSaB8PB8prVOb64YRB3IEyKuAvmfVqG20
qCm59FFx/Bhb3etZBr63KPtz2+u/b3QbaoDsjJDhS0g21/dew4ynGNw1f+Hyl6wY
vSHnmIU4RcqyqMp3ZfI8v5iKBlDWUAXii0uScDZV0So0jPMzsieQaqbVhd5PlSZ8
wLxnJGvVnqUxYWhMz/zP6mULeCksxbdMnmlKUuJ8ad4EtFSed3nAqIe1N3LQH30T
lH8+/HyPfIRiY24aHtJOQzijm2bIZykNNDj8Ly3yg0Kcul5cjgT7edgBdDvy67tw
9D0zTpF4cVf9UWmn/LKlanDHHMxZTFZHy9yJG4rtGyAM6Mz52vRlVrkHD48FmoQ5
5Qk4rp9E++tyskI7M4Cnjm7V4eOfMkgcF9mvqqC8O4hLctoGgrqKIQaUBN9fVJqs
0fQcrUDsqam2ODBt+eC/YQDBsMk9iTT1tQJJTsOIohZB/QePhw2L1k33rZzemB8O
samIup/nsQzp8JpNmJYMwchht0Uu+CekgipNX965gd/9GUzUa8OCD5khZzAnLW3z
8DoPwWUxqBuZR83L3+uMT1jThFUYa9qdts2h7UW4U68QspKwnIbNp2G82mv486kQ
L+9KzkiBEKrjRhrV5QGQVIcR/84hG08P7Vpw7IHIhSxT8qB2NTDAwPJYsrc7arGo
hfWmUV8NpA+fiw4Gyloi3Nj2PBFkFki6fCUty7UUii69zg4XKSasGRp1cisfD3EX
XS1uQ/UgAQP1H8zO/4ab3+5TepUz35AD6yryNrGLggu82tMxasqXC2WnZCFID0Aw
cFUv0JpCmYCPfMx+4JA5yLBxcVYKFaf/6QYLAn1EQ6xq4Q2oKu/G6P7sWieEIPy1
Dds1Qr3YZwL57Yq9/WHnDbqxJIkINXgRiT3jX58jsGnPxpn7/V0dPr1CuMqfZpmb
5C72uokyfrysYyma6rbALqL2+nFphDoIVPMYf8bEYNa/FPm0qBAxcpNc/fOazNIX
yPysw8SiZs0c/Zsby1OL2MheFdRl2UdJ+p5rg3Q//ssKMS+WUMgV2lnbXdC3Pn0n
ytNKkCwK4CwLEi7VBe63XBylQonXPeqsxp5EJDvU4lC9vsPz09juaZXYxs9aVGMt
FTaW9aUtPl/HWR5jWBZEjEofJGHZJPvwZnVhwLyWw18XEd4HZWk2EM/wgcLIsyPC
c8Qnu0R4KMTMxyJsNFcOOhHNF7Y8ZaphJhYH80MDkoebIn/c0MnYqhkFnWzjx0eH
oPhIoRpXo5Yk5kGDS/UKOYGNTxwFSQkkDH2yy4DI7OQepWWct3iOw56dg8b35vop
MHRoXuSffCR20FFuh8jsWih1orrLcrtrX7ui1PYU12wT8OPY4Lm+UkautLeSdx9D
IYckn65Z+5zEoAT+bMw3N1xMtkYN3S67974s3hm/Ty1MhOxt+lnfKO4UOpti9s0g
R3Pp9LF7gCc88yffePul1maRkJHyikJTvKSacRAekjZlyFLOYWun8HrJccbV3GmY
+Rmkvczx0iVDzdUZYm/ItxQjhywQqFwYjxrU1Ntbc+0bWIIwYA0198BEkbJESIhp
+IY10yFcSucB7TihGi3Cgi9X7MBuZCqrneLF4HN3piZd5MEMg2gZ189AEfa01p1G
7pGE/PsKWDBB8+KsRpEtlpudjlucGwG04XMK4Ohcb9FAhsFk6rrE09PSQL2tNDMh
M5p+0/fdE3NlP7xjOVOxE/IgU/sQ8ykaJwvx53jjkIUImRiu8ZCbxpw1fISS1L8u
CZk5sxyUwFhN50owhl9nb4OP+z03u9OMo+fM8LeardonRcRmYxjQ2cgXl5e67AKQ
8D4OP7gSeCjF12HgutZHJa0AuOrQpZQdoFGBI65Ze9lgzdmTWbnFrsuaBtU6f/y8
LXUDUk6ga9rffTyIGLFogfeqoYR/jzAM3D9R72DogAseVd/f1+9249Xdkx6MAB/T
TIXXXV/H759qvT7Xd7LcanyA7s8VVSKP/J2zuZ5deNj2nFj6lXB3uB0FIXw+ryFg
NWLGkVpFqf3kyyuCckZ3TIYNsJrbB0bXOEfrt0u2VdW8/1IA+2cJ0i9zDMedjKG6
xTyDdkEdqJDnHvEIDCxezZYnOYDj+qBe3fLtHruzWCGfQ/O4J4pMNunG2qKxc/ZC
IxrzBo2rhvc0Ybq5qLiBATRS8yRT9dlh0l0Uby2yO0hELgeDxp5VvMbLcTfL4Bx9
D1bcg28IKanSwOnaWaenT+K3gURrBt9Hr3RrUNgKIoTdxmrG/83aE4gX3qc3t8OJ
JM5t1H19tAtyiN1qqNfDDfBrnlbPsvY9OWLTLeFV5gx6QJ/fgfZ+FiJ2mmSQdZH1
A6hXJNNqAspPPmNKVkmqrkHoWkEjMbysGosHTpZBA7POm9sb5PBGWju5R+fxO8aH
2/uyGluEL3/iHfO6TvSUbBCnEQbhuy/OuN4S91yqj53BgJzY+qhE5YbaS9u1spJA
3hx42t0fOynuBhQNAg1BIpspy0t8LuFy6W+spOnAF5GNB9eYOaX8d/2WppSNLN3T
X+RL47wZHowlMvAFCgKJ13crMb/NJRYBhgS4mYxCxzp9UJ+QNIWMVcb5XMd+QwBR
7JSeFQiVTSXdX076McOIRVIGdEjvAq2bRhJ524t95ED68ob09Hh/6DBNIdlidSgD
NuhA1pAK8SFExfSqZ48cAmjF8zAffM16I7xJH1lKdaRedHGMjVbjbW8K4ubcga+s
VNcvBwYUlkERwGITUhvcXUZ/RfR8OjrIXX2ADVAUt0mosKJWzNC781iAppoLCrjP
RdnZuztAMzXKS1QGy4Nlk4FwgbjvxrVYRw+xGPS0kuP4bDqpDGuEG0VpGnjbf61y
2DOzpbeYd0zY6+HGukUxEaImDnHAjLt/ABr7YZde9sDABhK99Gyp24wZRnYWyg6l
tdPqcS50uVjmX77MNgRzjogjj6PauAIPcVaI/xItd+mGXuDCpdX56ZfrlwzLHiAW
5EygJpDBzmSI7CDm/3u6nw02GAxSBC+fHI2/7TjFbkeQFYWECqybAyvjq3xP4+LC
Fr92JNETfudq/aiscw/sMaqTA/oc6ATzH+IyfK+MsUejgJ0fu87Bz97Nl64/rEUf
FvGojVCNH98vRqz40SIlEbQV/6SCtKDHtK+7OZz0/Mz3EyYZA+q1Z13qivelgsoC
S2aP/UE0xTIymMl5NTPo2CKMvQamMxyY/O19s6po79Lf+Gmtkg88u8yAALqfbAKt
ZhH+Lfg8ijksldgK9paix7CJbPprmZn3Ez98drWRrLQ261QC2/PyU+cEiS+8lchl
G4CYhY3qs2A+Qy85iAxp2a/iqANJQTl7HXTWp3gCsvDrB230FoT9PRQtpyCnVlpf
HgWLOYTzEYVNXPV0wGUAcdwpT7gt21YGHAmL9j+S4RPb0hiUNFkmgLm80b4Ft0ph
LB03P8FiZF/VSnwQUOE6nfXHEQ6Edg4QPL2pMIVUSFYHeiS1F/Z/xl2YDtZf1xp0
CaAV+6Mq+2I1GWLzQoytRdYPWb8fcucynjYJ3zKOgZec9aHl+cV4EiGxJVVfK5Tz
f5t5iwfianTs+zSF/Et8mybBoKMbphQpNovXotIWnxzFkz90Uoac2Mso5MBF2RNC
VamseoXmd1ZzKmRbC1Z+gqXsCA8ZJCQ+709WMmoE9Q+oKCBcEOjV2qhefQUCF7rO
dd+QY3h1CzuOwMZOK8PACtfPG+SDkSFzzkekuFGYh8SPrQd8ZaoPfO3F0ncvZGyK
yym3OvrAUcHe8StXJpdhy14L7wHBWZ6EC7LJswAil7cfESXH5E2CICY3yD5GvvuB
azBOz1g/F21vtKZEAiOpilAshm/np7mOJvkUWEaB6CPnD/dyGPVbJlbJxFY+H6lI
C2q+PGl05ZlHRabjBB45ZG6swnXUrfqDwWOZqqTvEdRIpPlyJt7xlA66HeE263Oy
dWKbx/qvfD5t4VWUbwIVPO7cQMjNldKa+Mvu4qIq/CK+XttdVW7+OTzRu/m1njPr
Al84/qXQB9z1L2aZ+EzAjqdkHCKTNcVFX2sCkxD7MQPxPF4DqXha2rNs3UNI4NgA
vddnTddyfMMFXgZWv/KwQ4CkwkMeK8UtJU+se3z1ndDVxwHOMsenI16ig2IpwSGh
ubhziQI6l7FK+ocRPX3RRbtCO7G/X7Qwd1X5PRd0APXZ61+eV+ui+s9hfEWbJ1jN
beCjMc5vOk4qWsChdWdmMaHr8FvdPa+/Mu92ZATuxztiXRscZG6eO3oH6zR3ShSJ
q/6f4ClgMtTcaREjz9YwH6VuNWzG06gddyLLZ/HSQYQKc1FBKAL8hBprY38qxOmM
EsHmxjFJc9Gwg3nP6P4WC/ssTKASh/qcBTZTG8oD5TFGNHI/KhN0WY4Xh82yullE
QqPAtrq6bwXKoVp/LxKuG6aXGjPGia2iskj0xx7xdg1xCx65gOsQJSovZg/q4ni6
PrmbnoQnnz0jtqh8lgt8kuvly/KTl03eL4QW7k1ScgB2bpl5io+5a89HafItGNle
Xs5N4fYQVF36on5f4yXNFacWtt67rrJgP8RJvHDy5HYnkUnS+aeCYiseSd7cjsQ/
LrwxDjMZzZaPkFoWK9QeFpm95hy6Ior118SxM0qIvfwX8E13FVNDqLRhYR2V8HXl
zOtXlBwEr/oQX9S2CwWx36A+jXlBY0ighzjcMpUWgkNZoMByKCXSkk6R0YEfyCmQ
UBt3XeuwAGUPFFCkGtae+X8krepEPBXX326AaKstje3j6qiGv8ZIgXo0+0mJ/GEV
WpdQOxD5HDDejVKoa0wKUiEZd2mDGArh/FsBBbPLCBMqU8ccidGC07yWtnlqs93h
aPlpDXzWV+VsgsQHx9GNmG6SaimlNqHEvxs7sJORN74KXeetphIlApW/G3ZpQ+7I
ZjWWoxB00DweELf0AsTp2SKHb1pnHopDkephGXjiHxRijeGbTqJTV4/b9kgJIasx
iRwn0aqm5E+GUTmCE6L89z40jFwckvOKe6M3Iar93h+bEh8hm9a8UVQMiD/c9+kM
75JclMJVGdiB8ZJ+efVjimDNz66SCHS/etu/qipONXeZME6/95qnTyjENt/KLQmj
flY0qYOnT42DVpXcUoo0Ui58r6z9xTAa8slneUTE4mZIae6+shL0cf88qHo9hKLc
TnBvp5tF3vdyzDChEQdn7nmcy0bthzeYHIOhvt/ZJDO4DKZNDdYTswdc5xO0l8oh
+5uwOnjM9SJftbVj+YueurmgHB3JMABCV6vI7vvWb4RgO5utb3Gt2YAvsicQy7ju
iuiVymaamgwrul6V77hu+Q3+R3rYeIjAwrI3R1U4bc79/bYPyCWG72KfV1lQgtSN
5lu2x9XKiKTwgFt9PVV/i8YtB+KG0f3OXe3ALvHKak1i9F6vhuv6X/ypZyTHajyL
JAgP4KolvU1N8acg+NxVd+ylZITwpjoHjHI2A90lfRJ2Ga4w1rxbd9QEtAuRVHUM
r5ZTDwNECf3lvQ0q7mmyVvZZ892grh9k1GXW764l7xMtNfRYEqtBuxQjPhvk/N0y
VizuEXVDCDrZk1KWOtBLioR4FtM9Z/0ZsmIivmph3oVLQnBVKIf2R4x9JoP4pCS3
J24LYtb8h0hyICn55cmImtOU6uDfEGHn2Gh3w2kgMl/wDTfSalh7DbEu332JYQUW
D38UVdW4owUMmQF9UkXH1k7XJ7ZnazNqbWP9oVtwun8dsxBe3tY8/SqVBBhXVws6
y3d9ev4WzxjbrLdcR5GkY6khVwvU+wr/R4lnkqrbsS9LaUhtkrHs2QEdHbLpM+Ia
ixaGLNHCCX/R5LTmIOAV7aP/rQvWZjRsMjSu7A4T5eC6/kb0R4BZhhwq+92zePG5
h5pA+uPmd8PiZfNa9Ag8WtGOtUSCSTl+DTTR+aIJo5YssTpM7HO3u+eLWjUUupF9
c2UjJ0vUf132gPn5ZTdicofP1NrO+4CHOclRWnGlHQ64OMp8DZ9x0Amez4ruJ0Yw
IWRAVZ1vKScgF2W755lKEZ7GOlkdxywwsJFYKb6FoAIBANea1qniKhyt8+Qlj8OY
NrGRSWZdTUb5s034ROj3+Epv8HOmM+VMEKY9zPlrCl2Deb28pvY3jOiGk5M+10sE
/MSvhWG4N2+/DkyoOzIUFPZnPWF0WoRhb+O3scTv1AUWY/usL2l5GN69MatfISfc
MJCqYvbY/ZQNJYSK6Lbh2/JWXHM37T9/LLRvCip20i1h5Gg7s3/jZWGbp1J21kGv
8I0V2uy31vG08gMkUEyclCiBnZD7pBSk508IoUzQ/wClQmMP3/glnH0au6lfLqog
6aeFl3PBj6xQqkAKp1kM7Ez2VeYU97pTo8CN64i4upuJqKKObk/Q7E4bQM8tNGDr
8W+jt/C3Vj2O6fYIr1nhSe15shE41ZcdOD26YaWkdvA2bnXjsO+G2DISR3NV09LB
006uLFAm1dICsudHddr+8xQEhkJGbdW3Kl3B3R3g6zkYdlBhTTwBXvpuPD9bK8Pg
PQ2BQ20ko+/owE1lzkKbvu0yi82fKdEL31FnJ4crUgpIknJbRm1dvE2lelaJNmsg
nP7RtQ7A0wR/lR/prdrw5Ge0GE3DB63M6FXjL49U3StEhunnEA5djlgkynHdTPm/
ES2l7ghLdFWlSUla45NER2fi1v4hWH/Mikfq8ARMjoPREuqjcHdqHQNYBtO6k6H2
FRJm9R3sNdlHxz46eJpW2MneG3X1MbGwexRubGm7Zdhc5hSXtArqlQK8ODFa2WGx
vDLQtA3MuWqj05Sz0mWkloKz2g4yeIOzh6jftJBe0GvWFcVUQKiBasaXmmyw+ERA
YgREiMVoOIOvP1cZjhqy+djbbQsHOmmj0fnaS+UI00fLdwfgxGQGiyxKLaieuYcn
V7BQzFrpRKzx0pmoO35EQ2I/YNd0hzmTrhmXdOkO5SG6CYouOXX5LMfpqhyD3Oxi
q50uP+UaTRVYMzaBez1UYuvGNHM6lnXtwEqXVuI3p1yHHCjn9UNNq6mhPqYAk4Z6
6phk2zCkiNEEDHnb43g/nylu5JEtCxSPGaJtPYclw5+UQ3qFUmHELvHxf6FqdWLE
JdOe6DkznkFR+9tobEZqyRCVJ/5raBpfWdFn4N+3GNx7H5bvH1JNBem/OnEZiTNF
/mweihpk2mXRFNYqcvjABN28Pg9BxUc6Pca2nK7iEhV2SucxwtVruQnluyPUVN/V
e5C78iaIdpLqPZkDmS32WD74b+bRYnJx8scVxYxSbgssbn+IhWOxbnAAHI08/FH4
BvOY9g2fXqT/+YgMTxDnHs0ainOb8YqTipgZK/GtxWFNk6BDqhTtDqvqPrIHzAsD
eGNcmCchHLtR+kGjV4II5mvAVlFIQAPR9V4AtLXLWqikPtRHY8z1+3nptpELBYi2
MGWE4eVF03p05Nwdn3uiTYticpGd4mdmYajC+34poGyebD+7c2GZ8Ww6Fu3JbIg1
y5qYhivuY8s/3SS4KfpqcS8BI7oZVD7+GAWPb2DNKh6N2GFE1rclayE+GApHJgG9
TNZnl+15Hx5gdznAR5XLaa80bpvhj694CaY0n2cXx5TWh3zTENj0mzh1KVLF8nDN
u/GvZPXPnyE7kgrmTeJxpJmsb+NGB5/o7zGvALuJrP/9OHKrLw7OKGMXgl+cC1w3
q8e4UqmksiUO1vlbVL5anf0Sp6chu9YuxrLmCxwlJXdkRXL86NksQADJbBHSHFIi
2qX4Hf52y3GzAc6/sUWiU+wIYt6AfrH3nsga6sZspom6idH98PJ1itJ8PWrlAiDN
HXF9aVPi2bgDi1LxlNI39TxNw5ehnEqsHN8BTGW/Ns+S8i1QGOAUDvqgOXEzBGmx
DT6AQmHelx00BDi9VhN6eUe2B57ewxw0Yx6ZiL/yfkBFaMiHze0GvRP9+4dAjSWc
nq+7ggv2pM+mU3o4eZKykolDISAq0FScj2j3fHEYws5WwUeGK1e3Q1bMZNUFIa0A
uhw+NSrc0Z2lOaFB4+7jgtPsQOC2yN7LAmkIat5VL7ZApy79jPLd3+wsq11BBYJb
PZKz5/t8azKMb5yOUVT7yRBV96G9dv06NrwXL+4hWVtovxZMr4/yIiDaEsR9U1Ny
+eeOp2JWda2VWQXADDhUckJRWgHat52tCtyeuua6a136UKhTUwICkTOTKUnXx42h
0aLCZCwFL8w7foNIDFZDJUsAO7FWDCKcZmUk0b7B9aUGnYq2WATBHVRcyTWK7xk1
yBj6feYCQtlymETcqFnGYupfwD9hS+E3sZB75up46spojuEHtKmdTBKkG3pZgiIb
9TPnLEbqwHKZh7c01+84wjotVY55PYpUwtTWxX0YBiQkGwbunVzSXsUdoFGge65w
BD0kvc66FZ+PxZX8BmWfh+ao9jwRffUTPYS/KNCF9GE3nyH1i38BTT3HmqiIpN6u
noroYrgaWmxKxYda3aHw4sQGdTqMuFFLEEfF8/BS6EJeb6X8YNdIDCL0TXSH/I6F
RburviB4l2h/f6sugzuO3+CK6tbotmoa93xlcDLL+YttuD91RSXNtncfUUY4fR1i
YajBNZD5bb26HZV0vjBDqPJiFTi3kzGvfADnxPkGAwnCA16MpEo+oKY/igDo/+3w
cRdLQCqpRJKmQEuNiOSnzZEWgKEHZERuiMffinbNywjslKSCDynMwBLJ62Y5Yfrl
gjTGJF5IvVAGVJNVImhogkm6srIzTfbk4gR7aexHEyfku0xaFngwbwoWz4CoxDUf
RxoqAv/ieX+o8KHR9MbwgWcaiKrXPkuQr5rzY9WG4XA5PnWHNAdWigySEkzCJh8+
2pwUdqgyuK8IC7AwtB/vqfSg8Ww8sND4pKlcIs9QXtWu8a2yox5x2PLRvH2SZrwP
tINheCGobQXtFCwGmc92Jpn0rDuYHsB0KKyHHqRvJRSmbCuB7Law2lrMCzyPCwvZ
7wPrOMrYB6TLqfAZgxF0+XgN9Q8faU1LanjXuzJktnwcl/BWmslirlYuyEZ1Sz6f
QeeJH9JtZUdlo8XRFKVmoaM6Tk4xaYmQfVbaffbpmY5VaQ6Zs3o5EoSvPDWiK9z6
KkD0U/9zhDuWREbxfxlHFOebZP0Jo5TW+mR5Q1dLD7j6w1Sy+aOO+FyVcWHZchoo
wG52EhGda6/QKMJtnBhKB8RCNCNo1dDfq/xxSaUSY4TNbjUqukSfmBAHNPmChz15
hODUweFlSDM4hvt6JHaRXJAuwgiDBk8DcMwLFTzJfrSLPrrNenhmiXnq3p0+TAON
yNgGlAM19SIUCfB+9arv/w8+958+qPH1oMPjGdEgyvU51y426O8RqbssMWT7YELt
mT8i+zxGV+jEpdr+/WUTMO18IBxMMuff1BY19zeceBkQGCAODhL+DylMPfrOJLEY
Fb2gKdWHejvK05zmu0cew8cn6TxNhhMOWRsDoG3DrmhPHF/xUdSAAgAzLAPVyNas
HEqjSiBvGyVuBHguj2bcGhCMh4x7htMWzd3Tz/gmLQ8D/NE1iQSHZEiek9AH6hIL
FBRXKydAVhLw1rqiLHm/pFxtDO3lorJDASWWugO6piP0TX7rV6DZHX+AR40Ts0fp
vPUvA/OpYI5v3FyTrs68RTNJ5zi5LROVuH463S6oHpdPaUOSYaBCdffcEkmSd0Ka
GggqJvaeLIc1n6Oj/VGei23eX3K45VAko9O5eSRXXiFCGxn72+lF6G24KkNsNff0
ceMORP84bNPzAsRVcUtCdEDIbdDCKKelVvxk0ZJWmLSKbTzUFh+WwX+J4EmPxjtV
orrvO/em6L5I8264kAmlEU4xyucXfBazpa+sKydgNJOXl5NAaR0l0/wdxfFe5cf7
xruVcUMJYjD70mzj7qp7xxeOpfh19sU16U5L2ECwjiJVrFIFhDch1ZH7aRiFISrs
Be0bBf0b6Nmr1HX+R9Qa9250WbDHUJBwX+tostMktKY6PO3WPoRxZK8TWG+eRZuO
GmEHdNB7vCB3Dm+5COvx8Ajl+1n0YLSyLE5HZsq0W6wXAOA/KwrrKwGtekKxnxAQ
aJVwWcIovPh4VIqPQjuXMjijGsSGz/n0lsObOGsP8NPdmPaBGuI8IdqOx6nqFPST
tcKJIZGYNzxBtlNHjItcgVvQcLXdFImndEmBkuYPfp8gprtyyc4D/qG1SMGFsBFe
vrYoU1o6RxLYS3Qb6OO75sNVmZXQNuYeLQ8LXF3JQ4phFK6fgv0dcWl1YBbIc/sh
h83C+cCzbEa1KUGIjg9TYmWRuIlwdTNpWvhOamMf/dAsFQnmKDSEbM33fuRvOALX
0Sg4BGulbhJAvPZmzXkUHsFELUOaBVh4HKKut6wM8u1gWNU8zwoO/2tuGuhUn2xn
jGW3S4Ew01USrkgA1opb5XJ9Fas8WyUzuiaR8+6HPUAJbhLfwRewbJa52tZP4Pju
ybIW1Sd8qChpoFBG9JNhmfew/xchPKQmYSHeVQ3E2K6RYgsviFZuPNC2+nIYX1TU
yOiuMzuE1F8G03v0d/uDEgQG9hZrIZ2eXtyzc5u4t5qJ9QMgR4e260esemUAclhB
P4YolszZdCKjgN8k+ePgVLaeBLK7Wp5V9yqSiEkEi6FAcRbph/2BOG7V0T3p6vEp
xwGfXiZJ8j1LVu6CFGImAHGv1lMWyenU4I5igj6z4fMYHARRVfwh33+mLWFFcdLx
IH49YdztS2PGz/qfn9n/Cvy+ff/mp4BLH9SQx6ex4T6MHyyzYNrQzfRoqXW1y3Ox
av4LOz6518UhjHSmee1kTZGwy+ieSrBFfpeUiPsKh826yAt0ToUMji+XCXeVuQqM
FOpW7Bnggk07a9lLW2vP27hmnkIWznQBaU1UxBM6QCbsq9Eme4K4uhn+CDHYnGfC
H7tpb7hYDd4YJdHdPkmZo9PQ4L28KZvVbDAwSvUcmqJOJTXUE2lzO/MwWEc0jMYg
Xgb7jg0lbBrZ0JryRcReqEYupn9oYo7kL6sIsx1KtrxvDCmpVlspnW96HqmLohzD
DHpKZGoTusC0dfkei1M+KKCPfxlA7C1WlN+oeh51CH3lCk6VAxKUTbOivABPWfb+
JqfVHbID9Q2UEO6KcH8OFE3MsUSJYepKrGCO3/lt64o+Zx1+qRfFhO4ptHC/Vw9D
tG5nOfHHFB0fy0vnJ7PIVr/eAqRjJO4kYHrqJux6h8LauENUdjeKybrY2vstUxKz
yCMemhR2O4F1MJJzBEjL2C53TOMIxi4fzlOf/ligA1lkTebNcbP66USMfrZHdWJO
FKy3l6NffGAbZJu64TvwqZuZcN2kl+PKWz25KO9uWSapulz+ukNnQZ0gzL0SeMQs
7xGYbL95KJIb1SOh5d8FuxAQ8FDWaJyiWN9QnhYVWMb/tk1s7kMdYaXx8qyvYrGY
1I0EqqbCdQSTNPVZQ0KD6ab6T0O/tNSetEHgqTBnsrWCENhFM4fIgTf6g2iIpJW6
PCNSlt16pc/kEoLbBo0gXkq14S3ngdstRK6eC2g0Q9amiQN0df6uDJygZXxT6rwb
um2TRs2fTNNSSuGkAo1RcxsUVfZiGiJy18jxNxyj/0uo4sLq9HYIi7/+Vu20/0+7
Je4OuOa8OHwB7G4e4vmOYnvz/JlPYJ54kFCuM1mQ0FGk330eCAoAjdliyk7iQOko
n0jkANAZIZzxeHKVsnc2n5Euhw6l2Pnq04fTcObOYuvIEUuWG5YrAmJkNuBb3l5a
nIjUyLpQ0S0hKKe5M+X7ee1AxPNHcp32HlBlPfmHh/uL1To4/PcHMOA0n/+SpwpL
Ue0Z6LwLMaU36f6R5d8FxDWav9OlffTeq1BmUKhHLFNtq9J/8/GCy2bA+c4Jp9NL
rRTi4RqmF/yUnZFO7iwEr0nqruq0n89doz7JmgDvOmjySoGaNhbNmaH+seC4uEhm
SgWMoSqM6Cxd2Ve9C53kHnLITR1DPafkr0jr+B/6M40n5aHfEPXh+VTTaU904JjP
wSvl+dM2hjgFBebKEASww+0F3tygmFZHyhdqnhTTBk2y6Y6mIIyySpSkd9gdt5VO
0dMLI0wSSPLT92uz3pjF4MZIKsO3WrsIypAtnt24z+xxNt8V2RE4P7hrDfKuuAFy
1YRYwVw4Vi/VviKp/wXbrH2t43QpKzXM2Ubx5266oIBXF8IMZYAg+dpPcZ154S6D
QlVnwk1lAwdx8cm3DKfSYoy8mTbWvXozDvyhuVGVDOD5sbeTXmMpYpLt517aY1aX
D7W0A1kw4fK1qh65IY61f+wR5tcUKLf3SxxWhLjKRqA2j+FTxzok565tIGYSYfCy
/KGfkuODfvMbK/+vnmR5TSk5R2uEWMROuSUUFW2wR9WBk+nfCDCQ1f1Hzjfv9Tz8
spe5SS5hTamp3LkiT+AVTg9mWzEoXPDVRFVL4ML4uCy+ZW+AL/xbwo/IpzAFGer6
csYqC0oG1IuMKXf93NBDnV2U+22SJRr2+iR3xpBNicVhBM8PRe4z4dRaMpaVEmgy
o5YTDtSnuAFDpvys2HS7Y/4BBrKFKLrgEq8Ppozwbb9yKY+4x3xe7bO+YAM1kPAF
PhqY/ZARlzhS8WbQjqgjDngmnga2IqJ7qHtGXoy/Noo51JCPieisDh8qa+R0N1A0
cZ3OisZiZYK3Y5YgDc0BtHTeV2saNvzaWUUt58r6rOkTnGxXdPM2j1pL7PfM2cDa
4YehA7goWzRb7OwKyQaz9yyt/qEp6VEDZG2no8AOGh92I09PV4GXKiOucuPhemCu
k6keKl0dvEfmwxDd4S4YzV6Hjc1xniSN96NapGkumu1lyGZgCxfNzZOjESLdJG7L
F6Gl+PNMiV8H1tSmRkC/K4YgSi0Xr6ggv5735heMTcpUbEexoo/vIa8SM130Aqdu
tS0RgBF452mZYiatA/OHpeRlwOjR4IAZFQ5nN1qKs9128TxbMuBYug9Go1z7t5CH
iCCiv9oXtIZDQ9rE1glJMLqSBdFv2ih5ekZqMvcRLYQ1m62oO3s+F9m7YhQ9qxJV
dy6zytyQPWtFPNv82fXSZZ2ZyDa++67UYbhwLVGaEbWoshui3LlbIYy+HgLYAFmV
4C3CHR9g4Rf/3L8wlS7ESO9RpBNXU1miKsfc6T6hynfvteWWBG9zL1Fe8LhSAutb
DtXaJuMpwQTuWVD6NzGzKmWekSOPT4BSuVYXH/aogARd1aOBHDtSPBOL+1oOTY7N
rlP5LG2FwUfNRrolxmZKV8KVMDShl87soN7g/1GtXe/x1bceul/I+VnDBO3s3W/N
aHQiCj2+B+Bgmon+HqQAtKuBpDPUJpzpSiAZ5ZegIJKc6tMS/gZobNgxizaFHQ1a
KasFyd+cnlx6IDln8mz6Q/D4Tkbtdd96qbPowTPxAQER00LNtjAH4+Wwbj0thjSb
jB7WqMFv5iwEj+bWhJk/YseK6LvFWdUn4m13h9wVXr5nKUB8F0n62ZCfiJiQHnV2
ri/VgHKuC7KaY4+0Cibr9qR3Q90ATssf2rwUUB4dV6Hu8m8gPURKDkBBfw2HEnjk
uqs+wu1tsAVy5f3wXgNOvsjE+xhDYyBWZcpYv9ypc3K+FwJyUO7DxAn50KNN8uov
7SiUBsxurSzg4QqKuYH5mUV/APsUXBYFIuY8yFrCTm9kEr7ar77+Vp9JeuK7iCES
0ivQmYhaymUJboyq5Z7UwhmO+I5o8lCvzHSeyrzUDrHzVzUMC0eeDwKFQmUhAktd
ZjhQ6CEXLnjAYKZlzXAkLtPgO9cS/afQlhodOS5Fdi16eN/8pOXMp/7Jp7XQr9LZ
FpugPKzLhwlrmMWZMKKPkpFRfEnrrxlkeNQr8n4kL21wx62nm0R5adFwOSpkFFpa
RB/WgYEBQdb4TcioeWAuR/lQ6XMb6tPD18IBsekDTHPlkSEEePtEG8XU6Mp/4WTb
d2DGiIpy4gmuV52nHVdtLsmsQMbJw904KXdVRGKkmgggk45F3BlA5zvjMVp6NRRQ
GgNgynWykJB7Rk3OXJ6mGzQVquC+n3Cuocl3o/F9FjIetX862Lu6PlRu34szIWlS
kmRZk9Lsb9XB/btpSs5RoUp3IimUCrhmtpdthsBt3xJFeqwOh8PMC+YoL4eLoHiO
TKcGOz/o5qLqRHWfPAMV2n2mbuVr1f4E6D2DZGIck8D5RDy9BfbtbKck0Yu5WnQB
xeR6z3/tN14fT81UDJ4chGC9vwehA3c4YLYbFksMTsiqbFfoIMnvU+TZLmUE1gjr
d2lXxnGkN1mGYFh2TqVd/7SFS8/BvI6izlbeHoybBj5DD0O9lbiem/H1Jul4bUTU
BQ/4YI6Qgt0iNdU+7Upmtrq2foHn8MfpOza3bnoIzdofurtOcnXSDvb91UxZfQuM
JCsyBs1w/mUFrZJEGoE2PTDfYoU4cYpDHRdqbHeqtqON/GV/erpo1UQF9w6TCVT9
291PIK0olD78b3XGdrwTI5UP/ABWMHbMlyhKxYujv/4A8bqh7nSorjx/0fmYA4Kk
JnZS6xTB5NapetYAlDK7SDu+mz/DHawXk35H3z6ndoTETR9KYqhaw9vgPKUcXu8y
J67jQDu2gR1E+pt5DIkSegjw6R94CTm5E4rAOaSgDwVxUD31YgVJeoShAzphnY88
5LYi0oo7hxTzISrD5ctyAkXKmcdu7oM7AEOQ1m02vZZro8IxQioH0Lox/weEnUsU
e4YW1F8psJk96/Rz00TsUJNZo6y3XRsd+SjLRRB3KJYgr10Y/9AyYoiJMzn8nqvy
xthUzSv86UhZaEOU7Pznn/IcU/PGnDLoHNL4riny1aOi1B8irJp5MUVprto8YdRh
4mEPArSVCDzm7PhOhOftELO8bdTV+87ALETFHoA00YjFd0NSo1doV3uEVs3fPxfB
6iIb6boL1L7snq4n3qOijYtQRnkpM1MPq0Nq9Wu5TUiqB6aNm6GZtA8H2tiVjQ4K
3aHX8F340ePkgloDFdd07gfMwolOXvtj2A39iVyCeRFaxukljCl6A+kJw0hi5rtU
ssTx3kaI6Ci1rLwXWC+OZde/Fdu8SZlxFyf0f58jtQ7CHkfg2dPcJffE9R6vWfI5
qyI4YByVe9/NheREyeuSOas/gyVNci6c9wizy4Sy17ar+zJ14MRVlwBv8b5YiLlB
EJGV0RFW0IMXx2lMU0JEkYSfFOIDtS2kOlZvgJgchl3w88WQ/gZQjXa/38xwDhA5
d0HvzNHAVyDi1PNA9Pl1o+ZHvKBW2kD/0vHsxf+ABk5Jp2pRHa7jjkzJxLnOtNFt
Fi1jRYc+9qe+BHJwCn2sZ2P5uNgxjRP3Ag9PNQhZr28D2GpzWcM/QI6ZwUN17AoJ
/yaKl8U/mwOkmfRY7gKHIzHbQa4XNcuy4VhYHpZZwOIlcoDOBdx/kEaPJaWaHfjs
84gCIwSS85qYpPR4mMctcmR38vPOYONQJ9+Rmw3gx9cLc6hzr0faZOirFRZX8RNu
xKxGR5QXmSZ9Eq98Ovsy3q96+XZ//aP321ccn6UNYz9+aKpuTXaZXVdsyqJFeGig
T7a51hI4gBkj+5zaL+mlhZAekDItteomvpH08/MUh1tGHVTJ+AqAy13J3nYaOCO/
JWfGtHiXy2qInpcCVFG8ex7ldDSyCa6Xde1N2iJXKqrTN33QNcjfxB8jTSjjctB4
RQV7So9tNmAc0T1/1HyC7yCJe4iOBkjMkNA3UiyN1tn6ZJAEJvIV7yZZICk9P7er
bDh0gOWvij9XCGX9GLrpCIUppJsWDqqKk7bpg5njNuY7tp9twPxR+EMGgXXIfeR+
9gsDCZNsAvV23UKHxmd7GisFuqZJoDgI4yqSajJc7g+28cgvy4u+88mJ2ajBQW9N
txJo3Yz6pow+yaDDMIhRdMJXW1H6XL1wACCB6dOqbqB75fUPHSmWxIqwoztmyfGr
pheY3UzF4uIEqdFmMZUx/3SN/5tclBusqSZqpWaV9h7shd8XgenD1tvVgtNgOnW2
liD7bkJeRKs//pdVKfekRv+Ek/wxnWDN5tkdpUAOCx3XdB+4xK8MxLYybceeiaoK
5zu1uNE5qwECt2Wo0V2b56Lj1YcMdjhpoTXwpvXw8I24NziV3bVtjmKBkHa73RAo
pCMxnzsgwo7Wic4pMI0zlKoQMYkgyXZoaxFVCZaOT2evvkyIEAfBXtvQOr1q3+dv
GtDIRWxZntIn5F/E9edT31x9Rcn6QLmKv01xBe74RdhES/X/7ckU8UyZSvftq0Rc
SgUQi69Gq2MSg383JNKePM571cZtshUJCC+353ujjr3rSvi6XzfmPnOUIlYe8RPq
gOGoEgAw/Q97yku37SI2v6xTD8hWK9WgE7ZXzIIDXt5FhZGm7sAMHgo2b7USexcm
2ND7P7uEt3kHko30yx2ahu1fcN/fz2+/aYnbeCo4DrYT1DAXFGyKSpWEFEnxejb4
DivEKSp+fo2QzZ89mFHmJ1n0HQEk32otrBXQ5dK8ftFZHOKuj5XjHPtYgUA8oY/X
6q2iUy5rqKQbq6l8RpP6L1RBSnQidqnzASUMHMQxl2JwHB5Y0b1xVe3eN+05EmNU
gIZ20D3YZ4D2T1yMX528JVMVyCmtTYxuMrYrusS2Aea/5fMvea/SAyKkkjheEkB0
LTDhfBQgsLy1Q9EeygUBe+qKxG+Ie2ml7Z+wOKqLQo6jIXrwiqVpK1iwNh0eXsNl
buF3W4hoy195+g3bjFf6pUzWR0gmvx22bPEkpTTU9f2CaLNyde7w3d4pmJzOY4Hn
eicWeqEmTuS7LVxEdkThTpurDU3B+NRTtz/mJxtIrqylbgrBu+yxodFYrmc0xtJb
XO/iZ+cLqIh4dITtNPOHEqmIDx5wJF8DwP39z6nIV6eTq4BCXx0vfM49YvDDATCO
13Bozwt+wUrxv+auFEK8YQoPNSlFUjuEFsLxTkecYgZ/oAzxNKCDs6NYENMM0bVd
JRN8X9xs/nQ+Ti6sBwyIGfS2maiIJExysIDyORsXEhZ8VRvJfOgwweV0X4qXCXW0
9VTnvBgAyM8mVElhW2+QJCPqJVDQUW0wo9DSFFHQc90xjFcROZZGKPtGQN0gsDPO
k6H5SurguxeCpmaphRRFy1JQvzKZDkLdX36fpr8edU3rLLFzlrm6YTjdmHiACY8W
L5D2voh6qpr6rHJKhhTZ4rkIRhWLAu70rIKq0NJ1SDm7UdHmIBEjQTSCbzZazpre
Nc4bMV4Zq1AD1FNVt8tII3tvsQ2hlBP7BTiQXYF+CUhHET6bn4J08x+UcwL8+QDL
7rKFBHEOBiTJP1fcpx5JlPlux8lMR/r2ouFu4VnLn+zeZ0+gLjSSiiS6d6WvTn/K
zCB1XJbwlqo/ckik0ZLtkcXa/UmfYYtNx9C+5Q+DzgXrP+w0ZfuA18TZFPI2xvru
tbqBMpnmNyhPL+Jk6V11MsiLPfnVDVKpA3QoKygrQ+U1u+9vq0ZdLZBgqQTXxZ5D
rk/0ChJVQKO9GFhlfJtWknQPwC0Yv+HHcGHzQtVViVNzOE0d3HvqG56AaupmthU5
51Nap1AQLHQZ/qE76vE/H9SgL6PD63caMituUhEQwyOjJwMvrZoavKoIcAEpoWRY
XSgf4Zu/H7pJ+aM+/HXja1whdurFmz8PEUrVPoaszMWUecGukPEmuNnyI28ydtKR
VI8b6qTJ66SB+Pgyrw2Xj32mkVUFTszpJtqnBp/yTpITMOignPB2HCUdirbWtJy3
wnn3cnX+8xmi9+PJXcjI7JnwCKjLWPAYb+s6Pch02BhaVNmwjUkOQExQ+ilcOBWw
xR2X31i/BLC//zhgQlB7buUTxT04M2L/zlC630cd8+jiIqNJPtu0aQ64e2P+d2PY
ftRZ25KPyuu/E/hLgMLXR2OA0Terat1r+Nc6QzvVB9GBUYyJxw/3URS02b4zniPj
rK67kDVJK0ZiBnQrXuYIymQDu2qj6b7/4HoMg+YvazJ7rU2lRohA6L2Yze2sn570
nfHJI6lXrC+4TIw/MiTnGFmesSUl84uud78lUJwcCPXJHeK+nTxHPMJHhjAowr6A
WFO9AEDlAFWeAO9UScmOP/ORexzfu9ovppoc8nEGpTWjc0ayLXBf8K1xGk1JJiSI
2fqlM/S+sQJv78uG4h1R5kZnRckRvRAxzvWS+WfozDkuEHm4i1es8O8SA0J90bcN
aYKuKxtYuE1wjnomyvMiUJnjdWxEMbzMVzLSxPLl7GHBsi3EaCAboeyPH2Tx37wK
IIXCikGhJNuST+8iPEiPKkODESVrV8hTA8yDeJJ3ci8OERp3YT6wACGHwf34MCYI
DZf0TpPZLtNYiT3V4Y027Xbkii8651c7UQtYXWXDRlQ+LcDsDygDvYMJkq1JK2mB
9Fsfr91UB7hEkoIRHOMqp5gSMys1eUkYIkazZiDenGyVENVmtThMpk0B6YzqecQi
IWkxvvRBvJNfVvy73l2oMKpRNao9RLNXdX4A3D6gPjesv7qR08IhKfR1n16rtTsA
Mu6OCpxUGHvS/WuKuAL+7IAoMH9SiC+kbAMxC6BpnyE+Q1+u1AUXZtcgx0ieaCjB
2JRw39oQGHt63ST1AfmkbBBV4Iel1iWvR23quc2Qdxwn4iKCQWzXKRpItd5MpVyA
MKnrYsDvveSnIOCEMgaV9P73jkbW9whPn3FCrmv9Tagc7y6HlVGb6nCuQyd3V3LQ
wd8KCM55zCwRFvT2f2SBm54r7p8Ti9h/XaDOofLrZwjRI+s3EA484tUOT+BpyPR0
KWWaqzRxhMnpcERKgiUI2LZWq+eeaAwM4ubooGEL5ZQ1BODKKtS/3NQy6X7XgmIe
L22JT61wTYE/WOSHSpqR6xk1zxP8FqL6UUTWydXnglyrcjpSxwMO7NxqE7VYzNsu
BSEFHeNES/htAiD+p3iU0cLnnTodneJBHV2p7ybgXMVIbGz16U7Dx85NMy1Jli8L
AIYRgVbx8QUUxryA6vil1TWyaS/vH+Fp0KIljGHDhC4GXhUD2DdvhfJmSr1p0Fze
NxUxWf2GRl44ufQZuZB0kzR65Q44TzRG/Oy/XVm3vZDJeeGKvY0Wm9rsrAQKAi76
jXAuCYdsTt3iDREJLOFuLIrAaY+kG+nf3qGAsMDRfX1/Zpz4obHylslG90n2fZW8
Lbq3YrgCviGNCi71BfQ+vNxTjBuf33ho0EqNNv9Sw4nGg3BbXCuRQVcheSWXhDvn
brSrcrOMJETCkZYuPx3aEJB8co0mnhmcUBbfPplZZYbBqMY7u43vIViwI6o7DE8p
Q+XYT+J8B1HCJN3XVI139lmL7WW5+ZMVfhmytLgmwMTd+HT9obVp0ezWakbjkS7p
KM6YLtsq3iNghMMgwN7yLdeOY697q8G28LfljpP9x+wEzfsoCl48vnmGI6neFf+N
Xi48PknXTu55ZFx9lEESHdCCoYmsmx5VC33ORwg72f6X5y/rDdc6sm3wsu5/oELK
AioQ17UzW7qzgzuqHq44AY0rKTf903YJS+ggYOLZXrqn+j7+Dq4tgT+eivhRkWS4
RbbOw09CdZKWFZoDxKmHYz99kbTm4nW0lv77wdQwUMJAXWWHV6klmIQ9ovvFHy5J
7lnKUnlcHpSxbIeFRSdlffTrwxWykudpgD9U63lB6dbR5O1fOJHkmQnrvGcp+ldv
eh1nHQ2oV6A9lZzeXgfIM4dnIHz7CEagT4BrW70xri9DP8Hn6MMcBUVJB91zg9aV
upiwkNx8nSVIhvorowXRBpd2K1xMaNs7YHKmHE3lCJqNSYboU6bhm/1QNE50W/8Q
H1Fg4BPAaiKVtlSdaIpqE3Kxs6ZfNme5m4R4N+SUdYb8xqYJzgHf8pgzXMOEtnnt
NHyRKp1GJA4wwUIjbAMl0aSANTdlthpWIDxWXmK2m/rNZ5hamaij4j6aoAo2hoFq
mdCa19XRJn1DGYoJ+a8p5xFLNOGSDT6iukyr20jpMk9c6yYmLoGmFu7EfZKfmKlC
c+Limx+P/hcxe8OQePU0Ps/cHr06/pX15qQla2E33LqDFqp+c2eERaSI+R0YiqNw
RKVmptFuaiZT55eMAyGSTKXrJANkQ9KBxs9QD07BA/OtKHBrfkzTg9OBejs3xe8D
8/38yo1oMRXECd47hVKEozm4rn8JbFr9CLXgPVxzsuwlyGbXDHzRdeiG8lI9GJHR
xEhpds9m39uzhpUMiKckskk3nTAqxhWHH6tC6Q+sffC1W1Yb8RVawzvP1ZpBo0Ts
fDaX/EiOGT1lrIIMeXEx2ywlQQzJFvw/L0NdfbUS9NCUj79Rxhe63R7nd00PCzsd
fQ/lJZNBFK4cV5rPuqa6Zqae52Z4Wu1wm7fSlICPZJboJpZlVxYbHyzdHgT+rbA/
KkkO9ogADxpf0J5Iv7KPT8YtgXUIIpGvdQ0sGxh1U5tRSnT7RDo3gpjphiVspfKM
LhvJoBN8IN9+hHDoyonDeTShwbERvYv9WghDT5hstnbSyi1vahIAQkVuMmnMeK6S
ioRRpESQbBAY/cHU0zES8X1D2Ou54jbSgfdvUpEqInjRUgMQ/WLp+szVp65bRjMY
iooVE3B0PU3MSFkBOaYZkNvt5mHSu6N6xEmVwAlqJixjCJlR7tHc/Q7+fG83X01L
0k4ailX2bDFKkSo5psn0wYGv+2NXNlg++EC+w3pq0bq7B+U5aquQ6lma3VMl72Ku
fETW3j9XkcT3MVdOU0j8OiEC4x5uC67nWmWVz7Nm+ZWNtgsLEm9wMK51+fd8ULd8
Dv41iv5k8WP8kMPe0h3lo5RkLi3KrMdhIi0v/qiG3pa/uRWdHM1+2A72yfZPVGQR
7bKMx5WWvp6Zuz6lkV0A09wNZcoP1z57UR9UtoZpMb8uuJ8KUtQkLDsZPGARiyvq
THUs+Bbx5ow1I/vEZ9iMkLjr52FBefblefI8+E19ezT2u9r9T955oGbvevWhBEOu
DtGpZxpIwHLLgq+aC3QYWxd59D/qdYDN/nU32gnWGgi/WZqWZ3Vfj1eE9lTvcD4w
pHUciv7ZODfIqIeGX2Cnnho1HFAksbLxnl1qoH+tn0V8BVx5hxso+phB8LglIw3j
p67D76KDDmnduMLpe7gp4ZMYHBXQV5IwO6FrAaG53K/M2Sp+UhZtcJi7okiHj2WZ
VRlpRrS2Kq5Fqlql0b0j5ocJRU4pKxgT8otwVgJ7gubyzLVIxgZoLaBbqLkfvheP
l/2UDoEoU58PSlTwF0VBpIK//tibCrpULAAs91K6qkkg0ghW47Nc5FWYHHHwjMrh
qMgDou5fgm9bd+a0qai1sNabpbSv1odHFjVIYrDp09S3t/HbFVjPaHOd+wlt/hNV
sZTkVnxpWXf1QR9uo9OOsWQZ/+lQXyr6Logt+qTC9ROZsKd1scFPFTtad+xnqF2M
bmMBQJBWf7/3z9i/4jF8qN6pyOcJ+dGDvHSBa5RFJ+xDFIuXsF4b5d0848Y0lXXX
PWPoKVsgNJFWuAP0oCwxcIGFmr+7cCZG9I7aGzgLnDqVu1cmWsuLcGlAfd72+Q7s
v60hl+F3g2EF9nLAWqR5WZmi4jnih+aSZWkWA9gUqltnyTFnYS6i4mRUV9q33rH3
0YHlZwxR3vmeaWrdU6XZkByffBcpLzAl3SLzG59hToZYyqZhVQ0LGkXBcWeF1zwI
6ZYOsD0XvHT+oobnU9uPnpBs9pXbQfxrKS8etGo3YjJloKbIzXcIk1/wYN6J/xVZ
Ut4iqA8qvshBFelnOYCC9FGSFyUzHEpUunM31oO12HGelWdkHjJIb0ObN/3HE5dO
maZhO3I+9TyO15YoGKt4VjOEO0oW9BtcTEn9RF61Y+h2PuW7XwG9fSDZbQmCe72d
e+eQFGPWltdBy3kVU1W42+WmagYZxZ/aAVGVsPyQ5pH2jH6/WAr8S9ogpciHryzX
uXqlFWkb6YdJS7C+yeJOF1pUk5OvMqDsfwlEDKHtFr5b0Wf/6zYSv36Yswq6tgMh
N1CM6gDZY5fdeWlm8+amRhifkJ2LBAO6+wKxtMS22s0lKeEYobWKjyruEiv0Fq/g
dKWSbkBi5njKTAOldEaN6L2c9J2lyG9Ht+igrSfxDd5fDnaC9CWh0AmtvD//mudQ
eHcfciB+5nNjs2mdtRor3p/q2vJ1lRLmGDIvz+gau4PWLEUfxjctjMt+D0tFsixO
1riDQSZq6SH3hraTxRgA6Jnk2Rjs2jzF+gizPIZ0o3104VbDG/Vmw8kLLs/otS0A
LvdjbhYcjE0V+KdpZW3mDzXe0ts8x3dk8yk8GQSnGOZJarG56BKrU61u7etiGDoe
jM5eHKve1HrlMSvVw95Ftqosq+a93uN564K9uJuRhleCnijjBLWb4kKAF0FjTP7h
Asdj7WUb85PkhpPzlrD1F8CCBvJ4mEycA/+6fF9qEk58dr75BF3YzBPF5mA8H6WM
xFE9Zlnnce4C9JU8ihG0Ei5kgI1tYxRV0rJ/dbmZ8Gn48oHGSEyOmEOm/VR27iqy
+awz4xkJWyNmBkphTEFMGp5Lc05XVVR0Z6VTo14+8MGqEBSudbkkc31DVs/VqTZG
m211wszMxwTq843IbNZ6jke8njHsJ6PnT2Fnw/PaZHXtZWo/z5et4ShzgJ34/QpV
mv8aUhVdvzfeqqK6YY07/IHGSuz+b01Vtsr51Q41DNPhYPK7mm/1Na8WPgWF567p
cKL/oz9f5OGNF2v55n1sHV1YBmatv8vZA7YGSUBv+FLptBV8/vcR96joxdTIph53
UnkkYXrgNJiRKvu+7cd48GOI1Yy014MyACufjAYYwNvCsgtO24P9HWMbpFvDzgWw
aPLAmj1mda6dE/BgFizI/ef5WhRIvbOob0HL03N06+0n2lp/2dcwS0K+PKcsK8et
yB0r/wy/qcFXd+4YgspuY1B0D1pFRBtK7o2n2MlyOXPCxfsmVBDUD01TYvLv28tV
ceFJ23b1wCeWMw2gZW5i+Del0y6vul3kQRFQf5EHF6Ngo/s5SklU6Ta03rBL7VkX
23V4nKWNT5JsqWhilHhtq+OyhB6RnXtDmw5KslaHwLGg6HZSR/6+oo8SsDHHSh7G
WW6+Y6gVSD0DmFfJF4FNECTsDAzi++OJGG0aFQeFtJWeINi2R0y/6VN6qlc/gRW1
VxdY74idI8NJkRIH/KzsLhkeFcSMaC/MnlUxMsKJw12IPjDhN630D3pX62SZ/Tve
MVstmLFA185FDUxDho0CRPm9XCve7kqQvaIzOxcHt7wOEaHS8lP/6Bnyd1fhSuh5
y0CadL767/j1mo/Mk8UW7SeUgqPF2WRV00GsSa/owpuR9Go8sYbh4e090JLgqUop
+G1z3T/tkiO7c6fGzEIHnPy8WsMZgkIaB3mIPrZ3TszscLTcrHPzCP8ynZZd1r58
fQmVdZs3t0RNh/XDUvI0KOwE025He2oU2RyqrKI6cFz3Itt1Mz33bm4V5bOGLi2L
fhNCMqZGIf27uJSImC+TgNgG06zR4HoXpKXr2qsHlp+C/tesPvux2gO3O4zbXOwm
KUqTr23xon9cEUHlT3BF2d+Va7qDBVcsvVBNB1+lSKcnX9nDb45tVmFG1S1uSWHS
OBBijLO3DJ9ultWJAdUtsS3kceYKQNzmJM2MFWOSoOhT5teu1q4vUNC6TXhEhdkO
G53c6JsoPevMSUoV2uruDs071D0jp7xyAl0cwSzhq/NqeQRrWfepfn40Dp81qwOp
bNbcPnzbZCd7SrJs1IOFpRVWOILIQYIS0GKr0JXNl3jh49VGnLhxaRFaBu5FmRF4
HwUuR4cmRrfuWH9MO46+rehLe1oQ683Tm/V8EtCKinsE0RMuCwSN159UJ0rQ6OZf
8wUb0JDSeRGFQlvsOWBdEy2kx6LUOyCdElrNPssCrKlzkJr3CG4ZOpN+5K7GBY9Y
3YgHqr0Dnf+PmWz3DKhWW59nZfyTfG9KpYhPyfwhvx/DWQ8o+YLfJKnwbDzEY4P2
vIdQVrYyy/Rlk8dDvP7L/XeIMSwQGFWczE84fkrgIga7aavNGw6JwGMk89pPYKKo
px8CNWv2S51ZsML1eD9zzT4eIwsFaz1kgU5JG3LoFn8NlO2880sVIr8K8VLG15aw
huuOAU0Kki0CXilb5cVY/yZngvA1bHP+lUC7Hs8BrZ/0GSPm1x5sM7ixJ5vlo/wL
vRwf5FeyyjzUTGnxPE9ZLkL25eB9qXW91UPIevh6d6vJmgcx4KlBMe38BC554xId
ooz8Gl/V7UuYlo60lYqVBAAGxSct26iw5qsCvTxQDLIqgcSBmfbKsNB4wl3NMm89
xb7ImFvY8u9KIoiFmstqAOPIJ5j6tG4wgu6akbzwVbfLpYe0Mt1lFeWzEoHTW2ec
YSB+Pn8DwS2mCAJNdjrxQiWBuJBYT++L3z35wI3MjX9hO531auvAisqkweWLHNQH
0IGmi+Q+NNNCZfKUrR47mhBeHjI1itbnTrvoWOcqwlrzuEW3GP/oq1cUUBRUDNWe
PcEVai0w3n1N8xe3WvqHk+pWbFeM88QfA9tir5zJwZmxPNa+3gHoC4DaLI+hLk2F
VBn6wzyZ1gc0cDd/o/B4m7nk/FvnsscenHynd0dlLK3bmHWHpPuu507lp85iyjm0
3uj5eGE2WbYrIsO/cuhkpHQkhuF7ONYq1J8u2+E+0w4R+PYgYSlJYM3ZResmwhjN
d4fqPKlAzH3GDIo5JX9RBX/6E213HJ61bM8vBnn+IqUgfWVcmTjLK4PqC22F/mIR
AH3yejfY12Ga9zB8ILqqGvWjn6sV6W19Nf7GI1Ooizi3S1hRjiFzJ8jwna2G4++s
X2zrp5oHHajRntrL4nyTu2ttuoP8YcJy+yBYiP3b/Ywoe3KfAsiBYI4K+vtATOlW
QrfobI1hdOr3GzDuXn4Y2tbkTT7Yf9aYlvsYpMZgTA/5Kgmu1Fx+/jjVexclDwXj
FiN2ycu3VpFzyzKsiJlnoKyvUPxAgFU5GDTgDDAU0zSVMlBGxq59ppTIgNBqbDF6
nIzMMPBYXcZjlermKCdBIntpsBuytu4NW7WKLUYF7Tuv69xyW8RhqckInxS/IG1Z
b6V6L+jR+W5FN7urr+yhH9sRgHvgyqBVHykIzG6hhwrkEAz14emi3KJy1O/KJWGr
jKtH6e4lb/Uc4d70YSvoxaLR9Q5sv99hHHPjb0xiYfqRkrxSl7kmxshV7sR1gC0b
iIFBfPLYIt94mkSe0YKRkhQcM8F1o7W5PMyM8qqcK3MXvMAigimsFMUx+5vZfxJ+
vdux52Jw99QMOEyoUptFTvTQaJPNwg0G/KeO3oUIa3cm1IcY66ct9B3R7ahO5fTB
RqA05qaXWmCpBQSZLOx/lg4b2FuAawJdMys//BvH0yesSvc/SvcD7C3FJ6F/GJhM
xzqNVwIgAdil3k6wLoUUmc9GZ+WKcIyNaLs5eEv/Xo6z48/KPou2NYGqE74fA0g4
KUwkkw5d8s6F2Btpngr9jqBCq/dsBeJglkID7zMt+X8QjTLFRvJH7T3D2ZaEBkH7
N36IZYRY4LVuk10dEVm6E4lnMctMBJ24sXBnqF8H+EFOgCquDYzIHZm4gUKFVk+P
rqvd7VFhhxyvwagTexvP+JppllUPlvcczv9ORkXcQpZ/deFT6O75N9UwXxb5oSWt
DqrcbkTzULWZ8hFOrMJifEGpRpH6bX+vlSaL6gYaspEH2BsQqvYY5BAhLv6SR3/m
VF563a5ekFoX2cFMA0rH0AGO4CxYz1Bnnf5/yl5xi7NaenG+ZlrVbstwFkRErNNw
hTIDhI6n59Hzr6vs+ZGMjNkIbGINyu/r9q+c9Wa4N9ff9xzJ0rcXNr6FcShQKqvC
uxXG4bY5BqrBGt7S5TsF4UnwoYb+OrVzBfXkqWzF+22Kk1Ju/t7uAFGPP76sSnnF
PB/ON9ps4t/Q14qAR6dU3s78JDcH8pLvRgtjG7ExVOhgPhm9fiUbQUINriWKmmtM
ouKbkiI89VQh1lMjzr0I5FR+O7g7yHZYqbevlhL+oQzjoYaRxUwr0ZL4sN8P9Zch
jwYGrBxLptss3CgH215zFklvyvdI+qCHfmS31oVLOGkzSakRkPaDLeC6327z1zvn
rfpfDoEwM/EkOCNLHuoBSPCUnkpglfMXe/q0uNIpNLmXsEo0muZPWLET0wXoEZez
UKydOA0BFcO9F2nYPN+JZjmxYDGmxZ/eWem9gUXTsuyOu5Snme65xDqCeh+YjPnA
y+XsW1NAS/in209R4ACOjniDmQVHTtt6TpIPBqxdBOkx+bXoIDJqcrLqM8I//KG4
NK/0ywxmqcdHYw48wkzxXMToegFb+dUAI9wChkbYAUNuyh99qg5y3Y2HuYjayNUj
sz5BaOKlRd6UPb4z1bm1350uEPnMNlHH9bidkiKbq17OkHn0AZcz5dJJzf9Hycxm
UpV/1XU3ESbDDoCNsVwlDGitFM443NmF9nxMbGhVhQtiIWIsKhDm5C8vxwB0GSTd
ux0X7rWr0Gf4T1mggsMzFSut8Ix9Gk1dsnPw3F7893fNhxDhrm2dGPwHZOdq1i9t
evwAJqGrGem2L6n9boNq9kKayzSosOULn69cKYsVDtSgCFTcKK77A020rWeeF3ez
mAVQ8J2ucmqScD92yInTTWrUVsX5CWWJXi9xTqfB1k844gxu57OkRRMUomT5Chgu
bufhaY/0qtbdZB3GL5KgPpBTdI3TjIfsJBtg9/sqnmR3+Zj/kXsPbZUQO4NDdk08
cgilWoR46fmx/FihrgrvpcafDj/u5ksVABabxTSNKoLD7KGDQl2AdjPtyKF+la7a
obVLxSgOwjRegeDdyPAS6mzWOBg0Yj65xvLx8IbXdsH7ivurWLmh2qthOCPvmJEN
67PoUaXgl+eOZQZwc8lF/DVyQLsiBO5Dbdzx145042aQz1QynMXLZfen/lzxDS1y
6oy7zu1ymMahkiz8QYrLVDsstoHOTnVhy5PSZ1+V4OYlttMKgh72r+4RjxiGyXWq
D2b5k0N2dh6EBb2UZgdv1F+cXVPMk9ZKY13kwixpsy7sS5qxf9a1qTHrv4j4V8Yn
NNtq+60A45E8BCaP7ItidZN2zmkWggF0z4MEHucbdh2JeZO9782sDLNVQ7DXSFVD
L7KHOEWLwLWDpLkkQouw6+gFf3ig4Py/7/jnxmnHz7+v/tEDPqlpZjrDy+8AZj1f
eKyC6VRiwhOGNfILZ4yIdNzHW0X+TPvXBKr94xecWrlkiPtcBQwewJyJgxFOn9Nh
OzkAjO0eS9YE6FBPKPh5MQfi53N7zQMkVPTV42Lr86byLWci951OqBAXDTT4enAI
lgJee7MGSYZPSfGZljyUH9/gAWNEd5QjlewdC1yCzSrn7vQ45XQOJrcdmY52Qyl5
gYCK/rDFDbAoOCrLcqqhndlUf2fjyCyTrisziqcQ0QWIl4FfdQOhbwxLIUFS1F19
NOkNTUCAtmbjuG4TBAS/fyjeabDD8T8VDdyZKP+zqX2oOfCalW4XduA9ffQn/4KA
/u8gblzYqSpE2qVkKxDt2TstY75tiUNghaAGDyMiyvN2R2DEiqgogohTnl80SkGo
XQELEyjCeAr2V6pEkQl8jWgIL8ZN0XeRrzUCkv7QBbFSwTjqfctC/GcEEnQGS93G
Vo0YvfyzNhuQXoeY+NRnT9+9xuhY5jG9iI+RQ6dmKBcw/O2KjB3mMzOZVA2g/Axt
iOKZ0aZIaAN2SOFjfMHqigvryXn0G28iBx3dfopb7Wk3FKhFqSqpdEvWB7sAg6L4
Tg6p6cx/T1uB/rsrnNX8SvwakROmNwmO8JGmoUMX7pbOPjwrnciSDzdQn5jwd5wC
dcMhqJSwuX7CGTPOpDn6q2C7QBL/YIfAwZBGtNJf6G/muwzXvFh9JN0VIoLHded9
UiUOv9SAkUM6uGUJIcJSIRFCKhiejfc+7yRctQSTECXB23dezxFPFtCaA5fmMEdH
FzlAxrvu+jB6b5dQcrlHdpTvjSGmDqTlXfDw4lOkcoaKdstX/lGePvB5gayIZC7r
z5echosz0X0lVmNgBA2sXyLB87vRfcY2VUG19GoAK50LhL4rAX+FGPLZwHQ2znEc
6ALrqio+7BD4+g6wyR6I8t1TpNTLf8nZwOlyleIrbN/SwWYPuahXzNxWghOTCfKz
4oOrD/De1vctaqbixK935w8Q5fs6XLcRfKy+PXdZuyts/EpZdWH0Z0wfYYu6lM66
sUDoqpiwDLerzNZLl6CwtkTztqvIxTb31HgtUmK5E0NZOgiGOyxa9mW4ti6B13Nl
c4t2ppfKhNUoO9dlqSKv0MVS34BQ4M98cc5KwVZWCyVrzJHhn+plv5xI0XB/nPgX
1qV4uvuy99G3nVTQQOrnNqZ91uIb+FfQ8wy1njz8c6mzbKOuIVrCjnSTnkd/0Ucl
s6vAYtp/FcbRag3noMaF6s0qdLe5QzTnI9yiWlLNbpqpWzpU9vddB4Fb1jWCWCmx
KEyfMsJjpjFjJbBt/cvfjVcmj4GuxykMPcBPBUM9LwvINOztNesmwPsm9RcI9eJZ
qj8bEvFYu+IgLNkifU3Ncv3jVO/6KFBxlLdshTAdLsCY4RzQRCZOoC4Ehh4lWbs/
WRxAz6LA71R4dMz7cOprqsgY+XFcYuhrKJSIHNGkBSR7xGB6/f0YRS+q6WnUiNpR
e0ugZMzQ6XqddSUmQEKutMSY8pQlcLgSRDju+ekzsa7lS62itL+4w1nkVS7JRgfR
9dkYxAuw+HGnSbzO/Ss9PVuQfWPn4tEo/XMTPyM/KsOyLCpkVOXuk6OFX7MpZDDr
/eZZXecc21rBAj+d8CQ4k69p75iD+JU86de4AIGbtNQF118HhnEgaehOOzFsZCBV
Gop7sCEneSzF2DRQ9+//zdbgDCPa4m5QsBICDCbMVmBwzrfeHuGo0EvATTmnMls7
eFr9IYN1KpV6IcmV0BRqV9OJR3bruLs4aswXMPukNmxopcyG/jCAdX5OzMDWII0V
t3XrbE1yiTg6gUrv1BtKxGZRU9qWh1rtyxY6xKTv1eQeCAD0FlPEzqgAyInaSblR
MB7nKleNeznRxDP2F2zU6Tp/JhLbeVwTK6YvB9B2yZey1Goa5OldLdwg8ERuTifV
Cc2fvggc6WEAh99FQ5fncnbeZImmgJ2FWQapxjbbZMqLeRlswy510w5A1chhuAHe
2CscibGuRmDNfiC5RpbuSuTdF9mLXUs+Jk1PcdkJukYEnqg4kgbIELfvMI8p8tUm
wAIMxASfSRVSSk0s4cDL4worX9XEa/JqXRswEFwF48OmSSrjih69sADaZwE1YL7K
/GJ3QyIPwhAoKdDAZc4qASPGf0d+IYEsiSTu8vjdefLOjd9wQwDPD2057QDmaD5Y
SuRKwMUJeTl24r1Ooqrq29dheRV3Y1WD6OoaQ3IG7kcLKWOyIooZQgX3XPj/8mhm
0V1h/er6R6RNdNNulO9CHV8ClNCB46nb90JwGtan3F1hNLR+2R1n7YRbaSAI5CY9
3RAevPqTEhWQGNipyTuELKcyZYaYppUGBlaZl/m10q4uICGNWwkQrC/f4aIENV0l
zzSMoi9AboZAxK390z2aTlkndAHkzJ7tmG1Ir9n4UTUbEhcCDoKQxtTI0Hh8t9ha
1ui1NaogoOEz4wwavx//lqIpyWLOZ8TPT0bCo+tv+x6MCr0c2BUiiSQg6vIByk7z
7IgRR2788WbY2xhLCOrUsutbLz5i0ky1U6lbRSwXg8krAEfojqYOVdzMlyE4acba
TSlQavyJEGg4y1a0AQC9/wHga9Gj3GuoPbg2moR+xquGYBuf5eZLt6SHS/2z7yPG
hr3i01v78cIf+VeMpvUMGjFb3nSmsIDHIElDvOLaYKh2FrtZJbkLhMHhrFSLNPlR
RdQgRK+vxCCXIK8LL/U9V8+yomwo9eHQk8yOv7DFt9GyZOtUJQq9h1qfMcavHwmG
Iu9/+iW1jgsV70GFgfFat2O8AoiDzRxTnugvIWSYLf7kcRgfBjfWlJDbyuEt+TNd
0wptZOfcfTq0q4NGu6A3+GQXy8cVnjkyduBAkhmYc+KznXHEoUKGDAjWfioEK1SR
2jRx7F4cNs3ybiGQ7X3v8xA+B83/tnfS/1GPVSAsxcN1JLY+pf/qtzCWBzqcweBu
DoBKh6TqHOS1PIk+FXGjOp1BZ4g/14F/6B6nG4iKGLuImYZoRt8Skhk2d44NhFVh
DQ1K9fJTIwz9/R/eh0wxUtF6R4nweXrcbWkBpF5IMlL2eSTIZc+LngMzac06J4dx
j9V3pROq+u5a6s8B12Mg5Q==
`pragma protect end_protected
