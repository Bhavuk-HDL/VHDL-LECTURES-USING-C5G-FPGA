// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
mE5squzkDJ9fjTko+IvlcaQzoMyPJGs8CjEka/YJ81TInOMxAul2W1J3Xy4U+wt69Fkpu//ZtLtT
MScCufChb41k71jeE5R2Ig8oKkUMNVuf2tQ7rJGuRxAFtA9V88IM1J7XjwtDgntpxrIxKw2GW9ug
gAOTU3wfxiSFXNNuJGA54X6hXC6lxDgw68D7rnfymzuAiCjAUgiKECQHJtxslEzjhwPcfp4m/8E6
KqkqGvU2bxVpXCLvieBU09S1TlH6M/4tNBGzI3T5hFaX77AWZFdQJMeKO4C9fYoNdkUWsUit/nd2
HGmet+iHEjMD46o84Htu1OEYY7+NiKqPeIzpcw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17376)
sZYHNVQfHAc5LKp+DKI3DrfCTlZedR7AhaU8mjCZXZVdca8i2+QH5aqAXUp+3R9JlUePmnADK7ii
/iWw9ks6K9KZ+Fgdv12mtdydUUcNFD/a2hfzxo61Ub1lAe/On1uUqwFkmLwvs7jtZOs851Ew4k8e
7z2ZLzUGcgZgVJMJwKtK7gXR2CSTgD42Q006kazgQGBRAzqTHouzgRZpi4I3bNs4AWk/LpZpOKG1
N9KkZQ7oM0pe/dznxwSVhN58j/0D4hCriVvDDVLqgp4qDzgl7rl9PHIGd7L+7m5YHNd6/v2uJ3fD
etBicPgi2Yg59cwQZdEyBN56zVBQPyY0ujwsNi5JV7kZgl+G/GBZmFSK4vdB2ZoUAeV9BwZ0uC3v
VBvc/I9XhhdoB+tfTuZi+u2ndWb0pb39DSoqj5bbro41QkGqYplbkeih9rP3JtxM5Kg+/R0kg57P
MULPkV9BVBUotJWy4zmsKR+KWIeVqrVb2/EHg1+V1n9YyG+pxOYvO+SEs+rgxDs6Lv8ysqKKiHtw
LMMdtJ88mtsI54YcxcIg/XhSFYEkP93BlDmzZhJGKGejFg50ppHkozRfNGQf5h9AK5hk3+Ka9l/p
i3u/UNmPl52DPYzKqWjkRuPQtl5C3FL4uB0T/5xsWJv7YDlyQ7xgsiqKJr/+kKlIsLKaHLy8Arpv
Hby3HNkwQh5xfnZtMkn93ku8sRQjz5wfnSNO3pjdPqFY0/vZh2nxQ/laIHNcxYM/rstNvn5kDelM
uNeodB/5fxll5l3xN+lcvvNJxKnks/P7V9Stb+ZDCR44RG8zttKGLStrEvgndAkjPcoB9H5x44xN
AQP4z8O7doDqNKfCW/V06FyLGAYbZH7Q2OKsefeTIHefwraFzR7IwQGOxXJSfdi/f5eTwP2iqB63
xa4Z+Gv39XEfhwi24Z4sENdA78HIv1TisN3lMo8MrCeZJa+ctl3IPYHBugQTrqtcyRXJvX62SUeE
To1VlusRK363Y1fxrYsU2sTFptOHBbKwh+DKqvov9VKBV+HNynR7MbhSRfZ66RH9oSnyzBMO7pJR
92lO7zIbyzT8hGpS4/qb7vnc0rMuXFRdsvLxAN0fmg3rshlMnbKViCO7eD81aXP3UyfwddeMxV2y
SggWo9vkR84uoSZcgKB6KSkSYnYRZJU75ToUhRzabxdYMwZX/VcQMoT28I46xpsrmsNQIfe/rN+Y
reZnIAS445VtU/GY/1geAXyPGqewreJXnT78DrYggbPhBuG4eNBlicSXoAswRslmD2iI0U55prYO
jwMZIF0O7XPLzCEGNmQtxwE1Pnu7jQiKDj8vUopGp0BiYypGHcwbCqgkkpLI55iUX/7pm5uRKx0F
b4rNMl+IHZz9K0X9UjEgsR0bJ0fobNV0fgjGpPBg1CntGemT2UcQrf6R+XOGAtuuic85FPabusAL
TS2DS+sr7PmErDYFvp2UESetZL3Sf0WBP3T9WhD+aWL3wfIRzYWPRZF4VtRCZH6iIssW/XKW0LQC
rSm+rdIaMkHqSfluEwhL/zw69psCz1+eJjg4Ceuh3qg2j+xpJ4UoAW7EQuAf0g+vv9u2p75ItTgY
C5Hgyg6oJuGGVjtYRf0FOw4108muFZqrsmzQhWxPFx/EWp9zVQxIblCPl6O2Foe4rF0m/0I5h5bh
jIHsb2FgH32cGFJkswd50evjEr8ePUwUBzym7TY+qYtC0RWqcpuspExErXtotgWU/cQmjqHqNg3a
Picd7gGzw3cRecPVqKIV+hqWCdrtULN5PYsQUzwMvHNKJcrjhvJaZhzpq7I0iAtCnBaEj4Jl8mtl
UwpHdwwJBzeqSr5yQCit4LV80HRjknzX0FZyWyvhKCWK8MsZdy4rKRZxJSQ07HdGGECg0xG7Mwl2
w79rnTNNWTtSchzWTBpptCuvoK9wGTxnQ0agAzL7KOdWc5M85ohaq6fs2Pwguwei4UrTK9fFh18U
BTPWtkmxJuFVA1uxkm0SK+FUiWc73/F4xntgf0ajk0GkX26n2tiCuk2lvLIrer9Bb79/rvvScb+g
NzWV1UB65IZ2BmUWU53VmJyX6ieibfoKOZjF7liEzgwofz7CVZtrKaG2VZhCe0QL0k6SyffNVQea
ZaGRF4+UgZOWLf0rlJH1wiMDVF8qBNMsUgZ1RBitqWLa46sorIIrpu0RrjPiI0cKTfmaCqMN4BZ5
QHjzMFddhwFVN7fzrF0J3OVdEgjQOPUGjCJCWpisVk9gHNdaqC5pcPuTBflvX+T28ndvYn9bKuCm
Gp5qKLiaB7wXBkIXYZP4vzsEamb93S7fF+SRPqbpTLqcnQkWS7SVtJ5yBMgfkf5WRxrKjGeitHr5
WJFsqPGh/mziIRXT7XqRe9yVmcxjuDv0gQMsUYbnK+K8Ymy0AlAnZ+qaHgQA+cmEMHF4yGxLPYgo
4fbzro5/z0fV0wiNm2Fqd7KVBbtV8lD3IGZVQx8Q+wiv7lgfEg5glK4uWreA0r5L1AQ9RReZR9qk
abNEpZ5L4y0uCSBs1/AXDTBQe/80uxjVtbedbHUpgGZz9m4OKZQ0Nz61sm7qwweW+24SbmhGPlmo
Lc+1oylj+gKEZHeTA5RfeKwKEUGjG6e1Ag2TFWU6DkFEUJjIgasditW/RU3AdqtYhuTM5s0BToJ9
7B1/i+8VfRnIDXecpFjCRZx+6uk/3T/37r1XLCZPEn3PniBAY3S5UemvCGE1rnmFSQydJsFucgSO
r1dtqbOegeqKm/cjLe/cTwNtP1yBO/Fsf0eZlkJtT8DjF3/WLIznUGfO3XG3dViMc8hu/zYe3g3H
E4ZMMLxvkYnVf9cUv8WFEh7m2gPl/aYSQ0+mjVVs+c7VMzV9Qn410/sU4lAMFv1FGQL9UsuQO0jc
cQ67W0g19AA7gKvfEOXY8RgVy0sOI+1StBABzdfHcxoZ+qJOMNEzNyJrJULckUeGxj34B1AITcr8
x60EesY/NOC2EWzu89GzS9Y0Rtk7WLXWd68+PJq3HG5SVmPd7dQC6K0TnZ7M5xyyjKDCl844xgOX
Ojgt78pGDxbMzbll5wUMIJa/bDaqtdFkWEtXB+bFNnX/rDo+tlLbj53TwRKyWs4/R+KjtmO3ih10
Ryri8Hn4kZN7UoUVPRA1zyIDVNIDq2RrqUKl+aQTLeJLUndSnS2o0fqPmOG2Yu/bCafpImNiubJt
Z1J91xnU4Sx70rifFWbMlem5Aw5vBHfjYMhmMtoDjU0KAT++yVGnxlXBNwPJ4/WTghpvXkXhTS+/
mI1ALG1wDnbXs+aF+8X/HPJ1HntbHRtBwz50ZgMR2jz+g32Ctc7gu7x84qzmzJZ7vcb6rbzBEbMd
xOko9t88JOlgqK+4FidEvisirt7JcC8RMyn5JnRVRCe9muZFmb7stIiw6pHyPxAqxNoqKuGdGMwf
4KxKzFisMGY2IR72yfg0SQDmW6XI5qLKndUOQYE4Zu9TFXv2eA4TTJAjJH8y2gIo8iJMDhPTkSRD
uTERlTPIVbZnGzt3oSE8y8aYesJL88pQBfWw0Km02/0J3bRh5nICcBqg+ExOGrdf4Fw1qKZ7FJUD
TeUWGpVZaV6zgZnPO+Cl63bdaB2lYFvPAFq2qJPril8wL3NSNwUsdELHbQe4wI2EHaRNmXCIPfU1
8BpQ8q1d5I7zWM9FcfSJ3sdac4F3izk2vrJ1IGnSiwn6/Gt9n/+I7nH9tzjs9jVsP4JgGOt5amAL
uS3HpcTS0vvMU2dHHkeBi2VJLBfbQMUwjCSQ8AmIbzGRFRPlIogrhNMjKfq3vY6ViP2fZA1XaA+6
VAr3UIG8jFkKfPV1cnzYGmjWlzX+YWjRAFReYCjEDlQ/aUIrJ/YUiwb8wV8qD/dViNV5t5YBLAhW
cqEwQdRaMQtRtclLBg0EK8S7+RP3gkNa/BYDIaIp3X1bU3lndvBWvrdzTy97a1NbllZVuptouVET
950IbN9ZoJkK2aYWcRRk7YrWDqpBSqDdsCJgabEUJBFD4ln2ijJFX32ji1vId4aOPNU5oREOhIoi
OGoDpsBWISSwY5F37uuhu3REl6FInGXliCkHB1Z+3JjY1xLgxvhNauv1KFIc1QuTHdUSIkNVtjdA
FzTM7c7Gw7s/inOZZHe2zJ9kNoKTNPY4uuX8Y9StIOt1C1cDH8Han7NzTVB+vPMxubonCOLt55IN
uR/LrzyS0mCf1qC62s52Ib888PcTfo95K986q5BUZoH9oE/ftYIwkv0EgEopdjsdNkknc8dQYBMA
iAa6J1cAlIoUYc66+1kAgJDUTUBTWNxauPf4PE6VohOgoxgY3adyjbqixtUjCzLLlrQOT1J2Uirv
mGlnW8e8zkxyWu3VLF81PPhNHiwYIBS5eljr4mP1+TN0kM428edxwGl/pJ7x5j25CRdapCW4Zawk
jckaFV4zXxeG3jtxpZFItOrUqtnxotqx1DO7taHJX+2z+0rFfNCyi7ktNQviYRqjDFkDjDb1NBg9
N31/mPPOz6Tg/5QyBhQfK0YKLukpifQL/ulzjmk3gFxIcDl4jpf9bEDYf+THqOR02ls/HF39ViXP
gOf6Os+Kjbk+iRx3250iA2Y+7tPQCzQxqVXczEuOhtx7rTiMlqpy/wICddRW+3x45Oq9mBK+7sey
8+bverWjTk3Cut68EmPlcCGgSXOuNyzvZk6yzuWlfROa48+AQD9i3fNDQ/3vRw41XsSL1dT8v8s/
i9yVlDLC381ozldpRTYve19QHbqNITcflQngKi7MBzf3KkQpl7EGsfrnYtsGWIHVtgqWt2+PMerm
dMsTRVYFGaehpWgc3mFHQh/W5Kigamp7pX8Y/+D+TDrN/F+KCH2JYzVnbZ8JS7nffNN2L4tsaMRU
E4+xEJSMOXLNCyeYB+lP9qsFtQPfSAEMmsjW0wWvBLhLr4NbbmMkM/RUP115PbXkarB+k/2ZjJwB
a/FS7T0yJAkZLejeBA1ilLI3oov6z6Qn+lLsPGTsrRpZA4xd4dG+l1HV7fwiTK3FojbGs6/tNAqo
bZkKkTmn0Iys26cL7GL4alEiBM71JIjo7qXJ0Bi1ILkF2T3SbeEMzz0SUvyn0e5yDsbOWDYGIfOP
321+Iu3PzJuE4LmoT9zGF/T920D5FFRfjk5E3f+PEVDptInNnEOUsID/YC1dOTrEudq5K0buQQld
QHjOaG0W/SSiY1Z8mUoeo8EVnQEzdcNxTPQ4oN4pKgYuirmjP55M3j09wW+mmlgnWtvq8IrqqIc1
n4Ba/Q4fcDM522JuD/hO97fO+jRdFSG2pQT/SA2m3gQIesSIMvTykE9iu0KW8g0DAAx++ArRmlGt
nEgwiQrfL/lU3r8RJHz06f/EmJQnRhD6Xe+ipZMz/Fe6S0Dw5o8i26id1H2RDC4jMeKUVu/+ziEF
YR/GF6uUJWUOYWMohRIirGMQ7w022oScfWtuE3JkXnh2HAQEqLAU1SsJkbln+agPpKnazv8nKjSg
hDvMpgmTAkaKtF2d6IGdU+YIcYyiRNQMn2DSU6z8FiCaGWiQmET0m+ml6/vTtOi4i6wiOeIhZg9C
kAarPNSdNb1C+4tj83bNSBboQwKRN3zmQ0TXpNGmEf5s4E9M7zAUne6gf8R+hNEMZNR/kCfGcwbP
XYvoI37XsMcjYpyTOqJnBJ6SKLmzlS1RlQ0AN3MQoZO4CBPTxiR4BBHHCtoJU/RopIDt1TPlRF3t
tsZdoPUxmhvYef52LsZRrG6pYy5r5RofdIK3Hu1T5Q8HF4zRzTB7pjOSWqdScSgCFYZ1OcR8992T
DoFJwLmQwt+9f+7CQf8NRIAw1ua/L93MeqcSfbQrV5Ubzn6C0vwnPq1uGiqJj6m1IwM6XfXh3ItE
yXwaGcx5CMMgzwQCIw9e93Qb6yXds0HYiKycIsp4V1GyqW7JAnTi2met5XKxQuUUTgxEb7SdhOTJ
hKLMP4JhSgpE1wbfEM4ITSZIgEvLpDt1Mai38YRsWk7slUH976UMzt7Bc5o04bMBktK9WvMr/2Fg
5hkWurodR5uv/+kBni9IS2nqG5TLBOCZZRBncB7Vo9kFP13nv8vLzd5FrL44trVZpON2dWazo5KM
58tUE1K6tI8u2gJ7bT4fEBuyqQ0S+zPoUj9WWHQsjgO4vUf6Gbm2/BnO4feGckoQn+oIikom1pUt
IyOljfmWQw3CW0MISye5anCbyFEltH/KfS62mxBSGuPF88Dt7yBlDU5mrSFpBtjCkZCPWuhU//gv
bTUlWBTXzc8+VPw0OedVfL3hybEyk4RHF3lzHdTtOypfLkCcGhtNXBx0d05U9S9FvE5GUarnogDL
WBFAcvhcK9bb2UNEi4ezxJb8yE7Z4QbHme4P8lxx0oOIhyupP7cYVZdn5UvLnXTKb7j2x8wfnLN8
2N59hqSb06n+mK83apEy26IPKM16BYWtVVDzFmFPbydOD4iqULVELWeE3/lEwCtPyj60KDqhj9zg
4BFzjaqiV2THW3ravLxUkgT6KBHLIXiDi61gvD0kbgHPFPF+j8VtjbMhzcrnaPGCbnZT2rVAnWVr
CHtDfobk+nui6X3fxiFNZ1I5+LbccI2XbgiQrxxlqSo6eXam2psb7EiMk+N4bUHpGXulONBHLBCD
8nIZPPw5ygIKbxvTXV1UHW343DYhI4q7j4A7RtlfMPP/sV+dlw7eRDjDXr4eY38MKlMp/3UHSJ6u
qhzpdKOy629wJcZtqIByzpJ/2VJ78ewZxLBVByaNeFdRflOFDWmdkb1/mn4WgQgdIClmJ6bva8hf
RzI5ga5b5QdArp5VPsHUC5jqeumNaS6K1od1RbTymDxuV6DailulMbuIf9JgTFRBfPlBYyzo5IyR
CKgXVDFgAAQkEG8Z6QVe2RLNSqIsLObhGzgX9JwQs8f0FGBAuO3kSX4DE6OdJ6yxwyXltT8Qj2c7
VBdpukNYuX2KpRnG9KRjStwWe8cFd321cA3SKAYTfhz8g3VRcZWG15cPvY2uPrgtxErPtjpYHTcE
MbbbPPxz0UMfo8qdtcxqIg/CSFLjTc6I1f0N2y69vFM/sGkWECKwCHczEn5Ejj8HMoPHMGLZ4wSs
T1S1mX51NYQiML0kGyzH7BZjEFjd/ozfGlUxFS4G2y/bq9ubZycemCkhnJU/SYAMHJR6ydCvLBZZ
fmFk8tWhGp4HjxGeeqBbxRL/qoquRNwnX6AmNzarXrh1r3zkuknBv/2UF55Sb+bd8G6/3UbvpRCK
O3IesAJ/wPZhhP88EXB1I8Tb2BVBMAqM+H8vYt2WsOllogB2OXsDa0b/sqt+OBlSvmytnLmHRUTN
+QBs0DSgA0XD4BCDK5Nx5R9jJGLfQfu0EcLbTjMQNqQ5EY3YrlQYy9ZrqblS0ms52sUyy+pKIbHe
lD19h5Mw63o5u2jR8MzmKID6kbWpWTgp1AOdM8tC3V3/PqNjjQqle7Vq+clZWSHpx2bnfyjU7+m3
2IY2cL5mRg844J+eISSDXlPSisQSLkdcW+V6EL/8IUejqFZS+UFYj8PduoFGQ2/L9796BN3qmXHH
0y9I1ayspmOsnns8lwS0OqsF7t/sQijsie/pKB6HFRgkV1kl33aYVSBnOZ1HpgEBfCTygcQN331z
57h79HEJ2Yrtmd5/GxLSY5GLt8lTDKdIWXnZesaM4H+tHOLMekhoB3m5U5ZzFv7J0KS0n/N800NT
w1V13Zl8FtK43Owz95u/8M/IlOedN1RndUu1bXmLwr8NBAQ84VUfapxIdna2VWf31tKv+wbP2BiR
SK8snQ4XTK+FLkHg1vtduNxbnGhtmTCNcK+8Aw+LPlxaPtWaVmCcj3TZJ445F6szCLWGEH9p9t3R
YCYLLzscNFZrguzv78VVeQEH835O45dBdUhiZ1iNAmRp03U5k04bRkw7nWSCux3nkGZB87xRr8R1
ChXumCiVVgXnzLvqxhVIPYekedGNOqK3ywT9NNezep1N7DGTascxaNqt1A1f33FGZq5fE7gWhfAK
YlE4P5CedCitWu+Nflh6TfCIumdJYVmxrZXJMlgTnRzj14LExSmd2vXe5y/Q2e4E2kTAJgrjhszT
6qJZmePU+wmu34mRUdrGAlViNldEniwbPUHpr3lnovcH9Z1QXj+N2STpRDcpjvUFQEcyTdf+8ihx
44izrukR8hWNX8Yl653L9op6ecayxRbDQVdLuwUpEXkClfWR8XGzfVVvNLjC4t61F/TdGvxmuNNy
7gin7etL1XaQhVQSVLf0B4+fuJH3FXXwjXUaR0awN/g2kX2nMFqVV4guopiaguFSY7Ln6+G2xrfD
JU9M6T90keDYc2uEvc3Bgqllm9XqBM6BiY+bnl19t1TRdo1/bR9obqdOw/Lft5rJChXa1mlyKxNT
gCzQMDyRnRgSmI1jh5OzxVogjIcZtIaJDVMu9ipnpOHFbkcYvb+LEogBhFi5jZEpzVZD8EQrxjFY
UH0ydf5DvOlauwebmZKFWPZWD2XC+mMCfVWJtV++N8yAn7SJ+E7kg6llQ0oLP896E2ii8IFs571T
MRHPU3n2HPvo8vDX2ygr6z3nqRu2Ty/Cj0MBNQZZcZ/Z9+GHJeSoCl/t6kyJxgfZCnCGF34ogfm3
pEkuIhoQ693pG9ecSbGLi7XT324tfgbpqcex4+AtGFtB3ly48HHvSqlWnlviLQgiwwbSoBw4eqTu
XNH32sTJtKQI0ULhAgbGRzoO+rGTJgUCyW4z4UTOuXfBzs1bYPIVxjNfNojON089PP75aHgxx9d8
2DIAk93vDPmJCBaV3P6WAbYUoaNJ4EHVDW3TwaY2SxO/SHvbfBh6N14Cwo+onDt+MSEcKXyS2plT
dEVXmjX5o19/XlOzp3kcZUrgHhEFjS+xYgiya8Mz4vys3q2ymxFyrHZGu31ERCXjIOEVMm7rV/ac
PoQKSTj7UCMho2XT1eevR+DpQf4mzpEGKBSv0WVEH1ffSYgBibSXI+OHHNvkHytkINy+haGLQUiz
zXZ0GfZuMZyEFChNc6bOwoAzOffLwSbu0CPJ2M3bMi69oGniUsQaL63/+U58WGv8gR68swIAyZmY
pI34NNOYOfKZHhoBDwU4GI4dpZbfi2eMgyuqmRrHsJnfvHAvWEWEgebrjHfYAormgBTv25DAPwZ6
i7sbtX6i7AuJOibMHQTg3gxatfsBgFNcAhfdgJ5yDQgsCZ7sSNyDO8l7QeCWiZA1X6SBT5fZ+qL9
eTrYPQbNtOE+hkZm4kO8n3VFjZvmykzHuLcxie+nYLcKW0jKPMeOF8j+WXkOyy4nx0uGS7RWP8LQ
aGG8gsv5U36svM+Ryqc5bhZSs6QyOfSrIJJUqCENEgdcctHDB77VPuD+QTTduU6rB97T4nrl+m8Q
1G1zY3mikyHwgPiTQX3YqHHAYCrekuSmlUs6D1KDxd23Iqb/3LDi97N5rCgXvVnA++RP5VDxWs4g
lMk9GPwkl1XWQN3r1JB2MNXq6DwFDZpPhHt3tm5k8L37/sqLBQoPwvUhBXEDiI6a7q/u+GUffwRJ
74eezCUoStenu/P7+jMMBAh4xZChLTgNhAyz6rzqR/TrRJ/0GT90Ge77+HbuQmlpKJFTKp6f1Vod
kNIByTyOfNl8tNC3tnCLLcYmXU9EuAg08Xy5uU9tDwm2cvkKqvNC01CYQNdvGJed9e5wcUf47UOs
u0ALkEA+4FzFXV4T+08seIUZcFrMRR1YL0/CxVHIfawnLa74yB+YKV3FNK4vT4p7xtVJnEBfcOCZ
0Yc6aE+V4QluR3FJsC5Hi2WkB1IdVu+FiDZ2pxPKcNVn+6+ZAqa+94m3jkjgHSztmsRjto68WBVV
SrjGTuUI7bTbK72MVO2zv+mkmKlb71wDsC7wOeji51dcNMKSDFIcIcKx1MFOOQ28HsEMYFfHZBBe
YSobTRqBWK0r+6beZiRBpq1KIFU06dIUA0gP2Jv4Eg2QrYjUwa9efQSxANNZmawtBEuiHQQ1K8M5
CIx801+liLRPPcoSDOvFEb+sp6jW1V8gSqWORt2I5OWna44/EVaGXnWloK25HqYPlszSmgY1Y6RZ
7ENX7Z5JMiD8NEj4d21vTcp+9x+X2fafU0IhKmMoIRZuXH4zw3fjjpVxLE5gCI7HpuqLqfAWkocn
i4ZEOeeq6AcxGlOmhr2qmWXXLmNDx8V/hjAIdLq6oGHdIgLdnEt0x3i3oaeKRziqUF+0MDchusnH
ZuXCOXysGC2g3hWvNyRcoyCO2ZSXC7bwpEDAufzxMDZyftlFw2M3VWthMS8Bf8YQos1WHcR5jSRP
dOkOMuS/+N44i1DOlwr7KYXPbMxg4XwcV28g/KKu3gkt2B5EHsTIfwNqYIkwpldfqByjOTPhlPja
lUXSQRsQRNGnMJxvS/70vyzv5/3fhZYTmYOJOHl/59JyRob5cY0uN65q9dz1ntIakY+KV6Ox7Sn/
BjmLrlDHspCYC+3Ss51Z/BdyDTdrkEBCyVXVUKkJSPWGddG9KGdJOHEvcGIlqd+HLY/IEGTPRGUI
PMfm1RPdGPiwvDPN5MfAnZhXa11ie8VSqZfLyj0DNwEfBDb1fXbkZn7jfXELd0cRlNYl/jtpAoBu
0gXoYP+ZjgAsfZPH2djcjL19wc3NI2tweYIju6sGcpEjAsNk+r3oemvY7IqY1aKf8yAjQOj2+JqN
GSpXlQ90z2wduBTHP1ihpCl0q2JqKvCKANFDQFKr/rbpuAeKC5SH4Dgt9Hj4nthaOy+x03uyIIrz
qzScYIXdawJYDfJVoYQf3xMHM6sz1mKHgffeWgRdMsjG8OiJMkQSe79fQ3kwFQIRMPCI5hxNSKpq
jY02nwX6loL3lT5nV+gY5+DKuEgIttd6LmqBqxqkrZAZbgaDUQwocvvKJKdiBVPjt1FmcisyQBug
R1lY9f22ll+QCgxOcoC1txRWNV/3hsKhVgQhgUm5yzNjxbHm1yPJVm+vyfA7qJLIGaErz7Y5PNJs
lwUbpjpkPtCekD09UIjrvfwBh+YSYqsE2bSnhPdMTR+J64nMVklgIMudLG3C2cAwgfGhxMuOZk/d
a/jrISrraD11IA/In4W1c2+JhZrozUKImh42yQ/2tXLnYDh9MruTpL7DqmxsBkk40xBMmBLpev7e
GX9zmxsrL6o1kXrqCWe2O9vIvwXLZDQ0EmEe53prMFO0ds68bN0s+5haE4+YHuh6PwgWRLwVn4FY
/YjJer1w+PEcFvvrWkrHkjTLStkFEzVk5gnJM0cK0M+20/Ybp/jWVPoGo/JYC+xsxQO6Gp5B3vs5
gJmM//euYIe9CKsNp8XpYyNH3akOrm/+kwuYcEmTTcP4OumMCq7fRCzhsvRB2sso/LFO9UPSdczI
aEOoWkYnMKIC9EAb0G60ehRMxRZBRIMEp9hGPzdkK5XcRCar11KerN4PS/gXvus7BOUBBQysWchH
nWG8RMaW7LGYcLRVedogSus/zc/tzRLcdD9925ZA0739920BFYwKgDowqLxR+5MC2BbK7R7ku79/
0+ed+T4NSX6XjfuoN9EZZ3AiQn7NrTBrD5Pt4PLxuatJrd1JFZiGeLyPbFHBoT7h3trkfPiZSLlP
QTK5poFjNM8kqc1xIr9xwgibH/J1Xpgms6U/CO54DSzY+X0VEKlZNvCHYbLEI4TLrAKkXtZtIsH5
AD2BviiiJLyBMnsyRQ094qCuMEiZHeorNIckIjIJMOVs5tp+kTkKAELl/kAbF9lvqJphVOUg1kxr
fjsPcDSvf5riwr0BEUaqDd/LnwIaDoqdiFFrOp1+rr9ZDVsElcC28we1CE9hbAmOnP6qolnNh2+c
gTIrWAyZVltgFU+y9UlhUUfD/Uad57YmZqafYrw+lwCqTmF2RCpmwDiipSHLpnTAqPFdtjZp234v
OgS5i5uICcLfYQeeIos58Y+MdLg6AE/s47q9PiPDRsiL4E/xqbu24zFOBg3++wnOLYmoLFbD5R1S
yEs9T0tWrzFUrKSm1Th2AkWWrD8Onuzuwz7J6GsuwkZwED8E8BlJDYG4yB5oI+IWNm2Gkd2xx4o2
eFctvuXtI1rmmb2b12Uaa7YQ0XcH8AsADAHxj58VfbRchHHy2GnIxYKsYYVdtYqiZRS0BtVv/bZ4
Je22F484eWSUVTXhYXuW30S4Y2e7t+bt9rxGjbaUzEOUd54MCvTk66CLdWgi/ScVOaRwSZ+jN/FD
/2QQFjtH9K8TwzBqlxiHmHHgTjEcCQ3ffhkJ1XeP2GPumUsEjWoS022bvUWaoI6/ZpcZnJJ02hUg
9Ew8E8SQO5MQBTfLvejdKi3RbXNR4+vy57uVNfKXOhG2oRuNDcjQ/3cIw/VEVpcHJ39xYeho0OLy
jBhUrjcjUsdOmpUZqu/y6rJECNpVTXN402A0+6aweK9W5qC7/0bkg+lPHthk4RTavck0LdWGNm/r
sOYnkK8xyl4pf8PFfGlr8Decf+eknwjQ52gDkcy7ncF93AHD+uikSZGphMhKJrKeG8XQUffDfgun
dHMjsVB5MXKqDLs7SscKQEZbYRyZZ3Hgq9rwjVhtFt6NwZ0zY5tz655BJBGXgQKmV9sJeKUy6uXv
cRMQcrMr+WzbiPHrphUCqeW8uKk46/616dJKcd3JqOmk8aurdbAZ26VxnwB1L+ssZejCAftapht2
MxeYgjijPTm9Rg2sYHTxmCj2sNqPLOoKebODCKpXsWqHv3ROibeYqveSxCQNl3VtWWD3HRf7rdKB
nsUcwSNu86JbYGBJMwYmI40XKiXq0rlQARRtPH/s6Cr1p/lJr1DpQNCrQHL6hwGTkg4AcRWvNVz1
GdVF8JETE6HsIY7nVLKqWcRWqHbTUxGUy1cFTiT+AdBNpRctezYCtkTrZpMCm1hFP+xD3Sca4zN6
1MLKxkkL4AuHvDN2QFOl2y0XPqjrAENVRkJnidrzuE5wjZZWM704Fsc0BK99dhzFRPJaqdnqh24N
ZtD3CWS6kj/QeYqhf11n1GfRYJWl7urlxm6QOuObfb9DdK2K9ld+cgH87ScVgG3JbjNRF1WuAgdn
CAlUHiszV7wYYJJT/4+8XjzBsubngc4MVPowSDIJ6XYIq+nMBzgtXMQZdHRtm9zS1USk0bOtdGdO
iottRhIMAd0xdG607Xgo329uE+LJNds05S8jHAAYcw9H5iSjduMQFn63U2AZPlq0tvzYvOKvD6VE
QVrtJSs6G2X9/+PCBcIVFtVpM6+PW4e5GX8lHh6syIUS8umOfSaHsA0efi3YB7Naeze1sr5rYmhM
UKrIT83RaCQ5aS5HSu349kAierEab0VSPfP2Z/7Gpx63tM9VP/5tc8oybQQo9v0K2vt+nVuTbrUJ
maL+oyJZB73NcG5XAuabGXbCsq5FA6Kolx/spfJ1iDX18wXnnbX71nel9uX59iFBI/H+1wE/wYqo
mcdyfxzlqrOxvLcRCEIdy9fW8TE8dRsuug/8nt9te4ZJ6Fft4Y7BUSrnPGBzYgKDFUFucweKCm2m
3lr48i7HCLBwdzsEg2RyQv+CFbJeNLsqdLxhunvAuxnCB093IofHTzdhVhWLOzm5D4gTsoDPQFHg
NSsRopCDhwL4XBHRbGiWPc7hQi/hBM+EXrcfg43W/ZQn7GyEBtitB0VHN2sUaYsJOP39ZrQe3jia
U8/mpBwq0WTnYZa9ThJPzlpswYNnIQIktt/I9b+DMykwDz3qCfBcqep/9qC83DSlj3yrdCgfxyMx
E6kc5iyGoCSiyM93AuzoDvnnRQIFhcQJOZNnV1+48NqB6UOtcPvyuzt7t+oE9hfvsoXj+VX3Yg3a
lzwBmNep6K6Q61PCIhexRYX1oC7D2QcYvs8ETqF1VhD0LAbMSs7e1cXqrRRNjK003PYXGImkeZBg
210JrrFluwXwt329i7gqxHQmdxP1Hax0zlou2S4wkxIvgnhJ0AdSWpYxgfhieBHXTqkEGzatZM/g
u4s1NaFKcztYHA0FLqX81VK7POftnBhi3Yb9m9xAMNLs4tWhvtrttI0a/5QblPFkWwJfGEf8geEn
XTC4gH4VYP0OmSmzUnR6wEYr9qoWrkx3gqwORiAfZUyEbhNk+t/6IdfT09chD+3ogbZ/NOEAUZD1
VsFdQEVKU4CcKTg2WnSYkhgy4EQ4zGpUuJaQycYZT1wIHDMbuiCCQUiBQFYsUFTmtb/9dAqmQrq5
aR8r0p0J0TxW7/kNMS+8rfJgahjNSigB/7bUl7rEiQZYv2zeF8eRc68zrVo21yMy/CCRqeyYN/9C
U1cmyaD2Ev7yTFJOE+dQS2LUsC1VYhbJF06gbnoLafzuBLVo+WZTmr+OvqHoWlFBfyrsIbqukGch
dJGRNA71cpzeDJrpaC1EGN3JRlfmjnsggn1Pl6MlwvsrLXdjcwFLkUibCcJnjDEX/rB371fx4Ld5
gl156PgxnYx1VFpIs68K39wF5byZuP2MoLsXLB5S46w6WTQEAHOZue8asUorXfK2Vt9h3JFV+PZ0
/vrIi/2SH2QEi2LwOKaAdZjM/LE2Sr9WOb4pnqefGUBUO/0I5L1+bKYITSwdWVHAJwfYbcH8nyRa
pAs7YMw0IIaDuY/xUV4LnA03bcm5rZzjq8Bzsud58MB/Uq76YtcwCVzo9O41nBdgdNmkdzNoDmDp
n9HMDbktJnLGvzZnIdYl+NlPWHuxBuzNg8tskFFqi0CQC9ogoVGhxvItlcxUoqXrhyEjS+fOMJS3
w/oLiOpRoUQ0hw25FhqHO+YWTt3HqIvQt7Cl4idy7FJBjdIvWdghHL4AofnO6VRsuWHjgFT19k6n
jRTwsQLqX7AKeIO+Kkjk2SRtYmTOU7+4Nz0DLPvsdx3L1OooF0meY7oxa0aP4z8YNf+FRMQ1stsp
jlNHRnBULcC2UO06G1unuirC2WNHkbks4T9AcjPH6CSf5yHBvtf83fArBL8jkEu195rfIrBw0hnB
F89JfhKJ2t52kaPXqV7pyshC4Rg1icaZr6oFyX3OtsfDjLdZvKkT3+kWQpxjYbL4XpxFFFzqlBCT
CzxkCCtB7T/L5U2HBrdbXPz3rYkar1syrzQv9E5K2Pf3hgWw+D1IVji4NGWSppZkBv7URyjWnNre
uPv1z8hli5dXoyuNvg6KTyMW8/m/CEhsjFvfy0edYV+qPPueAdTJTSvX8HLJ1nrtUSHaSkZYmx7u
Vh6ze3w0N8KI/ovnwqaVuGhbkMNsfDHugv4atwRFFGkS5Laiv+esZ4trI7pUcC7oBD5ZfzhCVQ8x
XbU9+NpwDRWJzqPzjGDF0IusUfLvH+KHVf1OGZQ0Oum7ngER9jzQmEQs3ZeJ5S3B7rAWN8XTIcWc
tKI0alpIr35mF73Ap+Z3yZX1k57oOFQRnAgmD5SvmeBJIEDweWpYY0yA2mqGsrPz9/dZoDMrjyZ8
5lbePAL6gKWYITAz1OX0/xU9OczO9vP87sZR7hu+m0/0bqargS7mBWWRLRuaMxM+jY0xXWEix8eo
ak54SeSqN9RdHWnnU9Ab/4xtFdy+z6NvUzgZlimurn+cfEb9zVqWM2QpaDrE0bjyinOh1AASK0P2
Qjsal3JlJSNysDzWUBKm/ombu0f1KhK+Dhi+0LMfTcRRDgpIqkm+9UQAiYp5Vi6E6C98/qus5M9D
5ZYz+My4HTCR4akMyvwxnjQbtKOXZCGwCNNYqAvhCITRxH1ZL1/gdR53+Y6d8OOhooWwlwSq1xag
wYQcacU10EXJlECgneDctb1ye9LOpGODeDb7c1mu8ptrLUuqIfvzUPOjdZV56GM+/tNugrxY3jeY
DsOB+gNENP/re+X0os8fDqfXqFPMT7R9yYhPVzDb6sEYS5DqtbWRiQKmJhMpZnMPebA1hkgvdB4Y
11uDBTnHF8CGObZqjOGLCGJc9hffv/YlVBOi0r96jAC2hqsq2TobjgUZDKNwM+2L+1ogdIZMg1s7
PZNAzkCfJkYIbT8vWBAC21dQJI7CbXDGYfOQDQPCC6dQeXEMgjloNDC1S4xqQGErZi6Guk+d00RQ
cEaHD+jTbfmOysCHRFFRdmkbKvwBMKVxpAzxfZS0QitqadQ4cGkkXXVBTf58HXLwzNkFmEU+RV3l
r5hu9/7kfC7jRcosQRICKn6OE11oof7ZASv3XQyIkHaHw8Zezm4K2q7tki06n2hDzXuqsEoBZdr5
HCUbPPSzUKYLmylmlkPDqPlqPfIszC3IGxKbnZVlv/9Z/mogcYFduMeHgvLFi1tjeKbdos/XXG0s
agySCD1MmSHUnGV9XiHFLu/ApyaknFUGQca4VXeubXPEV8oJ7nkOHJ2uupL+JjUusnhvUuTyH2iH
E1WLVs/T8EKbjCdZdUYGNn+lRpFq3kfZe0JFGcwLjlB2RX5Ri4qydBE6SPCSAvVpfmaU8oEzYCvj
OJpM8aIBhJBWhNSwRGDNOBilpntqcCBtJG8pZPvK0cc5i35z3n8NnFPC9goZCJpUCQvr2orcAuvE
auVE0GB1ysqv2nWPt9+DGDzXpSVsieH/y6ib9sUxXC6Tfcvd/Ap6gSmwWOC6vfUHP2P6T6d8Qw9k
9fOPkkevaW3Atp4RZlmNghjZTz6+aSOoZ5ybboVceS8j4gkTYNyCnb7G4MiA9M1+4RO0IVLX4TI4
rl1lj/bu2pB9v5iumse1eDB2qvfnCIadR/EAjc2hUIS+wXEtvfWVSGy6/p5xrAYD+UpBGbqGYbl0
ekyDxQXBAxNg+uwaWtdz2GnQUvfOdPVsUK21SHnEgmb8FUQdXUP9yKCjuvY4Tp+o6T1MGNFAMykD
BSOsoRmos2/0o7uzz/2f3PTX9Se+s1eeaNQiz6M81zrS2pBXN6WLA8OeqRYlp4Bo1yWupVHVbcbr
fw8RMYtWcBcyj1wkoPtpcqrCZYrJxZcPcHq3CaGmT+AHSeEWHhnZB26TLqQgF/0v4RbURrfkyjJL
WjdBBvZ1eCOurrN2rlpdlVo4+dHk3tr8poC1PIM6pNSAatZu9cYa2nKsFhzvr8htkPJChyFbfhwH
VD/XQq0bccee1RSlhMZFKj3R43P4PUCTJ46C8h4qSsbDLyTPN94fLpyvRHIne2Vil3ZHJTCxCnGm
r8tLE1EJauaNW6cEcjW5OwVPCAlONOCzWxR/A4iDm8dPMxyi9QXN0mEtn1++6v+6lKQbvxmBmY0H
wcT4Q/tuiq33r/lSLjGu4Y3ilN3HV5dWuxGPDwdAhsEFOMrU7UB/DpZR6NIlgkNF7bocdDEevEsw
KzJhc3PPoGQhKncRC4ft/H14K7MoSiNJBy5ADmuYyhzPvOVUOxHKBW+8A6T+McbJfAt8uLfTV0Zr
GoxJgAyumSWFt7EU1T+xMJwQAGm4oxOsmnGaSC9WAhH6g8/hevUrWpA1FpH70h4+ErLqfbFXS7EW
MFeOeCa6tvifuXqLSZCpDJtfQmXAE1Nqya0gmw0Huswb2zYHLz34OCAA80VeHKHt+McIxDNXmF8M
1ru2u+FpW882PSW8cf55dwwyGl9bn+PU4TVCmPDrfh3gfrELVfV4vQi9s7gqpYUem6YL7ncDd3dq
2+8xSEMIVheUByo7AhJPWiMnZmn4ZS+bWsQw0CmGk9tiy+j9ePWzjZhpOOCpSeYyCClWQxh9RhfZ
LnHLdA/RS2zQZxpTPj/IaRjvLuZXqestnWOoJ4jKbtEU+uTjW/IX4lRFXXnQ054dJ7aOToXGiK9k
diLca5KKedZAxDtLCtxcxlrZNMeqJwDNNp19okxjTX3prD+KN4IKaQYCCrPXaG8rsZzR3A0Y2dcN
Q+TCI8CR+bXOUVBE9OQZUyU+aiRs1m2npUFLDGE3HuhFnXEPcWyNwHt7bYyrXIt1Kzf4j25SjhuT
QiVdM1guV6f7cffGDGsQUErvq9eepYjJoP40/ZNfDg+7Yd5jPIuYe0Tjz+DrFWkIQdiOLSrwiK6Q
/vMIfRNrtEGd4lJ7q+QkyU6EJRFr0alap8ADvS4WY0kMirfPtA4FoK/Jd5+LBxYGr8TaBdwyjiOl
PV5FjuuSwigXpDHBAGRRmK3tH0axt7rfN8tl2RZYUCVG0UhGiMhuXA/6PqGobC1yHi1/g1+RIT3S
6j9uSIvQkwjEvL89kuCJNTtKa3bD9DetJVceC25QIzBI/+piPmqXuZt08ceCEziLUXxji5WPzPwb
NB/hUXxlwy/+TQYB4CuW7me8mWD7Vsnl79gAqAaq7z0dDS3PbM8TVeA7Ul72JX5K0/tqVdOMXHUE
lAsVpofQKTJMi48LafoyGfyLw1i1BVIaMIgqutGZVxEF+Lu/tU7jrs5UBmGY03g+uV42WXpCQAkB
6FD6pT8ltKuuDE613hFm4lkzmbM26603803TTB1sPUeTu3PpfVYvuMRdekc6kUGlcWeNOaW18MRc
FKgKNHJg7HqoeBtLo4gA5SEw3XfKfbazxdWN7u1+jJW0ulkb+UAbUTQ/Hxx3n+HmW5D+Cgye+fki
qHNrvZMhNBz+2cJYTzFybntiGtj9oSNtjS9YJb/quOEojxlqoJDPiAdsUpqtYmTInKfbWOofVvW7
um6FD1TuHmbx35gMcGZ6gSQrrUKEemTgPPzqs9voebZHtEs9RSpxF+3M17HwrMcs8pkyl7nE7uN6
/Vt4Kv+k1Zz5xxFua1re2l8axUb0si6mVWm6EGBAbGcuwzKZldiV6MS5nVB0LVyGfrZ22pEaZpFT
7DvZe1B+CqdvPkpuKs758eAzD3y6bDncaLsLH+EB72DeTWdCroHZLq6DSoDTmLRWhbrfiyUGQnS5
UFbAkm9Si6ZAV7KF0zoauFp6lRCgO7PK/MPQ25bH+MyATTYAb9xj865bW7FOuTDyYjKRT7YNcdlT
R5/CQy+UbOsa/EgUOeaZ+PxOcDCVFWgHXiaE1o38aTrlmCBFyPv12ePUpBfENdDlx7olOEXpEpul
hWjwVp7LJEZIDyE6sqEAFibGe6sY7QU9uSTY8RGDVQkALCg02mAPgy1b2RhXQKRdOWGJc2uznY9q
nFN6aIBm6PF1ANmOYnoQtVYsJBvuO0CMHXywoA8YwgOI+w3HC3e93dGS5Z66LT2q1i+OPVr57Zm6
PAP8LuhcvnWQmYVw10ggSceqd6SzY1sCxP5iTyt9DMPjUC84st8Wb64UM9Vxj4C6zxLLvhu+mvTd
WVVfflEQai9hIiYscN3M4VicVIt5pu2LgX1dXjVmIGJ27VyhDac9AtKvNShsTbB/P/9sY4lnTODt
Lhw8hwkkFe29B+vr/+liroRi8GPHf/ja0QGs8lIcGXcWEfSBMPdI7UTGRTSolq42tBa9jRjNiwVe
jIQ/3nRb6p4K8SVVDv0W1fif+IEqthRcOwaigGCiuWLbI52nih7EgM8sWt6ff3ExEbHMpPA+XiXt
qPZ1jdXTrmJFii7dq+jc+GOt+TKFjL0bgmY1pjg5J9nEsZqnNv+LK7mfgRmgnEgnSo/MHtRxLysv
w8YUtB/aWrSLN5NwZAwOR8sRu6h3UV9okZ2zu7eTmCRZh/UZcQDIHeK8pLfu321eW6ZiZAitYokH
7ZHyR8M8fRRnEYv//9oHIDFrEiOwRcs2sVNOLcS8FRQWmjy1IcMEdjPU2rGXShu8JeWZNzMmtQoX
qcro4kRZIg2XnxM6wfkKEfcFSen3p3Yn9wb3KW3zyow2+6XSSU9CHG+jo/18usVV9QfMj52SVRJm
VAcG/12BZA+DQIGjbNrJGzT3Ub+Vqzf5nREetdNnOBoBNwKHv55/kXxONIEbVoFl4ubxuMOvRxgd
Uk4HElgjtPfq9EwSpeGjnllrzymtZbD9845nPmNd8u/z4dTqOqytnFaZeEei/xEA4HDptoulFf6+
3G+aNPpGRWdqX4CIsoQTd4LewVI5bu2D/1RB/QGcqYs6In424h5LgnESCeZ8U3MXNfZusgVixGzT
ZV1FHKCJUTbl0+YBPUJeDEwSZzWnS7Hai1Lbr39hs//94XVL5Xsl/Q0+HBBuo2/yqC9xymthBz68
UTJut0Y8pBS/pb3Td5Md8W1DEI8fXLzKI3naLAfqwXUq8Mw1kLPWRDvsYw1q6IcRfheIhdCnqgDl
UvZF4IzmQLym5E3+zIsAg5x/BA/t6rJ2/ZrT7iDaJsXVqoryBT5yTF5aRo/0CgUacrZdXs2+DpmT
kB3qSL2CkE494XqABVEMPdgVL4nKZTlmTU2FBwJHn/1iJqCnBFZ/7vXhlEHv9AEHVvBUfye7wV9w
aTyo5S1UwHt9wnVxr64ETKJ2R70ezGDr3IQMqWFUKlMwChIYHWzsCD7T+B+uxgSYe5Gldts4jb4Y
fuono+jRr1HfuU//QiEIw9eZ1dZ7a5iB4kW5C95vUtpCKyoX02brhTJt/nMFPLXGupYbkvsjxCcf
mE5iwXOMq+yVKs4iEBfAv8j8BW8PF7UT7ygRyEQtuEcMnxYwL6gVmBgoJWMvYK+O1i5CDYT1egYd
gJ/lcNygHSlBVWVqYNSERtEpe74ZI5McDoieyMlobEa5qte1VLXFnggzCKQUn6oWdsuA1nPhAWL3
ug9GXfsLcSgwMfX0pgmQe/izp1HIKOC00t0vjJxkc4EDFrVii7CK5U5ORu8dVAtkYimYGNu7qZEe
ZXyQkBX06mw6wBGeQH0ZWuDOPJnrlCrszmp5kfpI9tHkXv44S/BInuCS0cG1rl/iHuvv7Avd/tLo
zbjpAJ5XfbEnYZ9s6KRHHw2+xX8/vMxDDsQoM10ywo8kKuPS6cLyUjFmzsLYbi7rg3U/0rI5LVKV
IlSLIBfi/MQdbhMnXmiUWMtwXnrvBYqHekKRNon0d6kf/oSab4dA80G29x3ujaX2npZPZ6ABOpDZ
95tsRdZjga6rqt11jV4Y2Sg3MvCq1QY3zmwkbZprdfu5d5gZBlGk4CZsjWVhxW9zKcFuU9jdi7Vh
Z4je9pOO6XxmSDtw9kn7qi4iyx1dDqkbza5x9n7wcFQymLM6cglS4LDLylUOJY0Jzvz8CqclO0Ai
yrT01+ZwamF6Xvb1OGk8NRjjmiu6dmkpfVgqw8bN3f4qAopluioPeGfRmo7EI0PivRvhPfuaUag7
vr+qW5x4iN6L253L7MFFe0Fk1oo9bBJUbAagTVmgIkXt7+9s1UYBRdwI+gn+LhDG114cya8NLGhw
2k5eA8UfGw9j6qWe1usEfzZoiiMDykB2Rrz63ML2EY+pnodTXqHvINT3/vIvhpw09GbV2qeu7BfE
tNugF78XWwfKUhwwvWJ4Qlz1U9F+2R0DK+NwZDEfJBqcuBMd3D1/udLSXtTDrYT5gDsNB3mzeaVu
fnj6a9ma/sNZucn44r2XQR3qrYNo9c6deNtb7lu3kb2bmsfbIpiw0fg/hITGhNzqogKs0x53bIN+
unJkW6wcFwDJTJgkCLI4IfGMtYHSv15OFsMUb56yTjw0nfUtex5bzsl7+3wbSR9N7Unpp3hpco5/
JMmrUqHrdLuHZC97eeZA8DxhIY67sGCQLBbQ9qE7qwVJ280mUbNT5GYtLgRRQNBq8RzWOUZF2ZKB
yffyOOOu2hxAXnbU5Qc+Xv74vuP8dwnEFXNLkr/buiqzD6nShjUGVmNo3FPlbjRQGXS63V0Z5Pfs
VN88OSsVZVO8p2QF8EQqMs50ojouBXIg77tW+SIpkLHL0JhD5sEtyA5Pu2LBDz9ujTqs+ofsmKPr
1yGUQMaFhcuxFXvbd+yGzOuNBclNyWDDf3LbtxOzQ/w8yFLo/7LtxXPctGLomfV3DFZSmstCUrHV
76r9AInrYVi6lEK8nkViJqSEOBD0FNTqQ2hEak+6fL0LYszjx+JVKHQWx5fPnAzSrtnMy1dgygZo
GE1IRoqorqlXCtWuxsiPRKm+lxOcTALieBiH8MteAMo+aN0EeNtYoTYXiXi16rE5EdGeTjeAm65G
zAx3T1I989jsAL3p4NYn7tXqapIfxXMBtVFZiH9SSJfDRdLcazYBlWq0egYUNrRNQZIowA/c2cp0
rUZX+BQd1eg0ouHXQPfK4xTmHMvwLKM+Sp0Hn+mFeTCBcoYmzUe9XKP3PnNMnZPY/l6RTJUkXohK
fnk+nGZND9SWFImBhnHenZqbUABiY24VS8zsHWYRbcB0wzGYAUM+xforu3hwZq+FXvVU+N6Wwfea
SjI1McK2tiF/KO+NqpjZAD4wEAzTaNdKcVycD2m+z3/lfvFaoxU3UuiePD+zDUWKqicpAiY3u7dt
JhqYaURUSiCvMdl6IkS6m0h1U4nRoHM/u/+vpVjr0gBuPIhF6zMljHgsdtICbGnXSillEqxtFI9B
383t1B/ANxmQJ/GVzbBVxs3u5ECq5tDnoTYwwgvJqJv0NCBeXip+xaMi2GB71mIPzVbyItW56NDp
42NXBAkthUP/6KYckOgOFiteeim8qrukroybr6j1KleuqQCamGgNbv8It9TFUqG9uocHX1BoUZ4Q
HSJ2TJn7zsbHa5FQB5SwyI0SE1YJe//J78QJ6nZfYagPmP+DIcCfSfSUCN/ou8JugJywSQiCVGA6
LTslSEdh1tfst03+x+Y3pSTvwb4H2ZUnMRLf4Ri/XambV9LXV2hb854P6TyMtXQ+abe4WZshM2uR
kmv/zBt1KxSaYjlktVnrXj5CSfwjsDTqSOp/PfisMHgLbCDdJn4nTqIJs4RpWDvPTiHnM4Vu3KsO
JB/bx5kzPCfhN0es/EeWfGAn9fakpKWm5+ye7kiw+LFuZjzETKNM/9icihyt2FmL3+1wWXwuCe1p
uZDczWyh5kfOEZgvUcyn6qHPxZMvoHXryHwWny3sswnxgWnTDWrlfY/rOcYQFTZRDqC/ooQ/S/o6
/ha7UUR2vixb0uqyksOIx7U7p1HotF19hfFk7pOeKqeA/+18GpoDsZWeVFK4KpiGTpeEkn60pJkt
RamEzQ8WsdkEwbJdKCaa79YxFbENbIunkTd3wlOGn+8jhmf+GxbX+pOyIcpYgstHK6WOr9qRS8iJ
BWHbpQrrK/HuNBp3ow/qznPLT63LgZlBF1O6ch3JWfBlixyC5X48RwRjzspl3nhh+52AuTr97QeH
oKxCsiUU4nhcio4f2rJv/3wjiPepIp7a3zNha7hZCgFksTSHKW9w296DWAevmjEmvL5GOepk7hU6
rowfZNw1cSIEsGJlnRJi6PDlGmpNKY4CuFLA/raCZHZWpd4mOTG1bK6fMIAVWMC4UMEengSf8+9T
ievGEi2jvFHZ9ytvaeVWomp0EW8AjrGgLRFseltkO+1NRIjDVbn3s9+0x3OAGuYt
`pragma protect end_protected
