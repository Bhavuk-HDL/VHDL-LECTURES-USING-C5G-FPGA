// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:21:31 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
c+7h32+p8kar0tLQO24HBTcVjxxOgO83E6HB7M/YMjxd5gtR2yum4sSjCZnLJreU
1qmPtH6ATHV12j0XeLX6DktNgGxjqOgpeSgSw8sQOHKl6AvRhDOWWn16EIqynuDC
POCRX2c44f3tsV6c31TKUaNwo8SdkDGNWWTmexeyhdo=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7552)
PkST4eUyo0omB5tiyLWxDy870m4RpsaWf2mYwECd0Ozy29Vh1JocEECGez4+gjO5
7011BR3xlDOdfuhHL1LlaX9uNAYHcpCUn5MFU/0ScDfEo93w9mJgFr9bPudsc1I1
1cDQt8VJtSn3Tz7wi+vKYD1OSRxMSCLSNhDHB0BS63GhVGsviPCJoBuYTmTx4THM
eG9HoF7XEA4f4Ya4+53VxojOo9/RtOWUjTu42QkWrt5gAsPXkElcZL2j54k2BanE
dOdDCpRJAKVSS9pR6J2XSy79f5hgXUrYtsalS2I6UGrXEk4nMiWCLwlu4gULzVCY
Al5rbY71FqMBdgmMnjKXBfQVB6Byk8QPixOFlzH17kHzxnuO1GbpjYEDQcr0nbgo
uRTg8QWrBgd11cur3dF1hfr4gEvQo+ByrYBhna5riHjykWBth3/YRHiTJAyvLTyd
4WqaWXjBHmOYeLqky9gmAbDVVwIVF/jnmTTt/+MrSJFra/LH+/HAF1QKUUCaMKSt
JS7gCqfOsW5Yecd2GVVpSoKWLfIA2r3JLtvwVUlB6fo7lxcDIJMoCUaxuc2i8ksE
jhZ7QpFJqqUOBkV2KiO7Qp+EOES+aFALtDRR+HPme+sHR5nji3pO1i/QG9W3LQaR
0NxmKWoW9K5zfx4ik8c+wYoHTVMXA56G4EKw7CQkcYBBa2D+qNK146GahQeXAz68
vsHVU1EG9wQcFUvA46z0omXewc5Lc/eak14eg6xA/hRzDX650dt0OIl5GqUlH9bf
sEbNakGlGSw93tzZCq2b4iB87ZTaOiZt+bG5wPNupdSFOX6BtP4gygwjJH595H+B
/+ZyFvUdp3w4zZ56YzK31kX5CRxFXoLAYYE7tiQs3ycK1ZoFkHf9KODn9dGreiVt
8c0g4bftE5PISbPfr3jGeR8bsa8g0MPJ7rRa90CsqHjX/2X0RZWDam7IoF4ra8Z3
a8GcuSBLnBhztsmqdiHJfidCyRzRjVWH4p4lPntDX2UmiHXWPAiV27qXDuqkZTts
0+pXYbc5UKEfJVFZP5XBk90B4TLr2MzEOkP99T4RY/I+j26kfUoRPVg4GRwsOe52
WuuKICFw//7JRxj/CpGwgG8BSASya/kxaBe/v659ImaI0uAZXLTWVF2AccVoCsys
V087lGyMXcrsJFqkLDyoOX0/gjqL7EJDrtnYmo8vKaHiPvIoCLXPrjJv/gs44DWB
q36LnTfDPFjsb+cKuXrUGZhJkZJZW8dWroieqSatd2C5iomoLWcgLeSEF9wKdcNw
md2nPWzf5Yl02FerBn8h0kehfRF5cxU2vpDURhZ3s5G87ndCCj2B59PjlhDn/hyU
LNkJZdJLkflIDrZFeylcnEe5Pz3zbo11v6H2Hir1qyWn2zW0Z+6W57X3D05DT2RE
jLA+qSu67mJihsRTbheCtqN0N0c+bIPbk2Jq5olMTLiFLtYU9bnUHeFiV5XzfXgv
cPFiNIKxeXfFKp130GCyFntGNH+L0gNm3H70ZNMs9ouPwOdDACB8hMXqv9+3Et+z
5Dx23WzSojDRKWjpovBkikYmok/nq50Sc0yoSl3Qx3UGp/dCid97aFc7oeDyqcB3
sXWo9i463fnQo/hybL0txwKQGGup5RtJfMsDvp6mWYtJDeHB87gJLUkW8NbhwkMb
ndVs7faZuMjtXqzzUKoal0128S+nD4lEwyggQZ/lm7FpzZ8mjt5mZiD22GdA0xDn
oepNqaUzjOe45Odo3vXEELwiNLhn5TAZDj6V8Iropjn1gurAUDU0v9GYlsOOr+iZ
8fc/6C2D+havyXi5/ozpFW3yu0qxWN99DPyEfWyfJvmY8BqZZ0J+mgLrgl5mHwaU
IRpUlaPDIVnt6pGXPF9GIU+HYqYpbRGgN6VD4k6RC8nfqTVbtFsJST2+qahqpmMh
rpIlTl0VyG9noiamNvUfojT5CX1HoNkh3yS+cUg9K6o3VtI3/USveKUKL6Vp6Si6
QkA5P1avh3mCT4wzKTmBxZKfovMlwlPWDSkJhsa3bSuOnMkqPy3eRU5sz88pq99P
nOyewO1MYkt53VO1YUPqP1rzDcovLfunXjtnByxj5CdjcKQddGrvZ3cXWb7uNJ3q
zHAuQgVyA1CEkc7+ukKCfNKIbR6VSXmo6BKuOhYNog+iTB/8s5aarh9XoLGRFNQ8
F54vizx5Bcr1zeFoz4Y/UD1i77TsiWe4WHNR7XptkelLUWMaurzyWJEsmw9ZBqTs
U+jRnhwBiDTkGrK8wcrVot4oYb3VyafWmaiZF2ohL58GyGe2/xY1CDpyqB+XQuvM
znWfYzM1z+MsCgttWIOE0ObA+/DHnPCsQ+fW2HMYGnEEN64vu+eMpRdDWAjSO4n+
r77M7Xg7VBtY+Z2JhB1d/L3Vy595BblEDXLsZE1IOQR+/b0AFacwN1iPMDo1CgHr
JDjETFVFPZj1fBrfMOpqMfpE1OxZKrgWBW9Q8qapMfYWx5Y88GQR+4i72wOKLlJg
N+uutSK25gO9tD4e8WANM973ez7hP9sH9xgDzmqR1jH+ZysqZpo/V+G0KbBv/NFI
/ZdAkN7ah6d3OXd0sw9FGdyRkeeKMLFhaHgD6PQjiq4W5CrAjleX8tgCMEHKsle3
ra60YiCdj9CcxBu9Uz03PHDdl7DTED3xL8WbQbutT5o9AosZwWoV3Sic/3KP54T4
2pA8yUQP2uAF4qwxn85KYOYdpMd20wn5gNV8oo8Rc1lPVR6v9df/qLhRAn9Eqt07
3lQ6z+Gy4ix4UlMKx5buncrvvjp7DVWH/IDhtHCZBfOagOmnEvW5/4zijOAfWX/3
0GuLbWHQFKX/lHwlRfcTBcuYTgJdi7VxF0mOeX5c5dtQc/8IYrh/2kXt7Pm91zUF
6EzneTXQnrxP7uQjRDVGhwjPLK9TwcFCEWZs15JGtYS1/zHytojRyBnfDve+ce0C
Md6HrqQUW231AzrKgWtbmEJ3KzbYiTsdDBsDGnRfCI05nb1o+VjYE6cT0uegwyyu
NfqwnMddbKQbHW+JboIvqVjvdZzTutgXMudaJUbxBt+mRyIEvTBZi44Eaj1ei2SX
fZm/5PvJfH0mOEyBJYvmFsPgRuBVCoVmCmeZJjQvQ1kUC4Z1ErId+N9hS4q4Q+f8
Vt8fZarQhtBCaLrzBWvSRHyrGjcHVBnH55SvAEqzAUGukFr9wvxF31B/QponT7UB
XRJSPA2TjJvjfNbah/rHHgYAouQrHAJS7xpNIIPAuQUhfnD7UFD4xlZCXNI9FbA3
xMQtdEGALJuWeHBw15/xd1AGYIO/2qMZelsNYb3+PZ/pdLNK0yrGGlqzqT1lSnNa
oXJRfYZMW8svB3L002znk4/z71D8z5dk0x1KZ/V0bSYtpdLB2Yc6GOZK0NxGVAKr
gUjF3mDb2R00LHsJdNKd5Kc+K7Ea326+Pn2610MJoixlR9fg/qxZUoXbUifEBgk6
ML5fLaW7eh9SPtS5wdHriiorf/vmX9UzNXPijwLIPYAuZZepgDAE4VUKna+kHmxx
hcDudhAiUMmP1JPiDfI8ePrGqV94lVYv6I8py9KgDJbjClFJ30v2Y7r/lTDox09c
M/V+07HgKjIhHnVkTNZrjGQ1FDWtS6Xsy+kCsOX2MW2CWoCwIj2foG84vfSmoOpG
OiRCGndRSSTX/+g4knEo+WlkNfOJOfGEU3Ua7xbWZAiM/PAzv+7r9kDlU7d6op3P
Bq7T75b0qplUsKaqF2ws1Uzd1o27Ct7kF99x4wcbUFuqKlDrt/nlFZwIeIJ7e3tM
7TRU/4AS7P+Vss3iC9XcsWbK34QsuTfRqApFNpvLCLsNkgwFiaUS3gLt4a4vya7F
YDr/DM7HUjYwfDNlJSIdih/vmkcld+dAZuFUeBSAHaR1pMoG0dekoqxc4au4zSYi
XYwoLvwuihTXWFSadfbmAP1EtdqoLGsbrvYY0bU5LKQK7zvzJQSe7gAh1W7wMYIE
AIEAGaHygXJ6I/JB5Sq7KBEL3PzHJn133gQnQWnXRs+7QFVx2E3yTTkwJJwDpXUh
+R5UhA0brJz3pZbVpV6ApLwig9OoTPhZoF3gZ+OnwXNYKd00kt6g0WwNUNJ9arSW
0xx3azvETeAoxMFrFUF9H8lcZs4hbsJQgRXEkUsgG7U4twCEPbd32aJkMZrwLNMU
wabOUik+oYbLFH1U68H4jC3SBVccBZ8sq4L3zTIDLtCeGm5IalyAhoTvfJFJBsn/
hqARs5MPgLkciD1y9jUwSPlIPmlSFT5EEjg2u/81BUrX+ZP8coEH8ENIz3z+wCJq
nwSSCXkppVw0plQiZh4B0dUWvucZcGnc+YqqVNHGdTWRz4nMkD9jxcB4OdO1IivF
BBRH4TWdIa/3+d7oGvOn4JVVyzTQzbC/2bapuQE00+TFas2TQASmjYTO+sKqe1Hl
B1wU2GaD0NKnAQAX5BcimrK6gEKPTzEmjh/j9ev/NMTTV3yUGd65Q2OXEp1+s6+b
vA7T6eEl4qizxRI+qVQFBVMzFoZ2QYZ5t4xhBjJPK9CKqA54vZWhzBWN+TgelTBS
dDnBFV2pAgK9QMw6UTVvyl1w6rrm7ktkvivc7iLji+6syNbhiObCfjP0mWF742mX
Xtfe2aLosAwNgERLdA/4uBFbpPcG9gcaQt2Osz8HNHBekSVHr1KIJTsDRb9pAOEN
PHi+upolOsd59WOHfXCC2RYN88djQKih1l1XGdZVYCaV+KHc0z/ZcAcdY3Xpelb3
tb/9vggo++RggW5ExFeCocvxa/h9yKXWUlMCq0+ZNonnSYT8KGtxroJdJUeXNJmq
I5mXWOTVYc1vi3mZhnGv2MqxMroYTKT1Tq6pGuC1PJvWZ1qPRyJjVnW11yjn1mRh
iNYwR91VQK353L2f5ZmRL+JvadNthkguQpogXQ88xTRpTPpKzL0YS5WhxjZDyEdZ
5jSdNIj2+uoTyv08undDr0bWOlwI/1Oy1GpkRHoAqEZnSWyUIq36Wuqve/k4CUnv
eIgt3XKDa3RDJ+C7qGpleA0lFNSjRUND9vXVX5Rzmy6jswx21HW4skwaYJP0qWQX
GVD1ndZjYS6fnGwHbWd79BvZCkphI+y3UcDAayi8EW1vbhc6OdNXEz9eTxSMxc7k
mZfmV0YDctCdHIhlj/4aXci1C2PvIxkG4RwFuj4jZIkIgemlf9kDnbc5n6re8TBm
fjDZ/6MMW/WDJf/W4FNX1JD7lAmZsHTGmJzbwI4UIkc0M/YeIuSTCAmkmNRQs3Hf
614ccbkA7E7bsmHjtvOuODPlw69v8jfDFOBY1LyPmb8HDzan3i8ZsLG9b1hGTMMU
su8DLF6Mo6eXgVE6Crxpymet5m5pyL8fsn7u2UL6SmogcOtNIMgbAzZEidxz12fC
aZf1tcT3EzMBJG3yXJ0yl4id86I1sf74B5+MhVyPQ6vbkOtY7ZxVPI/lsZvHq+je
vlbQbogdPK6XGIMgWOHno5IiL36kg+d/5cHtaNINaaVdNotdgLc4RAwkaib5t4EI
Ry/vbpk/PWBiVAlI3x8XxleJrPSnyVu9pIH2tHBGfdQwmTkEGVRC77lf4XoyXugJ
wv3/bByD4TW5whb35I1hES9phLUdCsg8Y4RaxPeAOFOgtVqkjZdJUzKHZL2wOKf1
Wd9NaDhQCIbGJis1Tln5RqNtrx5PNyKhK/j6X+XHyJQTF9OKakHpZQ2N+Y1iqCYV
qJBSGkgcxxd6+Gi/l93S1ah0vivNx7nisc70EGsX7lUdzrauMyflGeaY8dxizQeX
1TzYH/EZs54od0vzUGlzY8OMcSKNMZpblyCkBvWnbLO3jYsAwZ6dUduWAoYo5DQB
aIlxD+d71KWogh6DTOJ0V3rolsvUcv0qJTAFGEFyQpHfN1ZZKWyz/CYa8kuFzUBa
Bqv51AHzNyerEJvCMaT9dJxyjlpmxhPEnjwbnjXeHInBcxbeumuAK6lhXBjgvohQ
edZaNtDzr2NvoQtwlCKSv5scqSlTWRiGAMcP3FPpFEraOVwXN+FGeFBi2JuHKx8v
jTZULxpPMp8RlE2ANQPcZZQBMatHs6AvWVEPyWiUJfPELNplpd3AuqCPCJOqpKja
X2t86jWhbDa7FszvjNEgnuzRCbFvm5oC5YqvdO3p4lLz7UHCpp9nm12GFy+KmK/r
oQ2SZ+y1bHBgsbl1Rf3FcfnakdeGpnXgvGNoGLOe/3cPQhszURt/0pXzJcfhwFCv
gqkZ8Kt15Oa+gFBByYFiKDxZFQscrnZMjOIJQkLusGONbNsJe6hIUl88vcZT0Irn
P+Ek8wxLC1neF/+Wb896UY/YIbzvoImBxXCw4+hLFCVTPV807kJhpl82Rez4psRc
EVWw7GiLJDmRLV8IM60Xcjz9WbUJedUGxPNRAmQAtuxuXHVUbBAXNNdMR22kR2QN
B597vjeMDSFH1Er33wQrlVJZT50F216glgOSyY0Km2P20V99pBBjwECGDDyRsg9K
oRmFw9uDBem65KjfBcTbB+/rJTP0mOrZlh5S4rkD6d80gbuwAB5tURzl9Ob4+CXl
Eks9n698z21jFFBnssR07UwI1Uut+d5ikspM9b3d9psJ125V12dsS4vbU7lqvx1V
jJqf7WVDj1+bwlJvgsXa4uDhTFuqcTd7fZYKW5cEWxSMPv//Y7CBI6IbiaiUGcFD
or4SOs/c6X/52J1tiGFGk5QOyGd0lfaZWdsY9XsZvdze9AhEbe0aKcOtILW6EnNX
tf6+2exmkhoV8cX8YNZVdzVTYznGcsP8+Oiq/SYbJo/R7XH/FBR0jQ4itVS5VTbA
ekKHwWQJq9ET7UFdk8lnYlFgB6I8YL6HDzrL9w1VB4YOX1fO47OUGfBudlLk59KE
GZI7HcTYC6k9kJEMDBGaHBufn0XeUGzwCW6y+6HkBhi4wVXDKfJyWfRHI/D/r3m4
tQnqjnalWxPMBbeVuLSI26OOVwARwlhq+SAOi3JRpRlWMPJUHpX6eDzAOwSc4ksQ
9qCZ7g2tTZtRFqNPPPJ5rc+Swh3goFiVGGOJgKG9Q8zSKz9iutOoQEGELRs2R28s
6H6Y0rU+DqyEWZlJS2VaS1hGMFjRSc0taT7PuF15yesMCd2EbkgAJ43uC3pJYJVO
Hp/tSo7RHDCMCyDexVXnHBpziYxcU2JDZ8KKxPCfvj/zKsDJy7t2mY6sln1qyxtn
xSdzJGEmMvss/3JZIMmGvmxyEjP7Hg6WLrNlt7Xpeea6U2kTJ4kV92fZ6uBR5JZ7
bxJndu83LJLGubc0KoyNcYEg/yHJyjci6NmfJfFbICxo5/imFSaWuS370QHIlLG9
eGdbemDUImYZ9/T6o9FCrROCWDrKrOTIuD7Tq7k0bxla013h4+9q6f94P7d5loLW
MapXr3zudoPcjyc97tVEsW4juy9rNn5AIHM+mqxFKRpM/rt1sVJhEAbaslgTvU8n
ZGGDflcd2KIpJ8H+tOLwfQhjzAyvGyoD1zCz6engpKMTxWT3AtfvCfqrJ02a9g9D
d5grvY5Jo2nclwuqjsOobooja6DQwgYGhC9ODCUuKYLatIoABvbXbuT5GWE02vCI
xjGC/suTqHDuXht5XWVHRdT+e3ay5uo5DKR3h5jM94kwTKr7r6BKBIlsTu0WTGg2
WnRgyErECwwHTZHobuCFajlX3PEgCFVhwdE/5s8c5kOnan7+7Xsdb8d6NDE8M7Ut
KfrSw4YvfhR4TN+2gfeXBHr1TqRt+k4JMJwG/y6Fh7yg3ZbWUphegrhc0WbH4fmA
xyymsPXRop0/P75wwgWNvxJVsEOEtq91hn0/27jXPWxRc5fAKlIeGleHdMdF1fjl
JxBJWLvBzepe9FDZh2g18SVUWbP0HIpTfWYDFY4qEnqPy//pakmuS+7+YcHZfjhU
IjC2ve75bTmc2vIQI0Xnk1zhg5WvhWSf3YzD65IBGiaNZxi7OLizBaSH6dbvNhUz
uVLN+Do609UWdZ53eY/ejdvV84Jxol1zVLh1Rx/ucY67UpLMcySlRITqPecVmEob
IJTr7dCiIafQ7rRdqvHijMwmP9rjOCDMCUQceP0KkyP2mnCuhDrMCPtC9y0CYegc
pV1KvwmJWlq/Tr2t8f0uNU1LQkDOR88njRc8RSOpoWQQosFUlVyLPA3H3H8Z0y+v
ek7ybF0BbPJDv9Ft8U+mErXaK72bkED2IApSscb8ZTWHkhJhr/VD05bLhqFjODcv
Xqj3JD6Ho57V0mWk0iX8YvhBpF8Lrwuf81FqwIwphl+jS0dI/wI2TR2hcgt9zzJ5
wPJ0Y8W+H0bpGlPhqG0i5ldqmgDSUCtC4tGEZMLNKs4RbTmTRSqDfLEQ6YaH0axn
0LrX0fYrQpWST6gNzwapAW/3dMYuQcu9pN341Wp+0klg7E2H1JH3d6KHyUe1FMc2
/c89Ywsxpmp9VOALYNLfn6lL9BIxsuVLkivhgASeirB6RkjRXXXAV7g7upJwQwnz
5GTZ7+Wra30kE08eDJV5/CSv8VEovPJloW8dDw8w3/60FD3DpWL+KY0WtIOWMQK7
U/IqY5BxTFn7RR8eM5KJrA2SLcmKVm4KaXVaaULCCEmgb7n1SdFOFYHvukZ0mSCV
W4HwoiIvgzWqEdxVOhqh8/r/+SCPiaNtIAQLTnvl3+IVnxjboiX2akYHgyP8BpC0
i2ttD0cvq9dSQJ+JIIXMolEmBt5fT2DhDtJBLtQ5jHtVEEZYbvSaSYM2AilLqj1l
OYUCmRpIjc0lD51ZWA/3HQdlWL49C5VYM/FlAB+18Jglv0VEu1jjxe969NRp0EAk
cBUajyQoQM21XXrGOccUTAg/WsfcUFXsAkr06Wh8i8C1RR1+1AFdouqMeBd7Ch5U
9lQQyEYztsgX+xsz5HDYnIyjJNWzhswl7FynVTFDPUZ4IbE+4mtzK352rgJh1ApK
PSbtMG8DXa58vwvBZPT9VwgSqBWDnrmcOdm8oc+0CZPToGDvACubLhaIgGNhc0w6
lIkYt+Kh4Ktbqd5L0mswyTrVDEuW2lnoJF48LQY+jQkKWO4iNJoCegkb2KiK2usb
U0fCdloEdYOmPI9kro10QMQPApitGdQo4W5ZGM7N7lbn51ogiw4D70PK4y81z9pF
v8K18Ni8DzEddmRRfNpPJlFehdLBChIEUmGkKrdrMJRVeluW51hln6uYSIozSKAO
pHsEpxEPuhn7T7vr6QE4+QhnSeoyfRSsrToxP77wSN7v3DmnnATGbjtdvzWc5tPD
VB0y2uzhird9EPog+0+g7jqqDcrG5z9lkhl+prr6eh0V6NJeE3X0set8Tx0M7br9
aFkq0brVDhSRU4us7Gyal8Oeb4gQj7qb7oMe5Ev8lV53w8VrYze3K2aLo6Mlsb+C
b2fiDrhT0lEaT+1MuEyuZo7XQ1fXZFPXEkjd0GBK9XmIs7aImlXdRQogh8Pj0teO
7FeHlfSre/iFtm+YlGu7RLnRKa08nG7Xmyz3MHWPyKWqtYeo5zULBVclUE4L6Vw9
+oiXjWjEaIR0JCq7127+/XXHRYi6igp2s7ZtORYfHmgfFynHWeNhDmR8PlbcTGJW
C6hgqqhDvxL7ZpJnG6zq0CfkK5qdOxJh/skv31283KxzLFuuA2J4lau0Y1b3wizS
yklFFwt9z2+gLs3VZHfmFJuvRj0LCXgDCF0jco9Fo5EwTluP8eCI5NBGAYgYjfXl
9MmOs3kZVV8Uh1OFrI3J8jxAjCM2E3bJ/c9dDIBwlE/pqEZT/G5uayjd2DokWN7w
q+LP8Dh1nTAR3dPnUG3YQpHFbfNdMSUoj9pG2GOE62ucYJqblMEB6p/MvWvaNzkq
xpIcCsOBgrL/1Z3v+j1dfolvk+PV8IzZtvKXZql6mg0QDL7vLwTe5C5kfcKuKA+6
TDG4hfnbqx1oRaKtnW9P5xP9GRqkJgsB2jt/tTCdHhqgALfLNof1lJvZmEZMZg+H
UGjCnzgJd08Uqr4fEJFYOeHHckQKaL9NE85KfjICXizlfhvksvPB52qthGdlOsvW
SC12/ZHYhA+heNfF9HWFJZONkkw0+g49zF5SV79jMY7m83m5SjOMmWtTWfx/pk6A
SONZHbUycu7H3Jb90HozdA==
`pragma protect end_protected
