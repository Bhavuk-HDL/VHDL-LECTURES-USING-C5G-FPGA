// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:22:14 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
dBj+q+ospWWh1q519TKfwbpMyfWwS43ryVswIRrhowrlqGZdAL/bZMzqfcn5KZio
lqn2ArXjh6rFrT293Vsdy16Mvj4evEPKhXB4Dw1tYKSnroHuajvessCfB/kX6lQF
e/MGsko1mrUKowXVcEBhLuU0HQYgPtY0+GXsqk+5qDw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 4352)
RGx8BARMkTcdsEDDT7uI2KSRVJRgCa5+2Vwy9NFIaE51V+3xooyF5Corest6LpPe
A7sShF74Auh3Vko5WtRf56D+c56oO07O3X5YCR0e4MAss1eXXH7Tm/SNPBxlqSuG
GtT9X2MghcDIa15Opj4cmWV0cPQBvSaMcWurj+EDOF2dBDGUxvk8tNl7BGCd+5CF
hS5Sz23NTELv6BXxItRRVurgQZa/xvNLyv27SImamslIUwUwbtPJS9S/lu8RP0JH
yp0nB05cYNf5QQQVOwuRQLki463SONBXWF7gUMo4N4Zu4DOoR3DCkjHzVZAp6v3u
5M0G404FM+LvpzW7l1ZxSs0itC72rNNGsHTe+zsz1y1qOXhBqbrVKh3S1gekqfxD
YNT38fbEXYjIEniRHkIguga0UKr0/+B+XpdwPL3WCJdeivbY6ploAW9HW4VXwaZt
8u+HZhpy8/eutReS7eTSRHYQoj5iyi/5YSimSdl8iQxa08bgrT7HriHP/sBKXQuA
B6Wjou8+DJqxa4454Fkd8dminpoXDY+sqIv6hknwQNy31lF/9THPpldgpa+DtMrn
1Pk8tboo/6fwvRSQnQLLoq8XXiq2VuChI6gffqR89trQMeVOqmh5QZIeMjwI+m6V
/njAWTfdh7zk9H/78gCSFcGZIKGOqRPCwiT4ZF1ZXnRAtPXxXO2qzLc4916gpJFc
tJ90F7KrYq9X0gxqapYKG33x6ZAqYta7Dm6lY0GabgpjZse78XiDaI3Bphb6QRwc
AbH+CEUBD48w13pErbg660yW4HUmEhiek/iIkQgVuOv6PDGQ2UPcZLcjERQsn3Ku
GpXWt7KPuQDR/Sd+y/O64k+d5lDhz8iAChwQJBwA1Sy5bBsMoh5Zw6RZYSqLXQSt
L9NOgABaFMGtAnpL8O1mNvrT1CdSMMNE+Oj361xs8NRF78dKc7KAbpWLbXmbT8L/
Oj1GOV5kxKun0jpB0eCYIhoJlL116bTLBbtX+0fHkk7dqtoA65+3pL6IZGVMpGYn
wfiY2tmMX4xUvCHgQ33qplPUi/4CPlYY6g/vg9WcrgNaYX/9FFlnH+PtjIsFewlN
kJ4Z3Q9H8vTwmJByklOzgZ3lNQE9l12w1e6uZ0X+l6vpksmfdc1N5+lSo0FfoiMB
B5Ja4Rg9IthKMOCpus7zPvevhA3YREY/hpMH95WAoIFf7VngctRvlxxcRPyPOvf6
KFIsGyv+3kplQpyz4R8xyGKI8iXOWl4R4xlau+jpOww6qZvHpYLpp20omAcwICy6
iBS0vRYZYCjSf9kW7TNGznGlfhMdb0iqO0xz2zWbHq0Mu0wQum21voAb0D+rZG+S
zvLUQAPYvzVDUbT9bPQNAyNMI9CqTvE72Tyil5Pws7hp2ZNL0iZqHYEUqiIt64ei
ixC5M+II2ebqCR68tNM4QZrGXdcaUmimPK4bQEAi6hs8uBWZ+N/71p99oiMCbJpu
iCcqPCB0qrRdMq6glEIk4EKZy4nj3s76/1fPHuXc8lnM3iIb8m0W+/jIEO5B7IQv
4O2OukWNf2nfwk2aWfHeloXYYCxjIGRZkVqCONiQFAzepfWNEsUR5RakPzcJD4Ax
DzcCAySxeIL+stfuH7UTPeMqTMk7TRTaHNN/r6hAhJKcVMf+z6AuX9LatU2BTCDs
yVfogoJG+UaMIZkUbyxBzpMb/rh3MwddeeTMkyz/9c0AzRvRKS/bYsz3h6919QBQ
029Qbt3YDbO9faq9XkHDdsYLpkzGf3h/GmkCLE/Y5IQKYvomJA2QFib2wUf5gNQ1
Rs4oCMKDtSNR1fyGqpRG+HXIvUY5XQIZHqukRIq7BSOkYL7YkyPqRqMjBgTeVl1o
KRG79k2pLJwK/SnY0ggZZNkO4ZYnhj4pgYbE2Gi2kBtp+CkxtDYFRGHMfT8FAXdG
j5+Idh/d2aZ0ymHiD/U5e7tvHalnI+/HS3XsAd6zk3QcqCyTboehOVA3ckow8RQL
VFCyqL1y9mO7FHa9BlJHj/Lm7iwnPZLG/AWbAsDs4CkWdZQOIsVuVjkyj0EXVTy6
WMcB9aqIRky8nmgWSaC+V8xd15n0UCeBYISprqpvF0t8JeNFWgzVXAvC4S7lgpNh
/qPLTBfYs+DTUBDALow7pO6mii0ABv27zMpFt7E5eN6MAYurJEAlB8bzQ4n9U2LN
FZvhPtedE6XyhqbDBReHbzGj926kE4IAK2Koj2etmV+WyDcmqwa9M2rwo837BVTt
+W/s5yAuLXTAoC4tarfIQ2S3/esw+volHMdORptdAkUHFcaoceenMJztppKZ2V5k
XxbVgY4dyjgK1yW5sH+lksOIaCmKPwntcf2mYY5omFIuDSI5NTiGJCcpw+opQF1T
hXuJfSHnju5GEpwjEsR6PH0FNv2f/yTVjSup+3E8OM/FcPqoog+XMnzxtAx3WA5H
O2yuwV6sxlNOsgXN9NXhxZjag4kNBrZ6sXMBxJacZB0nmmIURDkPyxYPb2RJSo26
WBNRQmCtkKOc7giDBZQQ+WTMAZyt2R03AN+qixvx29sAphlWRmAfQJZiqaPeeTik
6VbO+pY2mzfMTmMObS05i1ikYQw0nCStu1hluT9XboZ/reg902PazPDsqeENb7lw
ba1QvR+QI2mlnceMEvR0WsCov003UCjEKhVPupLDLwR4QH6VbpUvrhd0F/siY6Ga
kOfXYdFgCEEjC1gZfQ7D6TFYx4H+eHKtkfPgBpzUIzz2EyieU/LIeYphrmPZCCnw
SN3cEoVaCg40mdgd4LUTom2gVbNeMvAq/uJFzxIOjQ7clcc2tlGXw7jsLcd8OUsJ
1uys3/IRVTQK3Esmwx8eo1wd8Ff6l4IAIHwcyggo0m2wC6FFnxaPZ3/gueKaxTZx
vD9ci3IcjBCVnI7N/kbhsEO4rJRH7eeZzWRAMSMhVjNbTmRlQzmzFqgtAaA7TboH
uqdgqzS+ZxlZ8gqhbDBS1gNnZbcq1IeQ1uMsM3jhJbSjJyfZzIKLeKq+/hmvpdO/
xoqxKVodEzPhztBT8aD49/DzzLVJkdAHdLTfiuKeUlqhcBXRcfdvOycnxTqWpFMG
u1QDwcz4GSJzrhJx/Tcxyv18ymqZ/VpOKBpU9RrEHOkC4bLHKE+OuyqxV2NwNIrC
L+Fztn+52u2Eeam42XIgHlD+3XLWhlsHPc6ZeqVOsiVw+VPQ1IcN52HGkSb995tQ
e764yrgbRG+L463JvXfkoPZQsiFOcWeI6mbC0XEO5BZ47D9jKzUhpZcEKds5VH1M
olcrKCc3RYG/R4GJX0mFB3Jkeieq+UvXx/bJ4SuFuAIB35WWcU4oMILCplJ3t+6t
KGwTNDhA4uOknXJo7obndzyJXel9ugdFYGzG1OF4wVviWXf2x6sL7XkBd8zMkRun
HNa2W9kKuHzb7zfgLx2w/dmFoJi2ycotCSq/9PWt6JO0h3NB+HwZBh+03OdFmLrf
lelm1E/ky9uEOthuCCy5UN4pcshMDddeT1ut52R2Zf4Uv09+hQ9uvrR5sOHTipLT
CwySL54zILJagGqeEPg4snO5WAKcegRy1fc0yN8XqjtyeJMDJQO4PgUUtvpOS40e
9KdxB2iKDhzLFDGxQqoypWDAxMN/BPiehXOiVTc7gX4v331+DUgS7GAC644ctNRp
ejR2p9/QzRJEXN6zG2+/na/44xltS9S+Q7TDzsh3kkuEkRb/4ld8TqpNYJWHJxNm
oi7uiCu1a8aN/2xWSYiUOXzCD0CKpzWKjot4RzMbhhhEnVNpYUh6iGDzIUFr9gNj
DKGM2qlLCtYxDsOJVSLwktuU/i+k0cCQxm6JT+nczx1j+w0CLxJoBPkLXU8Ddk/Q
hFZpbjIHekA2bXHuOpqk5OJemTqUnWsLGdPY5hx8EoPtlwBEszWwFGgXhPmcQLWQ
33b7sI86PTg2zkd2xB16d0xtv5qVMR1M/xXv68dsWXJBA8z4iK5oREIEoVPqzD8d
1LaGG0bOXPvnUn0pOvsHSXqPaEnbNiz2UUH5vXkybXLcCYi5coiSlRWdsW3hgZ59
J7bz2XmpOzz4xqIRLCeQ2p0EB54w0QqaL1BnnQVEHppoR0/lGUs/Oo7iEU91iZrz
JtNpN1a/ze1JNI2miTk3M4pmrJVFbsD2I9etAmKbT+hKCpg7EBa7xfzCWPGPMJ9I
pK+6rNPqMCdG0+zyM9xgZ3mAO883PdBX5r5PGs6l8aNM1USQ6YF+/CkqPK7C5GvC
/zsE1/PLoacvOmT5mehJuvDLMTmXt6v64fpvhz6sg0f+f/8V+ofbmE0mq0nnSLde
SJr1OVeEuQrSHCPisAs1vu/G6Dwuc3TNJO66LD2i5YHbtGJ2qahcRVFf9REswKqt
0sHeP/CjZx064IhnHJfNOGoBbDOsWhuXTJOrD9UlY/eye8vlbmWALZMc/igwHldi
TWg7CE/AJPdJ8UtH4S7wqmwbmdGzOLkxNzKJY7A+tO8C22drCvOkSMZWv/GdCjIR
vxGi3xi4po62IZYYz6A+Zvm8RDi0PC1lby6GsCtWVNeUa5/KjUPlaygJoxWzZxav
3wa1XCKcppGUHfDUvwcaKc7YGwxHLRU9u2gTTdmaWPYlfa10Y9tC75jOusV4XIjH
St05tszYGtZdI3RN3zuZVbJNHDMWNhKfAqbMvuRwGTSZ4Sm13/Ho0cwPAU2Gcugl
llq7ZGgJ1CuWo/yHPCYRPVzPN1OeG5mWlOWnaq/UWhOtNoPyQUrK6WkpWWOOAHYI
adw6QLDGRxCbhHuKdvIjwfHU4vd17W+UJrI5t5ym1OGe1RL1oFr/uJO6ItQ//I+f
EH4kl5XhuTZ4q+5R+Xu8HU0s893rnr6vROMkz0veIT/SpdL0S82EIvFZTiwKiFmj
WasWi+9M7rvjwZy7z5m6JbONCaApdQ+o8LVUHky5T7mCEO7am8l5p9XTxndN4Djl
rZpPwlKax82/W4vaaKD1WI3W3GW4zevw7MQJx4kfZDK03vXi7FayA3OlHp/hnmB2
vUiOKqtx0nljiS4fx0ggkrkj1cchbX5OWKg3UyaEHxJ6AXH+w7wmulhCqL3dl1z/
X0TU2vLdNOtcyAE4vHLXc/1le+nSPhD3Gkh7vwSmuG6uO4U3h+lVlVsowQnmWrkK
MZJK/yrAMmiGbXUEQRCBl9CbPjNc9jEMsOvdh+TuF10jVdm/8ToooEXhcmAz+qV2
FSuLAD1z3xxc7YbTP669Zy3qS/kb9CbPWePN+dsLGtTmtGbpP9oeUlvBjZDx954o
hI229aev0eGEMEo8dMcXaWmGJ0R/kxcYqGzRJSNw3zqExYiECSZU9C5Gx86yAjvl
28O6S2ibd+eFN6lbzLzpKeQiOq3qH8A6tEksXwADg62TtnkVxpivL92c8tXefMFe
DkukP0cSZDC85OgSaWe5b0soZio4v8/8brBBZAWdwrtZ3y1/7BdPWkLpSUKRwL4E
M8pGtBzhWZHQkfDUNnVlBFZRsJQrrcqWH7OcP6UHTLmtD2ojsWexihvqeu4FU8i5
9hGeLnsfqUnqxCuVS63iSSZNH8TfaFUWhPx1Pu4BWZ50SIR5hNBQLvR0suTQUZID
yIs6qB/ysDOEFhtmp47T5WYFPw9Ar2npY1qP7QAYyo728J220GyQJVAKVUbPxf8N
K5j94POAAFKIHTQDMzgohakSVbs04xKY/fAnvr8EvkAcdo5UOYMEN3zE+J7xi+Hl
rbmJoufgU85e+hCGU6WitL2EusmfwGGLtFe2R9AOT5As7eTbsORvFbkLUPWu8Wex
UDnLvZIcZggVGu4uf7ZUpsy1R7WSfb8srM8wF9bOKv8=
`pragma protect end_protected
