-- LPDDR2.vhd

-- Generated using ACDS version 16.1 203

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LPDDR2 is
	port (
		pll_ref_clk                : in    std_logic                     := '0';             --        pll_ref_clk.clk
		global_reset_n             : in    std_logic                     := '0';             --       global_reset.reset_n
		soft_reset_n               : in    std_logic                     := '0';             --         soft_reset.reset_n
		afi_clk                    : out   std_logic;                                        --            afi_clk.clk
		afi_half_clk               : out   std_logic;                                        --       afi_half_clk.clk
		afi_reset_n                : out   std_logic;                                        --          afi_reset.reset_n
		afi_reset_export_n         : out   std_logic;                                        --   afi_reset_export.reset_n
		seq_debug_clk              : in    std_logic                     := '0';             --      seq_debug_clk.clk
		seq_debug_reset_n          : in    std_logic                     := '0';             -- seq_debug_reset_in.reset_n
		mem_ca                     : out   std_logic_vector(9 downto 0);                     --             memory.mem_ca
		mem_ck                     : out   std_logic_vector(0 downto 0);                     --                   .mem_ck
		mem_ck_n                   : out   std_logic_vector(0 downto 0);                     --                   .mem_ck_n
		mem_cke                    : out   std_logic_vector(0 downto 0);                     --                   .mem_cke
		mem_cs_n                   : out   std_logic_vector(0 downto 0);                     --                   .mem_cs_n
		mem_dm                     : out   std_logic_vector(3 downto 0);                     --                   .mem_dm
		mem_dq                     : inout std_logic_vector(31 downto 0) := (others => '0'); --                   .mem_dq
		mem_dqs                    : inout std_logic_vector(3 downto 0)  := (others => '0'); --                   .mem_dqs
		mem_dqs_n                  : inout std_logic_vector(3 downto 0)  := (others => '0'); --                   .mem_dqs_n
		avl_ready_0                : out   std_logic;                                        --              avl_0.waitrequest_n
		avl_burstbegin_0           : in    std_logic                     := '0';             --                   .beginbursttransfer
		avl_addr_0                 : in    std_logic_vector(26 downto 0) := (others => '0'); --                   .address
		avl_rdata_valid_0          : out   std_logic;                                        --                   .readdatavalid
		avl_rdata_0                : out   std_logic_vector(31 downto 0);                    --                   .readdata
		avl_wdata_0                : in    std_logic_vector(31 downto 0) := (others => '0'); --                   .writedata
		avl_be_0                   : in    std_logic_vector(3 downto 0)  := (others => '0'); --                   .byteenable
		avl_read_req_0             : in    std_logic                     := '0';             --                   .read
		avl_write_req_0            : in    std_logic                     := '0';             --                   .write
		avl_size_0                 : in    std_logic_vector(2 downto 0)  := (others => '0'); --                   .burstcount
		avl_ready_1                : out   std_logic;                                        --              avl_1.waitrequest_n
		avl_burstbegin_1           : in    std_logic                     := '0';             --                   .beginbursttransfer
		avl_addr_1                 : in    std_logic_vector(26 downto 0) := (others => '0'); --                   .address
		avl_rdata_valid_1          : out   std_logic;                                        --                   .readdatavalid
		avl_rdata_1                : out   std_logic_vector(31 downto 0);                    --                   .readdata
		avl_wdata_1                : in    std_logic_vector(31 downto 0) := (others => '0'); --                   .writedata
		avl_be_1                   : in    std_logic_vector(3 downto 0)  := (others => '0'); --                   .byteenable
		avl_read_req_1             : in    std_logic                     := '0';             --                   .read
		avl_write_req_1            : in    std_logic                     := '0';             --                   .write
		avl_size_1                 : in    std_logic_vector(2 downto 0)  := (others => '0'); --                   .burstcount
		avl_ready_2                : out   std_logic;                                        --              avl_2.waitrequest_n
		avl_burstbegin_2           : in    std_logic                     := '0';             --                   .beginbursttransfer
		avl_addr_2                 : in    std_logic_vector(26 downto 0) := (others => '0'); --                   .address
		avl_rdata_valid_2          : out   std_logic;                                        --                   .readdatavalid
		avl_rdata_2                : out   std_logic_vector(31 downto 0);                    --                   .readdata
		avl_wdata_2                : in    std_logic_vector(31 downto 0) := (others => '0'); --                   .writedata
		avl_be_2                   : in    std_logic_vector(3 downto 0)  := (others => '0'); --                   .byteenable
		avl_read_req_2             : in    std_logic                     := '0';             --                   .read
		avl_write_req_2            : in    std_logic                     := '0';             --                   .write
		avl_size_2                 : in    std_logic_vector(2 downto 0)  := (others => '0'); --                   .burstcount
		avl_ready_3                : out   std_logic;                                        --              avl_3.waitrequest_n
		avl_burstbegin_3           : in    std_logic                     := '0';             --                   .beginbursttransfer
		avl_addr_3                 : in    std_logic_vector(26 downto 0) := (others => '0'); --                   .address
		avl_rdata_valid_3          : out   std_logic;                                        --                   .readdatavalid
		avl_rdata_3                : out   std_logic_vector(31 downto 0);                    --                   .readdata
		avl_wdata_3                : in    std_logic_vector(31 downto 0) := (others => '0'); --                   .writedata
		avl_be_3                   : in    std_logic_vector(3 downto 0)  := (others => '0'); --                   .byteenable
		avl_read_req_3             : in    std_logic                     := '0';             --                   .read
		avl_write_req_3            : in    std_logic                     := '0';             --                   .write
		avl_size_3                 : in    std_logic_vector(2 downto 0)  := (others => '0'); --                   .burstcount
		mp_cmd_clk_0_clk           : in    std_logic                     := '0';             --       mp_cmd_clk_0.clk
		mp_cmd_reset_n_0_reset_n   : in    std_logic                     := '0';             --   mp_cmd_reset_n_0.reset_n
		mp_cmd_clk_1_clk           : in    std_logic                     := '0';             --       mp_cmd_clk_1.clk
		mp_cmd_reset_n_1_reset_n   : in    std_logic                     := '0';             --   mp_cmd_reset_n_1.reset_n
		mp_cmd_clk_2_clk           : in    std_logic                     := '0';             --       mp_cmd_clk_2.clk
		mp_cmd_reset_n_2_reset_n   : in    std_logic                     := '0';             --   mp_cmd_reset_n_2.reset_n
		mp_cmd_clk_3_clk           : in    std_logic                     := '0';             --       mp_cmd_clk_3.clk
		mp_cmd_reset_n_3_reset_n   : in    std_logic                     := '0';             --   mp_cmd_reset_n_3.reset_n
		mp_rfifo_clk_0_clk         : in    std_logic                     := '0';             --     mp_rfifo_clk_0.clk
		mp_rfifo_reset_n_0_reset_n : in    std_logic                     := '0';             -- mp_rfifo_reset_n_0.reset_n
		mp_wfifo_clk_0_clk         : in    std_logic                     := '0';             --     mp_wfifo_clk_0.clk
		mp_wfifo_reset_n_0_reset_n : in    std_logic                     := '0';             -- mp_wfifo_reset_n_0.reset_n
		mp_rfifo_clk_1_clk         : in    std_logic                     := '0';             --     mp_rfifo_clk_1.clk
		mp_rfifo_reset_n_1_reset_n : in    std_logic                     := '0';             -- mp_rfifo_reset_n_1.reset_n
		mp_wfifo_clk_1_clk         : in    std_logic                     := '0';             --     mp_wfifo_clk_1.clk
		mp_wfifo_reset_n_1_reset_n : in    std_logic                     := '0';             -- mp_wfifo_reset_n_1.reset_n
		mp_rfifo_clk_2_clk         : in    std_logic                     := '0';             --     mp_rfifo_clk_2.clk
		mp_rfifo_reset_n_2_reset_n : in    std_logic                     := '0';             -- mp_rfifo_reset_n_2.reset_n
		mp_wfifo_clk_2_clk         : in    std_logic                     := '0';             --     mp_wfifo_clk_2.clk
		mp_wfifo_reset_n_2_reset_n : in    std_logic                     := '0';             -- mp_wfifo_reset_n_2.reset_n
		mp_rfifo_clk_3_clk         : in    std_logic                     := '0';             --     mp_rfifo_clk_3.clk
		mp_rfifo_reset_n_3_reset_n : in    std_logic                     := '0';             -- mp_rfifo_reset_n_3.reset_n
		mp_wfifo_clk_3_clk         : in    std_logic                     := '0';             --     mp_wfifo_clk_3.clk
		mp_wfifo_reset_n_3_reset_n : in    std_logic                     := '0';             -- mp_wfifo_reset_n_3.reset_n
		local_init_done            : out   std_logic;                                        --             status.local_init_done
		local_cal_success          : out   std_logic;                                        --                   .local_cal_success
		local_cal_fail             : out   std_logic;                                        --                   .local_cal_fail
		oct_rzqin                  : in    std_logic                     := '0';             --                oct.rzqin
		pll_mem_clk                : out   std_logic;                                        --        pll_sharing.pll_mem_clk
		pll_write_clk              : out   std_logic;                                        --                   .pll_write_clk
		pll_locked                 : out   std_logic;                                        --                   .pll_locked
		pll_write_clk_pre_phy_clk  : out   std_logic;                                        --                   .pll_write_clk_pre_phy_clk
		pll_addr_cmd_clk           : out   std_logic;                                        --                   .pll_addr_cmd_clk
		pll_avl_clk                : out   std_logic;                                        --                   .pll_avl_clk
		pll_config_clk             : out   std_logic;                                        --                   .pll_config_clk
		pll_mem_phy_clk            : out   std_logic;                                        --                   .pll_mem_phy_clk
		afi_phy_clk                : out   std_logic;                                        --                   .afi_phy_clk
		pll_avl_phy_clk            : out   std_logic;                                        --                   .pll_avl_phy_clk
		seq_debug_addr             : in    std_logic_vector(19 downto 0) := (others => '0'); --          seq_debug.address
		seq_debug_read_req         : in    std_logic                     := '0';             --                   .read
		seq_debug_rdata            : out   std_logic_vector(31 downto 0);                    --                   .readdata
		seq_debug_write_req        : in    std_logic                     := '0';             --                   .write
		seq_debug_wdata            : in    std_logic_vector(31 downto 0) := (others => '0'); --                   .writedata
		seq_debug_waitrequest      : out   std_logic;                                        --                   .waitrequest
		seq_debug_be               : in    std_logic_vector(3 downto 0)  := (others => '0'); --                   .byteenable
		seq_debug_rdata_valid      : out   std_logic                                         --                   .readdatavalid
	);
end entity LPDDR2;

architecture rtl of LPDDR2 is
	component LPDDR2_0002 is
		port (
			pll_ref_clk                : in    std_logic                     := 'X';             -- clk
			global_reset_n             : in    std_logic                     := 'X';             -- reset_n
			soft_reset_n               : in    std_logic                     := 'X';             -- reset_n
			afi_clk                    : out   std_logic;                                        -- clk
			afi_half_clk               : out   std_logic;                                        -- clk
			afi_reset_n                : out   std_logic;                                        -- reset_n
			afi_reset_export_n         : out   std_logic;                                        -- reset_n
			seq_debug_clk              : in    std_logic                     := 'X';             -- clk
			seq_debug_reset_n          : in    std_logic                     := 'X';             -- reset_n
			mem_ca                     : out   std_logic_vector(9 downto 0);                     -- mem_ca
			mem_ck                     : out   std_logic_vector(0 downto 0);                     -- mem_ck
			mem_ck_n                   : out   std_logic_vector(0 downto 0);                     -- mem_ck_n
			mem_cke                    : out   std_logic_vector(0 downto 0);                     -- mem_cke
			mem_cs_n                   : out   std_logic_vector(0 downto 0);                     -- mem_cs_n
			mem_dm                     : out   std_logic_vector(3 downto 0);                     -- mem_dm
			mem_dq                     : inout std_logic_vector(31 downto 0) := (others => 'X'); -- mem_dq
			mem_dqs                    : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs
			mem_dqs_n                  : inout std_logic_vector(3 downto 0)  := (others => 'X'); -- mem_dqs_n
			avl_ready_0                : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin_0           : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr_0                 : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address
			avl_rdata_valid_0          : out   std_logic;                                        -- readdatavalid
			avl_rdata_0                : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata_0                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be_0                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req_0             : in    std_logic                     := 'X';             -- read
			avl_write_req_0            : in    std_logic                     := 'X';             -- write
			avl_size_0                 : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			avl_ready_1                : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin_1           : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr_1                 : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address
			avl_rdata_valid_1          : out   std_logic;                                        -- readdatavalid
			avl_rdata_1                : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata_1                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be_1                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req_1             : in    std_logic                     := 'X';             -- read
			avl_write_req_1            : in    std_logic                     := 'X';             -- write
			avl_size_1                 : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			avl_ready_2                : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin_2           : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr_2                 : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address
			avl_rdata_valid_2          : out   std_logic;                                        -- readdatavalid
			avl_rdata_2                : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata_2                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be_2                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req_2             : in    std_logic                     := 'X';             -- read
			avl_write_req_2            : in    std_logic                     := 'X';             -- write
			avl_size_2                 : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			avl_ready_3                : out   std_logic;                                        -- waitrequest_n
			avl_burstbegin_3           : in    std_logic                     := 'X';             -- beginbursttransfer
			avl_addr_3                 : in    std_logic_vector(26 downto 0) := (others => 'X'); -- address
			avl_rdata_valid_3          : out   std_logic;                                        -- readdatavalid
			avl_rdata_3                : out   std_logic_vector(31 downto 0);                    -- readdata
			avl_wdata_3                : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			avl_be_3                   : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			avl_read_req_3             : in    std_logic                     := 'X';             -- read
			avl_write_req_3            : in    std_logic                     := 'X';             -- write
			avl_size_3                 : in    std_logic_vector(2 downto 0)  := (others => 'X'); -- burstcount
			mp_cmd_clk_0_clk           : in    std_logic                     := 'X';             -- clk
			mp_cmd_reset_n_0_reset_n   : in    std_logic                     := 'X';             -- reset_n
			mp_cmd_clk_1_clk           : in    std_logic                     := 'X';             -- clk
			mp_cmd_reset_n_1_reset_n   : in    std_logic                     := 'X';             -- reset_n
			mp_cmd_clk_2_clk           : in    std_logic                     := 'X';             -- clk
			mp_cmd_reset_n_2_reset_n   : in    std_logic                     := 'X';             -- reset_n
			mp_cmd_clk_3_clk           : in    std_logic                     := 'X';             -- clk
			mp_cmd_reset_n_3_reset_n   : in    std_logic                     := 'X';             -- reset_n
			mp_rfifo_clk_0_clk         : in    std_logic                     := 'X';             -- clk
			mp_rfifo_reset_n_0_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_wfifo_clk_0_clk         : in    std_logic                     := 'X';             -- clk
			mp_wfifo_reset_n_0_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_rfifo_clk_1_clk         : in    std_logic                     := 'X';             -- clk
			mp_rfifo_reset_n_1_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_wfifo_clk_1_clk         : in    std_logic                     := 'X';             -- clk
			mp_wfifo_reset_n_1_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_rfifo_clk_2_clk         : in    std_logic                     := 'X';             -- clk
			mp_rfifo_reset_n_2_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_wfifo_clk_2_clk         : in    std_logic                     := 'X';             -- clk
			mp_wfifo_reset_n_2_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_rfifo_clk_3_clk         : in    std_logic                     := 'X';             -- clk
			mp_rfifo_reset_n_3_reset_n : in    std_logic                     := 'X';             -- reset_n
			mp_wfifo_clk_3_clk         : in    std_logic                     := 'X';             -- clk
			mp_wfifo_reset_n_3_reset_n : in    std_logic                     := 'X';             -- reset_n
			local_init_done            : out   std_logic;                                        -- local_init_done
			local_cal_success          : out   std_logic;                                        -- local_cal_success
			local_cal_fail             : out   std_logic;                                        -- local_cal_fail
			oct_rzqin                  : in    std_logic                     := 'X';             -- rzqin
			pll_mem_clk                : out   std_logic;                                        -- pll_mem_clk
			pll_write_clk              : out   std_logic;                                        -- pll_write_clk
			pll_locked                 : out   std_logic;                                        -- pll_locked
			pll_write_clk_pre_phy_clk  : out   std_logic;                                        -- pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk           : out   std_logic;                                        -- pll_addr_cmd_clk
			pll_avl_clk                : out   std_logic;                                        -- pll_avl_clk
			pll_config_clk             : out   std_logic;                                        -- pll_config_clk
			pll_mem_phy_clk            : out   std_logic;                                        -- pll_mem_phy_clk
			afi_phy_clk                : out   std_logic;                                        -- afi_phy_clk
			pll_avl_phy_clk            : out   std_logic;                                        -- pll_avl_phy_clk
			seq_debug_addr             : in    std_logic_vector(19 downto 0) := (others => 'X'); -- address
			seq_debug_read_req         : in    std_logic                     := 'X';             -- read
			seq_debug_rdata            : out   std_logic_vector(31 downto 0);                    -- readdata
			seq_debug_write_req        : in    std_logic                     := 'X';             -- write
			seq_debug_wdata            : in    std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			seq_debug_waitrequest      : out   std_logic;                                        -- waitrequest
			seq_debug_be               : in    std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			seq_debug_rdata_valid      : out   std_logic                                         -- readdatavalid
		);
	end component LPDDR2_0002;

begin

	lpddr2_inst : component LPDDR2_0002
		port map (
			pll_ref_clk                => pll_ref_clk,                --        pll_ref_clk.clk
			global_reset_n             => global_reset_n,             --       global_reset.reset_n
			soft_reset_n               => soft_reset_n,               --         soft_reset.reset_n
			afi_clk                    => afi_clk,                    --            afi_clk.clk
			afi_half_clk               => afi_half_clk,               --       afi_half_clk.clk
			afi_reset_n                => afi_reset_n,                --          afi_reset.reset_n
			afi_reset_export_n         => afi_reset_export_n,         --   afi_reset_export.reset_n
			seq_debug_clk              => seq_debug_clk,              --      seq_debug_clk.clk
			seq_debug_reset_n          => seq_debug_reset_n,          -- seq_debug_reset_in.reset_n
			mem_ca                     => mem_ca,                     --             memory.mem_ca
			mem_ck                     => mem_ck,                     --                   .mem_ck
			mem_ck_n                   => mem_ck_n,                   --                   .mem_ck_n
			mem_cke                    => mem_cke,                    --                   .mem_cke
			mem_cs_n                   => mem_cs_n,                   --                   .mem_cs_n
			mem_dm                     => mem_dm,                     --                   .mem_dm
			mem_dq                     => mem_dq,                     --                   .mem_dq
			mem_dqs                    => mem_dqs,                    --                   .mem_dqs
			mem_dqs_n                  => mem_dqs_n,                  --                   .mem_dqs_n
			avl_ready_0                => avl_ready_0,                --              avl_0.waitrequest_n
			avl_burstbegin_0           => avl_burstbegin_0,           --                   .beginbursttransfer
			avl_addr_0                 => avl_addr_0,                 --                   .address
			avl_rdata_valid_0          => avl_rdata_valid_0,          --                   .readdatavalid
			avl_rdata_0                => avl_rdata_0,                --                   .readdata
			avl_wdata_0                => avl_wdata_0,                --                   .writedata
			avl_be_0                   => avl_be_0,                   --                   .byteenable
			avl_read_req_0             => avl_read_req_0,             --                   .read
			avl_write_req_0            => avl_write_req_0,            --                   .write
			avl_size_0                 => avl_size_0,                 --                   .burstcount
			avl_ready_1                => avl_ready_1,                --              avl_1.waitrequest_n
			avl_burstbegin_1           => avl_burstbegin_1,           --                   .beginbursttransfer
			avl_addr_1                 => avl_addr_1,                 --                   .address
			avl_rdata_valid_1          => avl_rdata_valid_1,          --                   .readdatavalid
			avl_rdata_1                => avl_rdata_1,                --                   .readdata
			avl_wdata_1                => avl_wdata_1,                --                   .writedata
			avl_be_1                   => avl_be_1,                   --                   .byteenable
			avl_read_req_1             => avl_read_req_1,             --                   .read
			avl_write_req_1            => avl_write_req_1,            --                   .write
			avl_size_1                 => avl_size_1,                 --                   .burstcount
			avl_ready_2                => avl_ready_2,                --              avl_2.waitrequest_n
			avl_burstbegin_2           => avl_burstbegin_2,           --                   .beginbursttransfer
			avl_addr_2                 => avl_addr_2,                 --                   .address
			avl_rdata_valid_2          => avl_rdata_valid_2,          --                   .readdatavalid
			avl_rdata_2                => avl_rdata_2,                --                   .readdata
			avl_wdata_2                => avl_wdata_2,                --                   .writedata
			avl_be_2                   => avl_be_2,                   --                   .byteenable
			avl_read_req_2             => avl_read_req_2,             --                   .read
			avl_write_req_2            => avl_write_req_2,            --                   .write
			avl_size_2                 => avl_size_2,                 --                   .burstcount
			avl_ready_3                => avl_ready_3,                --              avl_3.waitrequest_n
			avl_burstbegin_3           => avl_burstbegin_3,           --                   .beginbursttransfer
			avl_addr_3                 => avl_addr_3,                 --                   .address
			avl_rdata_valid_3          => avl_rdata_valid_3,          --                   .readdatavalid
			avl_rdata_3                => avl_rdata_3,                --                   .readdata
			avl_wdata_3                => avl_wdata_3,                --                   .writedata
			avl_be_3                   => avl_be_3,                   --                   .byteenable
			avl_read_req_3             => avl_read_req_3,             --                   .read
			avl_write_req_3            => avl_write_req_3,            --                   .write
			avl_size_3                 => avl_size_3,                 --                   .burstcount
			mp_cmd_clk_0_clk           => mp_cmd_clk_0_clk,           --       mp_cmd_clk_0.clk
			mp_cmd_reset_n_0_reset_n   => mp_cmd_reset_n_0_reset_n,   --   mp_cmd_reset_n_0.reset_n
			mp_cmd_clk_1_clk           => mp_cmd_clk_1_clk,           --       mp_cmd_clk_1.clk
			mp_cmd_reset_n_1_reset_n   => mp_cmd_reset_n_1_reset_n,   --   mp_cmd_reset_n_1.reset_n
			mp_cmd_clk_2_clk           => mp_cmd_clk_2_clk,           --       mp_cmd_clk_2.clk
			mp_cmd_reset_n_2_reset_n   => mp_cmd_reset_n_2_reset_n,   --   mp_cmd_reset_n_2.reset_n
			mp_cmd_clk_3_clk           => mp_cmd_clk_3_clk,           --       mp_cmd_clk_3.clk
			mp_cmd_reset_n_3_reset_n   => mp_cmd_reset_n_3_reset_n,   --   mp_cmd_reset_n_3.reset_n
			mp_rfifo_clk_0_clk         => mp_rfifo_clk_0_clk,         --     mp_rfifo_clk_0.clk
			mp_rfifo_reset_n_0_reset_n => mp_rfifo_reset_n_0_reset_n, -- mp_rfifo_reset_n_0.reset_n
			mp_wfifo_clk_0_clk         => mp_wfifo_clk_0_clk,         --     mp_wfifo_clk_0.clk
			mp_wfifo_reset_n_0_reset_n => mp_wfifo_reset_n_0_reset_n, -- mp_wfifo_reset_n_0.reset_n
			mp_rfifo_clk_1_clk         => mp_rfifo_clk_1_clk,         --     mp_rfifo_clk_1.clk
			mp_rfifo_reset_n_1_reset_n => mp_rfifo_reset_n_1_reset_n, -- mp_rfifo_reset_n_1.reset_n
			mp_wfifo_clk_1_clk         => mp_wfifo_clk_1_clk,         --     mp_wfifo_clk_1.clk
			mp_wfifo_reset_n_1_reset_n => mp_wfifo_reset_n_1_reset_n, -- mp_wfifo_reset_n_1.reset_n
			mp_rfifo_clk_2_clk         => mp_rfifo_clk_2_clk,         --     mp_rfifo_clk_2.clk
			mp_rfifo_reset_n_2_reset_n => mp_rfifo_reset_n_2_reset_n, -- mp_rfifo_reset_n_2.reset_n
			mp_wfifo_clk_2_clk         => mp_wfifo_clk_2_clk,         --     mp_wfifo_clk_2.clk
			mp_wfifo_reset_n_2_reset_n => mp_wfifo_reset_n_2_reset_n, -- mp_wfifo_reset_n_2.reset_n
			mp_rfifo_clk_3_clk         => mp_rfifo_clk_3_clk,         --     mp_rfifo_clk_3.clk
			mp_rfifo_reset_n_3_reset_n => mp_rfifo_reset_n_3_reset_n, -- mp_rfifo_reset_n_3.reset_n
			mp_wfifo_clk_3_clk         => mp_wfifo_clk_3_clk,         --     mp_wfifo_clk_3.clk
			mp_wfifo_reset_n_3_reset_n => mp_wfifo_reset_n_3_reset_n, -- mp_wfifo_reset_n_3.reset_n
			local_init_done            => local_init_done,            --             status.local_init_done
			local_cal_success          => local_cal_success,          --                   .local_cal_success
			local_cal_fail             => local_cal_fail,             --                   .local_cal_fail
			oct_rzqin                  => oct_rzqin,                  --                oct.rzqin
			pll_mem_clk                => pll_mem_clk,                --        pll_sharing.pll_mem_clk
			pll_write_clk              => pll_write_clk,              --                   .pll_write_clk
			pll_locked                 => pll_locked,                 --                   .pll_locked
			pll_write_clk_pre_phy_clk  => pll_write_clk_pre_phy_clk,  --                   .pll_write_clk_pre_phy_clk
			pll_addr_cmd_clk           => pll_addr_cmd_clk,           --                   .pll_addr_cmd_clk
			pll_avl_clk                => pll_avl_clk,                --                   .pll_avl_clk
			pll_config_clk             => pll_config_clk,             --                   .pll_config_clk
			pll_mem_phy_clk            => pll_mem_phy_clk,            --                   .pll_mem_phy_clk
			afi_phy_clk                => afi_phy_clk,                --                   .afi_phy_clk
			pll_avl_phy_clk            => pll_avl_phy_clk,            --                   .pll_avl_phy_clk
			seq_debug_addr             => seq_debug_addr,             --          seq_debug.address
			seq_debug_read_req         => seq_debug_read_req,         --                   .read
			seq_debug_rdata            => seq_debug_rdata,            --                   .readdata
			seq_debug_write_req        => seq_debug_write_req,        --                   .write
			seq_debug_wdata            => seq_debug_wdata,            --                   .writedata
			seq_debug_waitrequest      => seq_debug_waitrequest,      --                   .waitrequest
			seq_debug_be               => seq_debug_be,               --                   .byteenable
			seq_debug_rdata_valid      => seq_debug_rdata_valid       --                   .readdatavalid
		);

end architecture rtl; -- of LPDDR2
