// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:43:28 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZDmvScyrwL3fYLzlaFOm4qdt0bVFD672yvKDhaYKwfb6Pek9s3hiZk9HjwyqCqPl
EdGUoY5DHJkFAZROdYVOqZV6UvUOVo1Q40brpu11cPnRX+V84PgtimQc/lFVCIbD
yNbO5B39510j1dEiYGoPc3jCpOWN2C5+vkQwEi9SxK8=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11488)
3IAVBm14lKoOyR0A5YERTvvup2PRs0BFIQRU6UxBj9lcC8bhJHYZckZOep+dDza5
vPexZLJhjZkyMu/0upyVvJmMWhoS56My5r8SpduPxvgns3c9ANr6+irWbODygzBZ
R5SvzbttflPtFsYe2BYes6STR8nGfA9aGFGQr6NKjddieKEmYmLxzdNmfyy7wi3Y
mAZDVD41omh/5uI3YWwTsbfQG+d4gDVLGJ7CNV1bf6wN9YxjXIEq5NBf8XMk8VPC
QV5uZoxyBEsL3Ya56jd+ir+DZdtZoN8iGYzfL9jfwDu//KPKgQSmZnxgOeSSsLgq
8jQ/GFpL1hY05muMmJzw/0lcaQwSwVYiFP1ueifNIWrNn+wOJ0Qmah9D6BQROk+g
n87bFMYvYs9f3+bMc72PflZjvzOa5fbO0KupipzdLkeBRyFkmQay516h1KTYnGjX
LJvhq6UG1KhKL/fWIAlenR6OWc2r/3E1apOAytM8cdv2cFsrYugCEcKqTWQc792n
OUNKLmRRUghI3WSo5K5mCwa77Pkzp0Cf7bfVSNnmJJDs4ntERczdAB+jt656EJKU
o/6I3dTSzeUqYJ+9Ap1XdeYKS8GAFiTH9wpNNfLMNfUI1ttxG8Y0tMHA05Ea1o79
CgrsOIizJTrkENEO1c5gnwI1GcqIOxSv4YYut9ZRxCDbbI9hZ7np4+Fk+1cXsI8m
CfXfSNnGFJGtG493VbRE5cQG0E8+7q+S1NNBKPICmiCyXvim7xewLKBEuzNjZ584
uXJ0Aq1ZLoDTCB9SYq5LjD35jbAz2nBRnhIy1PLIdqxJ0jZmvYEY6zSB10rAzZ4T
73cewLgjkV42ls9NHQOflSE4XLDtgmzDcdGxu1IBT+0bVRk402MVi/r54GyDPErg
gJJlBVUW0LVm/li+DvQmmdCRnQbg+okRphFevTlDtcPo5nJXv33QxvUCz173iQal
lZc5dj+qVRskP3by1jhZmrjrF52cbnK2xqC158DdEfHXt/oQCzbSyabZZC5jTqUb
GZ36IsbaUGnosx7VO6hesMIF/Zulr92V8EKK7ojggKw3lnx+EUh0CAneGu5HSHVv
JT5WnMxSmi8m+XPnHb/hhzCDOFOilvfOT/JBzb8sJvOZ6ANIyLUPhSLaoV9dChja
gXhQUiWar1dK1FaBq5cVYf9l+JAE2g6LFuY3gUkjADiElM0Rdz5/2uQHq81xirXU
i8GcOuUO7SJ3hQm8uOJ80kYxih52BJs0t7qEd86lDUFuRQ+YLlAcimWXM2IQsrrD
5oV/LL4v7RtXwfPr7z10iHfw88vZ8LV7dRZ21gO7y7AHpB1UxOpaMQEwWrjenfqG
ojsk6ZZanKYfZmAPw9dILj/7skdqbGdhCbXiYZppURDRpm+NoNMseTAV3Y1O1Aae
qFbUvNhAkx2MiyXdZ1f/ERy4fOezvuc2r6PmoxfGpLQvpdV3tnDIOWMe779OE3Gh
m4DTDgRh2o/wP0g3XiHn/9oISyqcPxXkEdUT+DNWiDNM58MbPiCVnZRHEbMkRTSj
1rxg/pmYHsW7RekDzogjp86YUEE3pbMwPy7RL9kRYjtC9gYs4CJ342PIlxlAB0CQ
UU+cnt4AIbssCMKyjajJvM4GSpAt9laFD609j5RxUEw0FuWeBqtVfPue4600OBDp
aPrBneGcG+YOyVuqiz3IL2mJ52XVan/h8NGi8kM6VfWT8XI8JRouXytKY3aBZXOA
9NWM7rTd6gaCkEE0PbA+z1xapFc4L8YCuuGrOAh9ryO1gKdY6upioWBnIbl1XyRm
yF5ETdhVWUnKPn05B7LWypQkAiDanWh6QDLMOnk2dVJnwyJT8oDs3JhFLhpI+wCx
SyZu8LM2th1+F/pTzXrT9QLZ5g3ac3BJ1S1j02AQS9Q4siF9PycvCmt4aekbWJkr
2hWKpnpKYNuHKA3rZ+z4hrM5AgTfENEZEhjrzGYoLMEvmt7SKkyLEJEkMInkSxDv
ZUL3AuRKIMsH1tn4Q5+N8yMvAMtzx+xrgtbweBeL8xkeHR4u1Kakbp+5+jxiNdBq
uuPBvvVcNo6gZnLhEqnFEmxoIxB6MyNR7lYaMQj7YF05MQilNrkjKcV0nLLmUtNv
P/IkEmHHbS1aCb67Eo6YiSRUe8+RYZm+MC7c3PP/KEtEWjPmwBaFtHsIFFE0MoqW
k18dVZl0KvkucmfVzstAI6uY6xdqJlNpABAy/gvTCcB3JMh76nsdPVsR4WdqV1R4
+xQRX8k/uMkRvv+yPGebSRs6g2Py1eYqK9eX7lPu1P1SblM42vV48YYvNCiIUZ7j
g9GZLubqNC2gvAS+QopZFIjJuIjaEeVunanhwHLyuLaHApTRNsoYFO/rcMmtIa8C
ylwMraPWUnuML1h0fyIlYRM0mxpO32HPkslo+W/7kPZWqdtYtOZpxabaL8z0H5ni
3tsLrsyPCsoqOCP6UpNu3/ycOaykxPhKl0QDddV9o6Jg1la/WUE3+S6o7wIZ9duI
+V1FkDejbFYOJJV7JwyvUNWFG72Nv4NodVq3yBlV/lknx8YTHQBwGgvesINBay0O
JpkuVbdNeRUuZ2t2mzI2UFiaI5r0J/js8iQcHo2DgQEhnsUkHF9elwOqbYYCFV42
qlIF/A5tjUznTolxTalRe8Plk572xwzBBkij8oS9B5Hsj4VHEe3yo/RjKkTnCWPX
oUuK89Lp95LAbk9Vb1jAEJ0SX8LbZSds/AMHurNd+ONV1sjsXzgMPPa4e+t9GQKI
ujqIKr+Yc32PCGx4bYDV8IOaGt09s19RkgpazKFhu5NiVbmUSUzLE/17jiWL8nKk
4ovVkW50xfYy7E3UMP8u3oALtU9wvq3hyXh2tK1tqcZMzMnKg2XG8eIjoY7vjrsP
BDABhokp8YFGKtSvH3wgc+ABOFipmD+7/A4WiIKHeKmPc/WT/MNAyTtORdESbSdK
zEjNqcM6d01acOD7sVSqpno0fwEuEJncOQ8A+Oar6+aDQUkLn71aVP40FfEyEPPF
ADUOAsOonVtk49F7BIFCIJ2vEL4Nqc9i0dikVB943U6xNH58T2OCfn8VeAnlXQw2
NnOgGEn9TiZGdk1HK6Y3fyiVUDXXBg2/BnuQHgiYTLdnJUOph86/lRS4cHdABlj3
prWh32+GX1ads6rgtufhABDCfOGhVUNYdC4lnvirikj+sB5AUk3R1wy6lQHMZuQu
lwSg5Q/qmeerVrYmfGnSJWEa3aGmp15AwnVbDcsGULpmM/2egsle98D6Pz57sY68
ICw+7+VKY+VDhfVam5T081RjQxF7TyMQatx2b4kMG9Vc74aLl3sFF0SFLm1KlYLj
f6avYq+B8INpY4dpaAxt8hInPFf3EX5lcQRouR4h43FdDG1NCn3R4yb61f5umGPv
HINYrZ09Jm5EjL7CLR1SociWYEtNpHoXy2fw+drQrM9Kys2lv5hsVxXDaG1RqQoX
ND72HARbHOEbHc2iB3UgWvZVjIDyn5L2gwawtDVaf7ME2NXqaz8k5Dl662fydC+b
+64LOSTgLSfMKDU/d9PhBrDo84mP38cR7C55lPDnGdi4LdT4f9Nt+pLVX+4RLMRY
wK6D/7VB5fyDRW129wPLkDWmJbqkZLkl6kbL/DHVtPFtBcjaZhXQFup1NGLdZFup
pwU8hagbg2/gu2GmxBvSirBmy7rnT0uoilFZRDeEMMQoYi0nMmC3sdDE99fdzUsZ
QuJQZyLqBz1XT1Rqxfvl693H16YAVx3lu5ZbZo2eUQeu8nE5YPWmrLW1zU39fn8G
/Nly+1oXilahxjrEzHxlYNNw21BVjvH8TKaptxmXUQLD5LuU1HPpZtBOsQPJvkKC
KE2TxzYOAnXvVWqKrZ/j57S6iXN81htGNWmBknmAYuZ5Dves+4F5+Mrwh9wZwDxa
NIqI93/ophHt1mROoBFAYpZD08dtGmM1pBx1M6OU6MgNh0MkH2mN4fvs/r+csnDo
xvg6wZuxusqsiTbZwIc9fxSJ+U1qGvZB7JW2cZRBf9hT8Zx42aPkuIt3yCjNJ3nS
K08zLA845Z774kDsh9bPcmoiyK8UnoBsYCKTK6LilWtvoDJEUx8fXXy10tSS81DG
I7EqnY27ZOf1LycKFJapR5uAxhSLKLLku8AuuRxO49MqfJhQsqGOIEwZdOLC/H0C
uQ7/SmzPCZYNwRT4dfiDnY6cLcEcEkhEogaY/2iiod5kXs4waah5VJU5h/hw6Zpb
ejeJms3iyJo8FjmL60uLH9A/iRY+qu98rAL8w09wGwXlJqFKU7Gz55wVDIKqaZwU
zwe3s3WaQimV14QcXBZj5yNOQwRL5EeudpTOFzSnRzwJ+0qVknfYTDS4HuoT8jso
48CHatnAEp/DNiQEVqoZnGIDiidnJe8rfvUQnFhM+JeZ9sRf23YhribvR1KVC8tm
TgIqV8gfJgDx7zY36OgGREbhDOCXlwH1dMA9kRj2nhMN0ZKg9PMKvgtu6OmBoxiF
BKbUZSkWNDNZo8SsY8ARMOhZnUydLcY+9819OE/Zkexyx1UNbmT70DFK+pj6v4E/
3m4MUQrEjFxnmTtztJhD9zhqKvFQC8A4xv7vy8IAzM2DACVcHvBGYU2P7WUquQBH
m5NtJaVCQftMN1SSRScpoUt85C012NamDO4jIlyu1uyDnzjk4QtYieECdJIk1/rx
0gRmTXBkJAnuZeO04hX8Y9PKylbtzSYfaP+EaNNUQTNXc3dmPVXmES5Dq5pZDAhQ
2WSk2Gs8T4cJW9vrDzjC+49pkE59hNr//472ZDCrBRz3rre7JuCAHjMg+Eh61vfI
Or8/YFI5vCpZ1Ussh3fIA4GtbX2Zm/TY6FRl0IfJ4CEd+V2bVV8Eu6rBbBfBM6oy
Ep/zUlJtmCjjp0dNRQQTtZFY4EHQ+K7Eyi8EhXBAmKCcew/lCFnYp5oI3oDZGU+c
zFZClhQzLGpV3ZabLzZ+1/NhwzeycOkVx8BQnxTr/OTdcSDjKnyHVDkUXG+NhQX3
FW5Rn542W0K48yvuXkQFrvHQAGyq6TjN/8Q2ixbqQagxIFfJouDV+6vuDAM/TCC2
ao8qnkY5kdxviMCsMnxEBSGhishc+pFaKAKmGab9SUBvDDWQqRnGznO2LXcZxzli
pfnuq8yYCVjLji1zkz4G68N3s3tZlMUyETHE3Y8Jov6WgLdNWILT7+rMlsWGYiJF
rY7hLWfy0yGT3b2bfShNJnE6UgR04mAND65j9gTHTnttXOy5dMrvsWF9qb/3jQsm
CRL+lL6TWRjcW6Q2tom4yMfb2GRpXOCXZ//cT1J4OYEsPHIRSReAxLoc6ZNPmsFu
vUf5PUIr1mChJd+KVBhBHgT9YcZXUDm3rPOnxtKecRazNnxkChfgcStFcfGcKAGL
UOJfujD/TgiLHOD3f52laFTKFYCjnuwyYZMMzBM7uIG7touS9Gorq1WwFloFyieW
dc1tckaScafIbFe1m/I3NLqtVOiThgT1HF5gJ6af7xY16Qo639Kn6WyCGW8W5dMD
H3Xy4Ca2clew2SHMQhU02I0kbpDSdJPrGdDSlzOUgAwq81MAIB6DFAmsL5MWc/UQ
9S6gYOgLROOyAjyAXxbb3CrlqtzrAnV1SToHTU2vtuwA7Dh8+9hEZ95qUAzpPA6C
+CsYRoaMXIkBqD/cBqQ2A7YOXjT/b+CGS3Bz4yq0htXNzjKk+aIrPnl/SuwQGnji
PoT7p94cM4T9QtXcNc6vJUzCPSOe078+Cji7tqEdqm6T/aD36xb5XdzBR7JRwuAX
0fBIpMwMqSbXkVxcvUB4paWv3m9nz29bvRoY3udMyqVgHUZIySx8e4I0xolG3P8s
hZgmmM3jJZVu3QAxh8TfWkyO65JcyADTxXKLaIAARynbySJHzxgQ/vFP3g4ZwzkW
JTSqWDtMDiC5GEIRJZFzGqLBVbmpNBIUfE47stNhoGqemajUnFjJdCt3RQseemij
qFUW/OhJJ03goCbkOBzM2RtkzhjZQ2OTFOIgMwNwth+h/LIVEfeuCGm04q/Y7EPb
W7qJiZz63OBp07D0Nw7kuUhZPqVCOUJXF+ScC5RJl3U0c920p0FuLlHYqwPhMm5/
I6w0D55xeDGxCQoeRJYP9Zg8XyLXeE4DL95LnfUHKyEWL7Acrse31RFE2G9q9RpQ
3V8zcOTiHhpnlJrZuux98XSK+c6Idp0FApPcJvkFYX+X5kKVKEmGdO/EvbGpl19G
XLv+JRD+v+FOz+zmXp3nTmfr250ocWB1uBCp0ft9uXHjV0dlUiEAxLjISEbHFJPV
hL5Bu3n+ixhR4Bth3yofcpbi+sHiYk2OeDxTOpTDMVdlJYljb2YmdAEonlVwou7r
7Mw+5PAFiY/2buv4ogHqLFJe3o1kadWhhu2ar2AFMyYpBLC2PyFW1WzRwxANV2TL
eYlrkO+qk6kBc61LgEoxzBiX33SjOewGeY7A25gQS82XIZijPVErMPFRL18oFpkc
YGTNDlQDKrL6ahhWdBE2OXb0aF5oMnecwt4D0KgP5mlWL9YQ0al6ZMlXHF1gUgVW
weicYdeCqOWTWRR/XXiH+cbtA3B7PjbRTBOnSmUqLbOSJUMzoKl8F850SDJkPMZx
Y2iTdFiTH/Fb9n+zPOjz2yYrw15T/jHjV7zDYII+3s8r2QlklkV4TPm1t7HZTM8g
cAMbLJHFigJgDiWFLPBtU/MSM3nPG+kxKuqSwsSE49eZj/oGpF1sODH2s217o4cF
2XLJpvx69x/lwtXIuo9AHXHiEzGgDIKA4sR5Q9vkkX4ceC1RGYqFqsWwp82C6Ebt
1HZ0Vo48Y1ipgn1z2gR2A2FfA2xnwhNtqrPrCZ2460WPNc5CR4Q0k80mi+rcNniT
Qn+/nLh9V5s6fWrmOyr1ZXlYlfBOw5xLDvEl5OiJ5HwDfVEz7ZbSGky6bL1lhATL
KgVkGfExSjTgzEGMvhQ01lBB2g/Xax2TaGi2qxJN7KCAWIk9CPvxr3BGqkUOqTCt
/N4zY6XFi8qM+0u4woCVQibwDL1GcXRkBre0ZwGTRApmOuCOIYd6fDPo5diy20Ii
1V/JPsy2Wkm1g/I9A8bQalBTKv/bPbQ0ygKerh1uR6rZTHeiy8NkOX2QucbhLUzW
skIrXhxYzEE15pPnHb64xrriOogT09FLxHLDVaNKPNM7QtAZnFpEyJ6RM+ypOCbm
Q86/40z6g2irOY9skfm0OGza57My6nkNr5oFjsvgBJmnjcW5iGNaV2GCxP7kxN3d
uCg7sCju3407c3mOBZ0adaryRT6d1haCtohiXdvY9MnB7PdKijOGTtQEdbj2239x
xo3DhkMDhURhUiVGSmsGbLhTEsrqYP/T3rRXf6ITwbQxomzQM/e+T1F3G5PZVryM
hEbxpIQveEub6NTAZ0YRhmD0VJ5QvWVYPePGST8qVsKNgM50Y4jXWfeo/VEJgUR/
OKHo4g5sUT1XKvkbOMDFvM/EhOaS8h8wyUhVAZ373/Ka0eIG6Nf4oaS9eETvmZaJ
xOPrTtut8QNM16COgkDY3IRAfvh2hzYK1NhatDaOHsfFEySxGB5LAp02idHQFT/w
zxbVYddCCooXfCjv1ZjdRCG4p144DkKWVKEBuWD4Nf3w8YbxQndZ4jMJTOqYYKrd
YHFsFlZn+P92lXC71UUjsZBD9OwC4fnJMT3G7BpPQFqRq2DXUuRqSLe6fN9zQuhr
aSZFXrP8SYEoiHmo0aQayoXgfxj3pV143Q0fLSg9ogITqU6oeouYSZm4GelO+ibd
iP+SVsmyqWpdRWQkbCH/zpLbSNyFw4vEPA8UQciZmAHSdXixbZEJBwVo+W94Sq4k
Zd8FvBOXYBhgErTJX4Lxbzljd962/8J4E0HrB0jVuaCo+i22TaJOiyPzfp4DkzQk
NYT5aTPc0HalrhMSpxjWdoHjJCd2MQdKu1zQr51NS9T2BEuf1i/vldd+Y61YEaez
9swwaXd1S1pqTzPNBLZ4CoBx9GWYyNrDj5VSWwfIiBo7QAK436AZRGsa4nF44cLb
oph6kRzjAMfzNuqW5pzuI4VYtInI6YuJDRZIojaWnuz32yOXPdZyF8vmXhzfM88o
8NG46+mo/heXg8m4RKwc0pUYiBsQf+HA8/Bh4vgZg+5vaZi0HTwWEA9I1esiKeXc
J6nUaecITFVXn+oydZmv7ByBIMdEk5lD3wN9/HkCO9kDmohhuKXNfQdqe1YCtDfa
47HA5pb/3t1jVuDF+PPjB6zSszIVvPabPsBJLQfXblSD9iRfdS77yayxuLx6IP70
mvlvhLBoQP4lQMf/oD7D2rkfy9uRgIW02DXby3qNNhejccsBa9KXTyX6e2rZUua9
/wFa7exXx+DLKDwA2DiA7RREvYNTI2ZAprxO1zDN4W9D9BQgjQIY4wyVUmNBPBVJ
3sjaaNMZ2plLyJmThsxV77i+K9JTaYuR3Owg6m5AQshpX7p/fwc1KSLjFdIycM3E
06tDXDS2qJwvGukHSO9kxu7/Slw2up0nCBUi0aOVlx881iuQUtOL/X1CVWaUQ4/q
2Zv9XmqirfgXbtCfRSMsjrGlFnr3BgS3Phj1xaObggX97PTPgO+zqv4wAH1Dqp0I
10/0ZxTZR8X3nNbm/9EMAUfB9cFbKbW4uHOj6gISxcp/UE+WbpHE8Zu31N6zScu4
uTxW8a6UHFxRBvArtMnCuETLMq3Kx2UBwyei739CbVQjgB76I0O0ZNswV3DRzT8d
yilpU/R/XHchUYBpV9mcMf/+ygJpL0K/WuaL2xQTNu6kPOE+hg7bA4AZdhI1iNfd
BmtdExZLn2Jj61Pj0pwcy++2oHeF/Qaz5royaKjI2IC5pxoOVWzMeF8IjSIe8xNm
062xKOQd3ngvZHw77WKmwZb5LnQBS1UOesfl50K+cuS0ab3IKxqXTQJ423xERADz
v8cYRPqvFD+0iV4HRs/TyOlnI2aQpnnZBHgSz3fWi83jfPwlVyG+kdd8/07R7IDm
0ddzuSwB1Tg/CELhghs3BJ6GJOpUXa81E9AtNhlgVjBcUqsLE7ZI3Gc0zGRK47Tx
+i1SOnYltiXjndH+5UroijiVwzXi8IwT8s4p5CX+E5x7EMXcs+fGLNXqecuXUiou
w9UnF3flI2mUSuKWodvzv1/fZ9hUWd9WqKs9RlVSOTb1TSUL4n4wMk9TrUS76ih5
e7g2ZL6fvW3SmTF7aaQdHquOwWey1qmvDfVJUVVopY6apqdH2OCn7C85bV0Kr/em
7mkP9EDN/R+LeDFRjFZvSzK1OljCGLwk6d2KY7cfwJNfhg1cbllCe42I1riyA9xA
gM0ok4+JfqWm+WCjKejXslKvKEZKJbDlX8xU2o3cDljDrieaUg6PkUr1yEFi6MLv
Uce907DErlRWkPF+S6zNNm/Y84tL58VF3+KOp6guQrJ+RFNqZvdB9/ZvqtK6Gj5U
PL8KW21YTFw04I1fxiBu5TmNITEvzJ4AJeGT4kUhfoUTWSlnKtmrXEl/8O7XKLvp
9UHn6wDF7jw2QzLeMsKd6aAJR/mg77DDQMR7JOo6ULijgymkQ/V5oWmFASdirNxI
tI5/VHNGzAOE0t2PtD89Jb50arflnlBYoxucVJI15YkYf3AaisO5+VuYDc+5h2Sf
chlmaSx5EoRnIkcdo8FHVlqoQbqOBkJYoGY6JeRIFMJYKMYKEHD/0WGYiNcNq8K1
FlB8Uou0M9sd3TCTw1II+FQI4KVnqgLed4/YhbFQtGcNZe0jDagbbh9swS/uHQ9V
BBGq1bAnfUOP1a5xSGz8E4Zm9Gzrg5lOzgpkt35d5vkMsRXqCxvw10yHqUuPCoiR
FdcVmReHTYdZAXSb2I1np0qACTO8oqNb243NcCRh6VfYUIBYqUZ3a2iDopYfeLlw
MtLyuNnxW+Sf3AzVdIMP72hqu7HsWm5mLScO4fu6szbso2dsMyJqk9rxDdJcYerX
H4M/IT0uKOVXURSrJbPFUYV2MLddR/hCpP8BwN9CfSr6RUrvJ6hrZd7XY6PWM3mN
+cifhEXQZqZH2HNiIUm5RyrwMxzzO53i9qpH0fl1ENAXkI4MM4oXkohfL++GnXXW
ang/hwc80cdRRg5nxItBTA+8WqJaTycFHbr/iWU026TiImIsCXn49/jQUreOkbpe
T1fQWOLJ/RpKrlS+p0pHMggwpzxwSufus4oWUQVRUYG188yfB1yyxFOVX8QI2HJ+
htKd85+rGScMK7zQIuxZoQJLVAmpvaZbrMCN5H3B38h0mhRsezubQnLRN+Y8DVuI
kDb9pCX1qttlSKm3XHme87T9piVK6XGyhIJGiLurMPmRV83d30vE3NaeZgF0YBu/
cEFTxkYsROjecv88cfllbfgsAUMD+44satrz7tBaVe1UmXz8Nok7Xsp0MlZdm5em
DXwxFOBhO8KBfCL8VUIQy+52oEUE4w8rQj/uoLlEHK997hwhI37Gnia8s7fZ3RTr
JaI0FZIgDDxilZcU1uAPHKhZ+LmR8YGCd0CxNKhyXCxuGI5h6Y5knB5+sGcUk9UH
r/oIXqMOoONTI8Wa0VWcX2Spt7y8UXg7KxOZ9dfVX2376ZxWOkCnFykBcCqA6cvn
jutdvtDm2LzBRtnDyLs9U1T8za9G8XNocrCM05q50xe+onDu5RDvqglwJh1FgpBo
h6M9duS59gZTB26ynyn+WkErFGm7QkdGyE6BVDnGaVSRUwOa6BSIz2eLQ7wKHd1e
PgaT5wjG1O01TDTOvCd1TQhHmU5WolilXZRR4JXU3FXaYeoCpgtQiRjz155xhP+h
41T+7oSZSwvWBbrTqsWqnmOz1tsf62eD2Gr86p7PT5F77hIwu+O9hryU/OsA1SpZ
oWYogbksBpJjelPDWpRgHaULDcJPdoYA2cWr65/zy33ZdOrD2fw4aod0ruAYy70d
m3KG/qObUiAn5OSP/mYBt45r4KTn0meELLkJJOy5yXbkCiAML3IYFNggzWMrXKYP
VY+ghChz34doFsIaQBqqwinpWKyoGDF2kHyygVrefQUjR+Qux4mkk0OIQ7oy0Ax/
aa6eVpxq9/LmTVajrFgCvRqjnpJd16UcNJ7fCugkXF3U9cpjL1GDf29oLiISTYEC
2E6Vvmy8SE7QUNIqjmMDzJ8wDknRswIrpMne3EF5D3bw2NDB3tuwWq8jnxuTu8R/
tagzK1t711B8H9KQbUJafJosuHGSLXIhES9dRJLYq2uB/oIVNd+IcW6klUyAGpdd
8JiR0wlSjEss9/svP4UGmgxV2Cz/gl9cEnK0YcqRlSOeKo+QVLcshkUwKy5LRAa5
ijRJ+2k7kylCclEWDUPwGP6CEkYMhd9EXbzHTc9W29ApQEJ8+I3S9neq+pK9g268
DYHi673W4FFkdLTkOMwRH9MIWKml9kI+qUVaCRXnEqbsooYSqXqDd0TylEAWPz7d
jSYurWGWKr0u6A90Qs1yJ8kwe1zHTSjJ5MJea1NWIH7tznfBK19+CPpCxDViOaWo
BJMssTfJ4i+Qf7NthHGVkuVjNLBw9TKvn/qLFHV83LW9aOb6FMSvv8sKHMf2EGux
/+nb+zW8mbdB8W7bwAdCqLR0fHBdPAiGAwMZ3/wc97zmG9cWf2jFkes6wGUinodp
QlCqTH6O7dmrSVOexWSk3LMPzbb4D6TfI5QGhd8OQRW1sK61y0UepBdjAXKVPTqq
4l4vepkMnGv4vdVRk0mhPV9waSOoExH2UBLPU8kdeoLoRhNOY8w2CsRv7o+vuPug
XwfIAZKWqcbItlkv5L5gw4KEpQmo0FA51dLcgOLXgnJwSDoeLYaZLp26w5OKH/IU
/+nMbu+v55YKaOAAzzmcFzM7qsf5r9zJwiG1KrmwgtGUDQR9T1k8N3xNQIhHDaBp
ISdivkx3gY44etOLLeZdngHmQy8kpb2qNQwTsM18Ayr9W7WciS8GwhaAKTIPc8rP
O5UAq+ZA07J/3mBW+gGr0IwKjgHU1M6x2iX8Cg5A1bTkQK4JaXZ3DKLy4s8omf8G
iO4zEabb1ZSTGRkVYVPyVtJeE2g/qH+XR+iUXhdXiqOZ5GcZtjx+rZDjwz21lEO/
cgMb9W/BhoFEePcToFO8kDvy+C+sZT1xcAJ3K/Tld16r7NnxWyYtS/cV0iY5LvoX
XIgttoyclHZ5PU36brusF+BwNUsoXerYMOHF6tIFzpASj3AhO0SGf6FUCRWwboPN
y9edIe/iAsiTa2zFiSNDdeJZyZGnnP3n58e8eyhjZoNv4X9qu8r8rH/Z0m/Y+ExW
RCsFO0zQiOuDVB6xbCz+DJPBc7N3SsVzDC5D++9QqikFvQt+Pn+uqLFNYK/TuBir
6eoEgC1LDVIqMmYCt0SeGJZRahXrJMPZhoODrwXGEnY4HNTc+0v4sNuZZmCRn0OR
I0XLTF1SjJsdZ5US4KRhgZENXmsGtDmJWMokRSnH7f7RuZRgN34ZQjOvXQJWWysZ
+WC+FHse15kBhfqJ+nmpeNvDVT/9j5OHoazbLIRGb9KLV0nhBhJL+9Yc44/4LeFh
kXJ7jrlZ/DO4jJPL3Lsd3xYJJ8nCWq1j/FY8cvUBS/+yRjOgUKL5jx4OZwIQUZQj
VmA/RRh+X5kEn+NuYQIgbGqY1sw66eAa+8YgoY0lgMp0H3DXhkveOvoeLdhedVf5
3hEo3ZlXNhh3+Enn9SGUbo5f/RjUcayg/r1ano9sCFn0VSFb3Pl1kolyEpB6zmD3
WOcsKe1M5Ybzww0KS9Rs/5zcoFPvNzXgbW448K0po3Fpp2hyFcpzvlW0xUJEhd7t
1H4BxDd72z2k01srriDAXEz/KoJ7C/kBFzhlC5FufP4ArkqrSc72j1ewIUM7CZUl
SKe618W+xbaUzICCy/FBKfQafFmcFQ41gO1GwQYqGXbFPNhdEmh0SCbtJ1gG+TcQ
5Lcuez1bs23vz/CCF/XJ02t7GNNf22XQD67KMIRpAdZczD7ODXZYyTO+9vTzuAMT
e41bv4tBh0Z3vSIb8c0Av2QiNP/xpQU9F5M92YwamJvsL3/4wiCb744TE5mhAFFw
GNexzlC3mRAB49Pxxi9CEUg3pg5QOgOnggrAzm1+GkP7If5a6l6mPqawhDZwoQhx
ikqlRzzG93JyczDGvUDLxoJ2uT+e0ykFnG24i1texpW1TAhkM9ICezbl5QzSMEym
tH0sCyJ13YT27JqWwoFWmQyrPVuqZvVlPiPfLvCFst3kksPQddxDUjy5KYUVze8Y
oIrAegJh+jD3+ogHaSOa4shXys8bd1Pys1AXtRly9G5+2pbHKsKp6Wid6jHvQ6Is
tFGXciAm+MG2CaTpXLHnxuauF1Xn2kY82yGnwkOLZ5Xpmt3ezPWTQ4K6XMfVA1yM
TlvcGCy9kAQam4y7yrUhGV3ry63xakRPBD1GIt84yW7daQhGZunrIC0T2YEzSahY
rh49FriwCqy2lirYFpEU2wuXXUDGVg2e+SO3z6Ah5gRKVm2SPEr+wv8rRiFKR8qM
S5W740hBxCZpPDLO4opuVphlK87Ksqgoh0R+BZN5qQXfvLsORSFq3nO8N9Y+5rxs
B1OOP9l6xAKYvvw2LJUZ05YBiJOZlc2/pumugGZX7GxhwIghO4yAERcbhpJXvFeJ
/FrCovKGx5BPOl1CLoIB+Plfz5uh+axMCE+Xt5M2qqCwqh6Njm0Am9g0/8EGqhnm
9VRTs+z6t2auLlwxG0JjPK8dTzEBRaYwYKvZ/TtVsvYdU8eUoBG2ajbAikH/u0v3
VIUjvwPgbK0mSHAo2WOT1yDmyfQ9HHMpDJi3IdHMt2fc6Z6CEUQLRWtzinCZA9fT
Rj03SY26+6XGXmYqswDV1nB8eAUfBoDPnbokTl68AGtrZmbhfnqnVHK6Ihk805wY
8qSDJUoY76/MzhDcODpZCJKim7Cj00GtFtaBS/UBVGF34d1S/libMEN7e+LXsCvr
w0ypK8ZVWGBsQYm2jqjN8FlyGA2AdsX5etepMzwc4HuFoPRLJNd5Ns9c5EH7a663
24xMI173vocfVthpIS3RTBgBKkV8IS2whi+YtjQ+ZjjPYiBL80t7VIQltn8C1xym
a+3dfpuEzz/6wlRHGbZSjGdso0CTe02XoZGPSR3I6RFXXRXJcY9deJ0eNT1oqI86
GCgiF8G4+mLJoVK2zsVQNAN9V9xwHAyl3HF6X9s1zGZg7/C0+4O9+uo4u+YIdXdB
1k2bLjPKmvgIBl7BAe000KVAsxqsHQttdkAo/b922dX99h/+NXqRnQ4yBtFG4tqw
7R646gbrVQVJmXoAm8JT8uiOIPTPrmgqo0O+U1RIGdlHQuFqMw4KxG7wqRSTgv+J
EyukYJhOM29pU2qHrrpXCdHhK11l0jJfH5C+nH87ALBCEwEPdr8q4hSuhifxumUE
mgeQt0A7bRzqBvoON3UBKOuWhUyPqqLv+p4maUQR+JhZbGVSP4hiI6mEvLmpxyh3
q2okkVgDigIgAnLDhTM+uybuj0NSFsXqGD/HOHEYxY3KaEFs59edFxZHTF9lCGRu
D+8Eo+xhuUcGYOHOgQz8+R/x62EhUFbEHdj2O6+CKGyRZtw6uNmDHDxq+polEHa0
Fj/TKc1/cg5hF5/uiLMq+pRlS6KwaRHx2tRa1cngJR1zWdheHXIUX+ovqbuzhQ/W
Ud8Pi2xZo0FbuyZQSIzs4Zu70uk1k8IYceOb5Ia7n0BBVaFEhzbBkbqmEHpm3HCq
HUBlDHZVOwQrpGOj72zPTwepUhXAc4t7Ncaz1hqC9o0nCp9VIBcCzAzcBHTrOlz8
qLUFS9HHOte31fzSdxzlKIgO2ZE+qjijzbCfZ43po03qmmybIVNgNs5rOnaXn0g1
wdGND5EOcBQHiHvriDCdsqd13dE0RFH1nMRU7kDxUaQ4q4Yz36jrniD12BVdLLvX
u2P3Onc3yrLU6uDd0zahSpRS+uXAXnwWX8eCgd/M4sGtfWtmPbxCfp+w78xGmMrM
LHMCL54kAZbu7AzMgbTDztDGRZTVR7ZNIWJqn+CuQsIaZKBdSqomG48FtmGGR4nd
ch2POifXkUsfHc3AKg96xpN13fvRloMBIYYow5coNKeTm3BovgaEUNA4qEooVBGl
EcSX9iIh6UhmDeiENzo6FwdlZZHkMSK/vI+G4bwqbOs80Hopk4H6WAKLL+HlfUw5
5nG2MjE1uUV6DQF7Wiixct5HPYOozRcko8ZJm2u/XBRgIa3hC9g+QCWH+ghNrMf4
aid/BOyGqnsPcvFgAONnzk/nW3PM1j49LT8Xc567l/+IIeYewalJ+eI9npb6LgdA
+Mtyhi2ApRaIekNZ6xZtOHQtXdxoe1CVBEXmWDsUdCj0zgQe30cILWpfi68giPnN
jrBW6kgsbu40JGLJA7McRA==
`pragma protect end_protected
