// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:21:30 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
KycDs9gXO1FetPVchHV360LLFNhOd7ma5E1Ws7GljTYEMfYFeHgbrn18WrwR8wWq
hFdoCG18Pn+xLEKLkAWzemF19s3hJNbKQkFzY/RMW62QFVZgitvCfQnBv8r3Jm2P
ZWfdhTcF+xrv2NpKOnGkWa6hzplgK+CgmHft41IhMy0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3200)
G1uv2fj5mvRYoB7YqKorLY25LG8yJVuF4MDVlXlPnkC5p9a41+AHhO5pULelrm2O
s51bcBz4DcgQJfs7hrU+txIAgDv/IuiFrtlywmFuiEwB2DFZ3VV9LNv9ZchkfCZ6
lQ3wCq+3CbUXr9n0+9Mee6kGrmOtDhAa+ViJUyJH0P75kzKoNT6b+VG/xHQId5T/
kMocjp9/dZidYmfL9aIpbDIM9AYmFngN0sCnoqAi94nvBjOB//ZFUrkUs/nroJWQ
+Jw3NrAI+/OqR7z9IIQafWofyuYssGfgirN2bWh9+LQBWb9QKmu473KKCzSYwUV9
l1WBvggvBxn8Mb1zjT17kRVVNNQoZgX+6BhgEWDlMcRM09FxHTBHEqMW6g14naBc
hZ+q3sn89V420zRaC2G6LrxVpa/XETWP8baOdYo7OrlukM+8jS02qZ7gtaGVHppV
05UQObXsxU6yrYzoWwk/BleuCi7Rp3UtymQRFjRq/hwBQoYafP70dlMnLY/mgK/3
0n8SqQdMVnJ167jMlspRVGWSqZ0bLRyRM+jStPLDmiSQZjjDIHadgFxEsz5G2li+
8QkqTyRLybwQHjJ1BnNv2aTlrkHJqykWCXnBbcJs//2d86v7/3hhh2BhKoMSksXU
cKc3A762ralE93SPpLGhqSA280mQHhaQ4DvK/PEAdmu5UYG/DTzUcfZnih4YR/SF
g8x0mImsQ++/PLFn3pf7OEScsr/NWp7bLHKUJe8BpY5NrwcqkZPAU1e8Uec1WMY9
lxj29XTIBv6zYyiOp1AvwP6okib+f/G3WWf60rFDPGC1nkU4wcdKu08G8xra6215
REYHqPXIDSQPN3pqesUQqoNFxCXp0IcAPjrf2m3hEddZ18UIgYG4IJomOPimjOwy
ouJ88Tb91XswsM1RqOCWDJY3baLjyZ0ILMwOcFH9RGblwihLRwZcG8FSd5HMzFng
S3NRuc2NC+jjEAaCIsmWHJa3jzxDZ61kFMQkaX6kxzyFCgnjkHeTne3iEHU56TfP
ianeQk++woFdPEURnsfXfsPY9/FNdj2aFwZV/Sxg++IMEKdVc9TAk8xq6ZGFJdS/
pJsYJnaer4BV9lT9p735ZGUqcDc023Ezp7Zc5V/xlLZ0JscaN3w9q133pnlk9AWx
gsPzFPjy5nlMfwPWSBxdb7QJNlUNnPdfsyEznZ9s9IiME3Dxg+wM5gfpzlS++hKW
oVHqeGgPb2DC8jyDH+2dEM6Ze6TWDZz5r0uF51qTFBPUkX8Ddr1z9wAboAqhwX12
NlmSrgT17RkjDBxBOfVNcdbNEYGr0T0Ic/yFzJ+ZApJUmJgn0lwdAsuCNlSELCMq
0OKQ66Q8BKoMVqHkGmB21UJBm7KWBWjiEdrQWJ/9vQGUXbY+EL8JfE8d8yw/DOm6
3ce+ZmXCPvDRcVdTKnZ8MECaT3y7gtBFO2WNG4gmgF/tEcgyegVLBrvGo3pSYff3
+DbiOC8Q2LThdKocmu9nmbK/lHlUfGrSxFg8OyeljQLkX64Ppu5RErlTlLHVALGt
Rk2QfXGZ+RabMgTFZ/q/amMfZ6377yTtsCS6aKobQDytsBPZEBElyDw4xU0Cci/C
HpwP8znntQquiBLITfTWxC7GAd4xdN4bDpRVVz1ajsvJPKcYmBKYuLg1lROHI+3/
Ih5xbsTJxgn9Anf5kxoblChpW5TlVQMa/LM2WWkEOYEmVc1WsDLKgN5XTXUUDvT4
0SgQBhCrzPa2xgU0nngepc2rXK9To1mL5Yvu5Q8Xj/9tjZ+nWO0IJKwnKQoRq08V
Y1ECPBDWf0aCsSHQOs9lTp5RnTzK5oz5kRyk5W5fUVSBhe655HQH7MEtgZaD+G1X
UAl3zcyjbOM++HsJ0HN1x1Xl02ZzS8Ed709rjHpk4rPGNJgFxHjihKKrB9M0bo3D
P8cE5dIO0aPYS2Oc8qfCsSY45Z5RRK2scPuZsL8VkyPannPrgQY+z4olarF7mjXN
LGTv42GI2w7YZD+x3MK2r24fi7sCOwuKugjfyNzX6LHfd2NxGLRGk5b4SpeWVdhL
5LZfc24AeBeLBUcJoeUDQANtjEr6wUifpSWRxnFKhHpEbSaPu0fvmRVtxlgxGOds
LZjkzNhzxfeA3uvltq7NUKMpdtixQZIyFnX8NPuO9iRMX0mpdkZ1u7MxaMGDBOI1
kn0nstA+NB/7imYquVHNyqXA3nIgd1LnxHtboU7/r4SfmIln2Ef1BibE2tZMDs5X
rLnMbwjWaHViQHcSPt0KCZtMEfLXLJk/hNODH1Wbu7kGQLgfX0xKlviYtZM0WU56
/FZ9omtDB1fN8vZBJ3eQi0daAQmNaw1B7hg0wUFqrmuVjaxqgAKiefPXiTkS/vz4
yBsPfA7fMMDp3wl3GaaB26mx63AAqNlMQwK36M3jYpPkpMQ6D09POaRTcOsj4o4f
ADi5VnKHlcNLvv641dta/XzK4hkaURBVK25NJ6ovrv0TKCRNdwlKcjB9oja2mgcq
4p+xtM9MqEwEkNODiX/tOUvKsjbimMl4dVGO2Zq1yRnalofb6Lrer07zjNsddh+x
uMXcuYZv3IP708jXKPechUpSI85dio7vQTwIzwDtVW8m252Gu3LRDEGxah1D21zj
pYrV2vwaKVbTj3PfZnjg+RhmW0rK4mFHkzkhVruQuRfhPVWTzeBRsabV8tw/WaZf
luWBvXpC9mqS2ZjAVtT4KNbDd0tkJgzd/dky7Zr9w3AvFnEAO93+PBjaJzC6U9Hv
whrmdBpAxcHu3oGAp6LbiYU9QrWwMGOp7BOw+9IDIbOJPQtBqiypNsK5QZ2W0igo
zOfB06Y2g5FnZsjLu1ZC04Sv/ryPWnMrK3ZEXA9+iqFaSntfWKl6+G2zgtF6n+Ck
GcF3JrvSrUSHJGTQcMmIakOKAtmBGRY2sbJ5KRLuhBhLSD5QwPinEB+ezEiXaGA5
yqIpXFiheMdvYksQg2iNHb/Zq/E/rXosZF9skA5rKK3M+wwR2FD0zsuxrTP0c7dy
/OLy/2PjTNUExFGVr1pzGKyenofKqUjXy+YBZaqJq2xHwInMtz+iHW2uGTToEJqK
xfgFCgi5nTPxRiFY2r4DZZ5vP4tqjFk019nv4tPnxhsB8P0RLvIhZ5tS07YydQEI
pXYlicRzsxc25+sVMP9/g8JxaLH7C6T3w0O0/WSQnc7PFjhjdJWdM+vlVuKOjVGK
dw+Cf3VV97FUT8a9Bz7xxicDwv968iPXdIrfgpdbFRKOnfhrhH+DGwDrs/IGYb9/
vyMw4YV9ALNEJkGKTem9d6pcWN3eLn8mZaEy6ut/Deg+nWOo6LmKlT3F8mZ6Z9CL
NM0VXbWjM1/+sM/zaOJhFu0/vl0zmi8qW1udzIO9OlvcX/RFXkLHWy5vMcFfsNLT
G6R4y0ldi+VdF/ovc4LSmOHmLqoRINAiIWF+pQPRKNghnpvd/h0OJtFj8Js3weVg
LD+EWozcsvSPMkdVDCH0Ak67jbys3Q1WAFodoSKKIVm3XlAwbyBzRbI2iOLqaQCD
UmX0utcCLNCbJVg43Bz9FTi8AMOdCvIGdzL0P1Jm9iboyrOoZKR7gRnA9bWEd2Im
UsuwSjdilO+QwAoD3p/0r4FTfoXTg0cZstb8f07K6y+b79tj+8i7cjQG9VYOF0A0
CFHdY2Q67VUyEMxryJCU4bVUTerCQS9nQCxYh6zZyqtVpmYpItsWpk3RWGEetj29
vqjw8nRb3nfM54gEsl3zvZEaO0wfdqk91wyo58UrHEr+mlX1UmrzuBoET44iIJKw
AU3B8+5NXfLUFGx5bLM/ebRpIkXrwFF59FOptQBonFY4rl3lGzDzzd+uPrwAKVbC
HKI/3va6DGSC7eFj///znZSxJort8w3MfwJEMx220zOAFqMaHIhj0TOFy5BawILx
juwGbWljgyMKFIY2BZEaSUM8DpgfwCWQsCb1srnixPf6gF0nrI2pGTokNdrEvaS5
gzfYbkpgW5QdAaoyTiEyDTvTAD+aGHPL++WmPeblIzy9AA6nN0J7LBPk+XY1zEPs
RqefSIVcL4a+pA6lDZ4AHRBcxnwDmGN99Wup69W1G19/wVMvxSVHlCGyPv/9+Axg
ophd6iMSORx63cjgIfshLz/gvGgwAK5JamIeaGLZiEy2huxvH9/R3mgPivxVeP/d
ZboFMvwRANzWrQ2pp/esCF53sna+yjwLPVVAkOJhaOdJVjq/3k9mO+vdBPBTqYgc
ERCNwN8gEFdI1mwloP2CI1CPKWRiRJA2s0YJS6kgdiY=
`pragma protect end_protected
