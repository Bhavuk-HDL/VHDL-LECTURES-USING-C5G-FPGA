// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:21:37 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fwI5/SOye5s6uewDhYNfIDz4eBeuDsW8hU7zU1ywQ5epnfIwd7epL7kdC0/0DQqz
625Va//MTSU9b3GMjLNd2r/RnOltY40vRaUfAOzku/WfRuU3CYZwlCJ7xINygjzd
zPF5Bfm0OeIJFNsAbvz3zOT/KqrBPrb4ZpN+nizgru4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 184976)
gqniBYNGdBZUl7RrSvNtVBAo176eRETd4iJG+SjAIdjm+VY2dL6t+4yn5lcUt5MH
p/wIL15bkLolZBw0k5G/2Fa9GywrMshQ96M8bzujwaqpxMAL7ZvKFpJv9CBY7OOp
tTfY/IXd/AWQmS3y7dGM5Qu3HWxT7t1mWc6fcdb+/lcm2GjAQKDE2JSSxTnsxJxW
Eix4BGQkePyX99EwqOcmVfz4V8RPqvGwiMPaVqZbm1cc6K4I8a80Hb8QRRt4oL6x
1Zj57L1dbPFg7oztQUXjjcZz8/pfisJyUmYSsQpxeL0KO+0YB3UIuQbU76B/fAMB
c/QB8AxPUjhXFlezwVtIKdzWbtjUhNXCWsoVKs403xhiLBMb5LAckYL+p/Lktt+B
YnLyeUsdnPUHWqdALiChDn4CMATWerykxhsuhG0q2mg/i2cZYB7966eIdyT42Wd2
Y/aKUx/OvfvuoaxkuhkMMqRB/9TGityjVxV9i8chmRu8blvT0s9c0tU0s3UGqJ32
oWizsb0eZipOrxYfB4KLN3rVtKU4HDwTCJ8bwTiWFAgVqlJxHSVG5xDLI95hmLbf
w78J626M7N30FojL9Rts5Vaut4hnp9UAYx5tyIbuTr9+tH8ktjFlo82k5EvaqMN6
gL8109xsabVrwLZnBF2TWKQ3rdG9oDEQ+hlQPs5W73pSgWmeaKl9IzaYNlqc9TIK
yRrEp4sQ8ZstfcKr1PlJ0mdTMvXcuSp567dx1KIc5fPd52xzm+UslKFcwAvy+5Iy
3CAT0fOGwKcKUHqisviJDqHUUx1DTFmA8rKJ3InWYNNRYQlWg6unAtkZWEkCH34v
iH2n5TOd2pc2EieCYaaIiTm6fASYjO0fq+Ld5opsAdYfPA8bmTXTyjT9vGPCdt4p
+23RG1O7TXdb9kJcV1UXcYr29MKj2ftP5zM2tB10nMYgIoo3ZjsRhIp/r/Mi9LpW
1N3L5yQDknEf+TkgyRqpu1BZDTVvQcrnB+CYZmAXLrQ5MNvsG5T9Si16vsvyhevW
aojfZ4JtZQSx6zZireB9r2uZjuIQMQQ7cdvQpWUwM9VFgEkZVJElcEkhfaT2tJwR
BWVGIWU5Rd8I+isf5NaXSFC43FgSONR7QtYs8WKXihzX+FAEUNVz9dF+6AXB8oG0
qGIpVWlu6vNMrhgpVxxLPE0nqGCQwzptVNc9ejSVY+OFOMwA9ki5t3tRhvAWahG5
WgyhV48bt29m0q6/nRX2LNpCkCPHHvoWt8bj5T2wwNsrWFazLMGx/zz1hI+PX35t
pzLGxD5AsCB9ILcgirKH/zaQnHreX0CH1QRuyB8q6j9ox+U/gMWnLOKBeK7jekq0
wPtVi0fcQk1lVK4JWADrKCHoDH4Ws9cLqqU8/A2dLS4L/vqrnOQfbrzXX0bytSMq
RZ7hAoeAP9RDryPWuCnZpiM8w4nFW1O/+9+D4ThEwbWyJOXE90KdPMBQ9A1wnPhU
aaesS6dHxYe3GVYMkE5umMVvhBAFpl8NlJ93/F/6Rfmw+tngHSAVf+LtQxrVwsED
oAEnZuNjUDuTn6RuXK4ZbRTGYkMoMIhvHv8Ip5A/+9nkKRrLzN615dwGsaBXfy4U
T+dg99tK4NTtLU8wdjPpTSC1vfu/eusyac1rYsg0eWa080GJT2+SoIjQ6d2w4+SY
4RXyXpgp4qgNtXzcNiOhHDCvhM43s8ODHz5DYnYme2KAeFJSgWWpfa3mAXcTStJc
v0C9bFs0N5ImYSJm4AhMnUSwMwZd5CiK5Q/IdKpc9XdY6lSEwduIXziUw9jES3uQ
DQZeCPyZtYO5NqBp3OitoI38NiI7dmsgyQNEwJancWDJ23Ur3G5Z5YBBuoS/uRKk
qyotWU/UDh5243fhivrFP9Cvfq7QVZzQePh46NdlHUjCOXrSW2F4EXQwrayqL8hX
ziirMke4//jN7vDBEC6Gjym7aQw82BwTWKUSuge8EfksDjcCzGcswjSYzAjKtDJE
lq9EvZTxxy9l/+DYuzECqsGM7CyEK5AE/yJg6eu88fTi5PSj7kquz0rNt5DtCubF
nwUYrgPqQ4UVtbPFZqEKb46cHeMih+e1BRijb6mnrLsOptA8fsXgT9WKx2pnmkua
p+/SDOFISCG9WPoIIAWYWwG5cMK+3j/enIHYhSwI/d1dRM84AI/IFP8V6sXPz/5D
M1OOWxRuTc48UZOnnwYgaS4UVWeOy+FHtw8KfaGbaNH5qA+4sIiJ7GG+I6LcPB4c
jFxPj5PzZ+Dhe5Y6t+u6zKGaDJUgIm4gGaJdp4EAuffsUMYsywljKC6HBgSx/nsL
Uc8KYeCVudtG6oJP27wjbbFgDhAR/alWT1QL9lrWbUXOL2Lq6AVNrDTlp6vXYg75
11IzfE5p3EBW7HMLN5UWZF1eBpkcgAQ8TSRa5fx0/dnY9BWBHzy6NL+Y5q0W7q32
OzcdtcoE/WXCRIYsiBeP/wjVL41EKIDTJXXH3zXxIYSym116JyKhpqSBmygrIvxR
Aih3bpwNDp6ZMjk4gwGWe/cWXNn9IMSmoU6dgpPce+Bth1nZS6Xipb8/JeA/YR1x
LjY8Ge8FwKRw0g5gdQIS2WOS6Ziuwuws3R49dryFTRy2MAgGt4cR5r6Y6GPj9oyO
Rb8RLGE8fyYVBZhMPkpVRaZ0qoP+J7BvuhwkmhajkUGTrsiD1JkLlClLOjk3sOB3
wkQul7Q+m4iAubASjjX7o6dfS99tkKY2+1A8A1tIgtyrkFYmvSx0Nm9tcuZrHR4e
YyJ6cRpcWE7Y9rJM4l5vnzKQ7gwiL0jOcNgSu4+OKCLYbTmRAtmBJEF4gimn9Ffm
TvG+6OKx50UBggOXtWxD0O516yYRLDgQKKZXgfRRrB0RQJBhu4WXbkNY0/a/u9GX
NCEMFtvfkqvFwHDU7HaDfC++bn0bJDxjo37dzwdKEuu3A5WG1Sg39fhDmsERupBt
72K1vesgCUGvCsVhdA7maPDm0I4zkXUFwf5TbEV4NGX4bDYk29e8vakLwsAnUDPe
0y9vWjORTF23rU9esxzVG+vpPPzXEXjy6QDWl2Bp04nbmhzivOfG11ICGqfjojEt
ehxKhtKUZuJEL9/Wz+sxgZ7AYrrnBqUocPAq9gyq5v1FlHzfkhFUe00k6ywAaBWa
zaupO0aDxpM/h1Bl9ruF1DlEfRDXf0aoEuArSd3Lw173YquaAhu3wozchAtVMKBc
LBWVC+L9ZTn8c9hpZdXC5p78V9JCEeoGXIQjYXLzsKR6XbztsssTWObSeMP+vpyI
tWRNxHI7Et7OLBkBB8CAH1JOTbkGT1Te7zXJ7AuwX3inV39/mdacHLNCMkBF+wSS
ptpngqLkGWrmHHpbEYVEhh//s6IcVZjibINMprWr930Dh6zM+7Nt5H+81gySvZWM
QTSZeUpHL6nJh466IKyY6wDCWb4L79N+wRRg4BPjVq7f4GhGfCpts34jjW2adSZy
R0bG0LJBXVHFdNRdkgMtL61FdHfP3lhoEhS7NveVoC7SgOmG0MaazC0V9dqJxVtm
5VoLmGnTaZ0KrXnMnv75LFfGsViAMwDksY8a6pv7mADBkYj8zapwPCfloftlzhgg
WshGSfeQXR8L9f9P5LRK85tfSziv0ThbTNz4ftiItk9bZpWbv1skIfFsumU8q+VC
cKqVbnLb6FBqVZGbHtbBcjXW12rs07LElRgy5CJnFk+VB9emuccu5bgIijlymtZt
GgOpJKLcFVjxwBy5uNYtSMrgfEF8rO1lqA07oZLdIIUXM3OOATJ5H3TOg8egq+gY
iik1T+Ul/laqx/PaMO0w7zluGE2h8e4jXAaXhJKUUzoZpVvp6pgWOi8OnVdhtnMx
ZS/X2LMaKfHczRUuAuyQjzd3nhh8OQA+ddcBz/bfut4X08nuHXaGM/l3o6tKBBuc
o217nelhxMQCd7DJNrL/IDUdnWxARtKDiABfYdbzH0tWjI4PkVvpstjZKGS9xLOC
6j0cejtdPx9fXFdLBwad7rq6UFJWixJzd+VNcdAvTAZ+OhoVolyHDD8ho+xvpLtA
L24YjgM+tT4foFacJYzCI84+Aiqx3SJAbFiN7x2uCwkrh55qT5Fos/ytclGc44tJ
xB+YlihJ1IDgqnxdg6uhj6JWzL1OPV7YSwb+QwM0KU4dkwh9p6DHMTAuIapj0gDD
+yYurk7GqTABoiMVgH8+uu/8WLFIoIGAv9HeY7+1+t/TkZhf+4DBIanJKy+TPtj0
zUhca4Ne1vkFJaUkcA33CMBdhTv2t0eaF5BWdGAapuP2Yc+fI/fMF8/8kXwEsMC6
nEww5P03eYwyMQrnQ1ohh+LrtV4EO92y6TaTMLknn+0/lBMfVORTj9MXhPhjLaV4
yI4nMTIxrVjiYdlWMxnhJo68PEY0curorYTBy+6VfUh78qcCKzJ19m2luGVNv7FN
ui8ajhobRxotpe4pQ7CqD32izxKfYYvp0/OX08A1oebd6T5mWgxvumacMgGOxdqj
N600V1Ic4UnW8toI49jOt6tEYNGafd3ovv3qu+NAVnFRyZRb+mnISsDumfHyYS1b
9Si33EvcsuBAX1xhfFtCH55tmoj+Wn6GkRtFAgguShJuz+/Hr053nhlcCqyXPWbk
sQYgnly4E5/Tp5K3p0ncTBjrwAZPXMKTY0y3HDXQthTYr1bFlEgI9yROVYuqW9Om
4YG1wpY1G/dFHyZL99rHTWvOnoAe1swi9crdPo+u2yhO+PxQYWwjMlqShnjbq+gn
4+OTdK3QdxqbDsGp0wAdFrxAHQCs339XhKlSBLcB++VaL+oeBeOvageAlGEWiyNJ
JChTNxJ24rHHTyGbAMpGGh2l44ixNz3qZ20r5BP9JkQ/tc9RzyDyqvXFAm7txqtO
ERH2dUjqHd+oeGCsBoyoxRFpHmrosPGKCxYBq4/JkDI/CMV2ziDYXs9Q5IcapR9v
fiDxUe5MtbjmfxS2X4a2hwcE8MPQoxj9Wa6M6rKma93wWJjRAvdbwd/iLTikUPej
G1hgc40ITWj9fQ7JiB6L+cnPd9XsD0kVjOnvwQPDdm41RYJXPkA+2Fmn5/3bSrIn
8HUjnfkfSUpruzmbYfVXDgubAo5bywwe1iX6jYnERZOERZ5+pUJOTucq2ucBbJ2C
wy2kOvBu6X/X7C5DBEc7A0gz7XZ4iw/0cMzlCn5/yCF062JiWEAepaV6/1r4cEfz
F8wj3bEmknKWqdRruKB/XGTB1bOfGhAo6bLXkmzFfe0YZV6MGcEaa4vu30OAOmqQ
p1fyGnPtrFfGNcGq/UpS+x7TLQyiy2Ak5WZHjs6R6h57XB8znGFwqBwLpLJQyr/x
jIS1YZe04wmpVsGT6GzFW4562FZWDjoEOM4t4+JNM4x/GkqXvaeJeC5p5Q/4t5a2
PEovUvjXdZ+YHelCzAG85W/8dVvFELkb3ogQqR/RE6chBZWVD0yiASJAcB1rXt3r
VZ9UBnjzHo5XP77ru3xiQMKygMUDf3sNOEDPV5MIAa6FjZJOAHL71FO9VKoe6gbK
j5qJV/JDVffq+zdtTiXfYTOd4xSTbI1UPmtr2tcMSK77ItrrjDG1e6VaKR0mDJMR
RUpZmcfTOGs9+1eRahYQXhP45a3gs/wixE0jKgFOVBjkeizpaxNbeXii+ZZ3ldCJ
aGfTNVQvqerttDPxLfNinrZ2aIhHWzPShPKCHDSrh5zXSwunPwUe6WHZaExj6NHd
GTwyHP9dRyPFCwEPwoj/1AwgpRo0Dk+QHW/hOUA5q1KNE0hifzrMfkCl9srg7Tbx
bBXcoY/6TNGf+EDv7Iz+CkJ6SVuCUiJgpA0HFNT5pfFuMnq6JX8N5CtlfSI0H9Y+
r33lT2Iy4IDdM13M7h9KcFQMK5OcD5tCKawXGMvwY2WIGqkEnVisDB2lB1etgLul
TgtWO/wNdAYtcRbYoK4X/BLplPmwr78O3GrSgyd5z8D3D1poq1hFeUWpII3lDnJr
foRGgWpm+icEq9UNk84cAl/8Dnq0dd1XJ9ACEFD710GhLYyJj8wyflZ+XgJpz2/K
JNVPj7MOrZpNac4zHnNakLUuKqhMIRgXX4Ii5LdMhIXxE7mCjzjVS6YIIDT2sdGB
jin9js2QENAD61CxRK8zZFjeukzldsRrsLDys3hDXDu6uNJyao0QaRJUPVuWVacf
chclsbDk/z+1Kq5z8zp3WAc8Lih44FW0rlfKv9GSYndNtXKE79dDIRT4VLJ/hlmY
rEneBwGkydXjwiNQcvGnnZpJjYlEsiO0/g6/dqj0+pCmZABwP0g87Z7G7K6e20hN
77IFlOY7+yyLFNTNrZTeY/BbwboL7iESeeelimDGb/9vp6sUie4JyLgcGbL/QtQJ
rzYPW4Uu2JsPic+bjoaghsildbjHwBjP6qwqcTQo8dpTChrJkeOVwnRYXvXBzZ7n
sQtZETFsYljxY8prlyn8AcLWHAwxcbdRF8wKVjikzBHtRAln58bFdEHDiOXHJkLM
qHJDOQKeT0db227TuQBe3OFtvfRzbB/PT9Zs0481QuLw5/nP7vdy/kvbI1a5x0r5
3zLDH8qgoabLGRH5ozX5t5dGDnIMI7518ziVLkWvt7Eppb07ClLJiLxp4IiJzEHG
qbpGf4vZ3BwwcYStjPpKZvGwznUWVX1nBQwtsHabI7fH0Sou14l/CXuyARr7Fjf2
ZOiJNapms0ALoBtXGakBl7TuBBhM/AjyUa8Oz4eqWP3NqadZDFtGlW+bycbewEeh
E6omqpGqh5hfe2zwM0DXvSJxCCBUw2+29w2iNYVHiBwXBapheBn7tv9xxHDyhD3d
dPKy3S0zXh8j03bEclDwlTUF8z95tzLm5Pk/p0sSlTiTpurq6rooNNRUAzfo1RZH
kSY26qJKY0SlMxrckwJeD7q51H5elGTFNl3nDWMvmHV5UhZ/RcbZHDc7zgRzSNWN
oPwssoId3aoLINMGv2ZMwULDYPYijOV5CKwv78JqFOONIiWoCmYyOL6QTG9ip7aT
UXgiWAi78+lpAM9PUE5cw+CugPEt5Yyfrlmtx/fn87LoBswpjFogBT//AWlZ0cr/
+BfqCZQd7KSmPjaYIIyV4eI08YP51JkX8iJTJLENvnYZQz+Zx4vRL5fe9Hr9CgYj
yy/m35bMXMXw8oYe2chJmEeOuuE9priwP9wIZyQO4CAtkOkyS6KRIUlSFOE+00/7
nqsPtawvFjLFUUU9qtiOD7L7LCDeTPvn+uJYJK0ILts93DWbjPcFMW9BoBCORLIA
ynVYRGOzwfvPUDkrNvBYrmEWizkbxHO2nxx3XWSCZAaroTEw4pp3oagzbNDXN4K4
rvjmI87E56l09hQrvjBVpwPH6eSL2V6/o9nI2iI2j4VuIW2wvNoPZHi5aqRSinDJ
Z3fFDah/GXAWoq4bhN/txYHW3B4V/5dlNusk/lTtEAZuE8KrsRgb8yJAdhhfsmxk
T+qO7wjqxZ0ItTlBVNh66TtwppsKa2PZqijrotWX5MjJ5I3UQXXyApe9ZY/SYjO9
T/u9DhE0OPKdg9cqvxV2MY1wXaDE8S0pbAVlcZg3Tn4TPt6fhRxde9yvVzcXVKdq
WN83Blij1scoVh7vHQ2rteZgDmeiK82NyPrMWmfYadL9967PB0cW7g6Lre4nwSX0
bSODOFuKCUvhDzAH5M8EU+YIWqigVZKpi05pNdexCY2vOzcM9nnvnweijyislxcY
EZvjLFL7/mSla3m4sUYRZeT9uVG4eqkBMvcjTyUZoG3ZiSY4zYXRaZECzgmvKkEB
uXozMaO7V8fiXJAs/H85TuZ2Q4CKCBv/gknKE4V7AmfoABFY1+kZ+zQVW8XJAsXV
qEXfOnHXvr25bMhrQ0qhxzIVhD34uE1PHKlz6jn9e75YNiokSQDO7zUS+PQTJqhR
VSOjQwtW358HGF0GzC0wbZBzJbbnAOqaKg37TexXQxPQ0IiMF+ekPU+Dp0Znat8G
Ei9I+6dYqUiTH9hKQyW/kCgCAMUex6iyfywOYAta8CRJrtUvw7SeGVhjOQMtR4by
SFoueaZt+OlnkmlZ0hlXNQ40Cfykrjk1O1kn37hBRzsBPbONCbrGHgAVm/Gu6oA/
KCsjMn8w7MB9K2clYZTkYEmls+ozTApiAax4EDoP5U8BMxFu/Ky6qSZL2av6tali
bOV0s4dP4m9bUpAVF6ugMOAXSlIxar2gcBIJJgVWqeUptZiwSitCmEwkKUqaqPuT
hw+F2GHDhKh6FBqvCMZ+A48p9HVCipbGtYocQgO25P27Ot7Alu8K+ajCLaGsWJi0
RuBE9iIKCVPeb2cmhBteLw985tMfX+O/3Iig4MBWMrjUXKfoNWyH5DpvW/mu4adA
vs0+e3bIQIhz/Qh0A4eP7krnrjNVnFlMYkCFIZvN/T1rdZZgJKLinqjcRJyLCnTb
1j7rQ5Pd2ybsonukca0DFVnFH2tFzL/gYcmknDcBR+VPbBGMNFmF+4kdbTHlYhZu
CtiUtZQjBHEVuyi8l8BJViOSBCaKuFFjIUt57MNGE6oP1W/XTdVrN99Bi+M2/86g
QEoyMNakX1olkUjMJZ4wWtWHIBTEW48CeigQ/GKo73E0UGEZvLRfiNmUBvvpFrGL
w3lhWbZcJ70gKY7OuxNEzoZhItukpfviXlOjojbBakWzp7/UDc729hHTRIZYfsEJ
nwGGCArSbWNKCUpdQSCPfafUOVgjfo2hK2R6FemuKl6SE49F4ZvBWPzKfJsVSqYc
9kFuyENLawzOs6SmjunjJXaulx5GsK6c86aq6Sb8fZ18iNBAW7xONBLR/1fLhtGE
ltnVaXlB31VqF0aAkZBxIDnCau9QY3YGaLhhUai8SqDqZzUoqTNx43YL+K1nx4tr
qbC69QTbm9i6eg2zbOgTCD/IeFqG0RQqOLsF0O/dLtQ8VsdsyY1FwNJvnrFi00Yh
DrYHkk5kk6JZNPtqTaC/7VDke8r+sSRSJYe9E6a7k60Yg2hjN3nUYBasgaVDJM0y
fQHRSsuvRq2+7YBKz2UbM+rSEhr5XSL2Pib/ZcTM/sfZOfKYtKQgtLfLDt5mf2QU
LbJrTNOmPeejTLz6lWemvYeBdO962y9ypwgN/FzHHBZr0vMIOS4lcs9TYhd+r2yI
pmsUEfySFnBNM3WOsYSJMTjHjXarxcAVrUDB8s2BD+ZP2Qw9zzrbjww2d3yPHtnz
LUmktTQ+hCkdieZhaaTMelFCh4fAL4tUlhc1mKU/MjirYIhYv286sEz9CJEHAsUN
eI+BtcHorQm26NKsHh+pifg4RF6q79auanbN7fVaRIO7AITD+Lj7GXLx4bgJGtzM
4yRQV8mzdL4zSyHvGy6KOvobra5NkHeIwMtvy1liIanx4FnRlV89SXvz347oMdoq
4puzB3mbyLvLlL5gGPI5y3OstXYT2xPHs+oT5BraXQK8qgChwLmm9NVyrbD7xgCk
vpO6JWwjpqNICtPGbYchyGnUaCat4lc0xd126SvAa3H6ullNDzt4RUEXXia07yoG
zfXQ9Ggq0wwzeP0bAmj95Fipem9ZFyY5fd16VM8EbqLwdS4EX8jZhiB5WcGMSMcz
agnvHENsrigENbo6qufQ5v8qUK/m3ndSIaGYd8HMOVmyjlvg43812Rx0TYgwv5or
Z3N5SNNia6/DsQ6pc7LBYFAqjrAM1dk697L+im79zOhxOvz7o7JZG/+INiep//Zx
MBWuMA4UtxTgvyMZvb3NjfqTkkshZ4OKvGpSVKVeW3P8U/7M/AKKsGoeyVSmqjI1
4RHqjWoGhLOytpvJ99gBGV7Ud8dFJ8GXi3C4fRImdcn6GrI4oUcDHlV0u65FTnHM
GhO5zMGfjBvmEm9pRb4HzqROdNr+iCCCDsGRb7N+GMuQiOG8D7DIuppDvAunxLA4
mP/BbqtXXaUdCdF0DE6P7nJMZ4Dkei3CP0AAi9zCNb+nFElw37VCNpM6/FF7XyFw
6e5Ce1iHMbhbBUTnINnCTxlcSlaFpFRnNmlLc/5oiukuLUB8QJRKBcn/CXxGc7tD
zo7HHqLY3e8LrKm58MzuCw4D3wpmp9JZtygQlIde+JZtKENnuhLe3zhoEwXPEDo9
LaYgk76PN60BapJtkOyLdDu3CMfK/ytgKspZ3U1v/ErBfJRa0usuSQXsUfeURZH9
8IjgiugxOYInDgiU+EnjdzVRGqc8AFG7sqj/RCY4RsMPQFqAM/lU8YXAIG/ne5Fh
ozsFpqlkYQqp8oTzJXs2xuCITKxU3tyxmk64TbUsv3Xo/MqQY7APkfE2qmpC1F8q
ZyjpB1u8X0QGZVi9O4MzprUYxWOjMS8Vrg7ILseR+/x4eefEPRr1q09OXHlrRhYb
ieUikiKmsQ4X1MUizDV4kSEqAcQwdf9BeDnCZj3bFQAAGq79b+sDn4RWXyxe+MfW
lWTbVz247T7s27rfEFVs/fVbp1cVTrTyMCZr2B+onRP7D2bCCE2zh12/eQJdAo6Y
fY6pfyMcu3fdvyE6cXYmqg9foF0LL7+K56U9WdblL6/3P5wiaPnx8GIdwZlbw4MA
ejqmhGHKxehjZziJ2rwW9prPMC0HvizkNz/8ROiXtEcfIy4sgJkVJtoDRL1HD1eM
W5NKTOpRg9hc0EY0JDSyQar+16x1kvbKJfQIoa+OyUJkfPzEVQSWioJxCNaLD5n9
CTSetoMTBxo7VKS8sRdIR4xvwNJ6aA7PZ9WYdF4H09azSnhxXAFR7+yt28yoVbuA
yZsFfJj9NrPvEti97ucWg5aDCYGCwb935AqbMswYaJqmDCz8aQwtfJ0+6nmuXq9P
2MNWNm0z+A1xA0YsJPEuvn0nrSKMukOJzdQYpq+eDZP+IG4ONsrhwieBD/dA4+Tv
2JFJRwXU3oo2JQLuNPTHMKqFZYO4EMGldIpnFuhqDJ+mR4pH6XskasNGbiiirTVa
ZsDHKASOwCXXDt712V8Hm8ojWZNTuJLlAMLtOpmNJKH7xK+5k27Ljt9D5Dl9RaMN
gZuDOf+vqc9ee4IcMfNPgNo90gTQCTq8t5d69Nb7AZ3H+SPEUlH8/9yQd0cIwPuc
7D3eEL5f9c9McjCX60LN+93Vsl8fOofAWP4iWQTJie2a17SQNlw37m2Xk2JTpWjU
kyPLcFoGHJCPooE/3fWxLz5U3jgZd68I5dvBI4YCo69A9d3AnU1T0nnL5HMfBPDe
mj0xVoCSmOL3gidZMT6TVDe4XS8Y7M2KnVmsdFAvhHB+bzvQJFaMOpllMNZH1mOK
bEgrIhLVwBQzUIBdijaNTVx7DORF/PEo0yb5NOQwmiQFMFhS9To9feiqqo0z7gO+
zDVpDBGWAVxsBn13G/h/Y8BjlEsskMAJM+JjiOK5PRhTanq+TkaFXS4YmyTQIU7n
I/eDYJ3F3fGn8BUMz+a11765KRsCKbLo4vTxC+wvV63viI9povA4YhFRKD4c2av8
L6AFbI8E2clbbEuKTga4NN3XB3QslEG2uRLISewvtuq+HzedGLhMuIjBo2qdEQf/
bEho2utlXPnXrl780NsjU0nUwSXckE2m+0uUvpNNUwo8GL3nEDqUQAwBKgYRlJjV
wcStcmKl5eFGblESvdcQMlUoxsfYqBz9ht75w/HeDPB6gZxamzIUpDH0VfDUlNcG
/k25PwIBMC8cpzLTwP8Zd6OIvusb8bI9XSVWxfNatBs3LQ5hUn30Jg5rXcjb20Ja
vlQt0oQe1qRPiCHlvMeKNtdBQvO45FVviEWvbqtTqEenXpLZe46zragHHpAhbimf
LGtz2d4ZNTsqPeHve27adUNtf10EgDATm0ZKY7Ps6SB124/Qcp9/EJGFlVmCxH6F
6fhJijEIIehHtebzSLB97t9OfedWtuzDndzOiRF4RFgLUYcwLvQY1GNXQA4tsQtd
HOHinom2Oy1rdnanxVeB1ColSDof/OhtGEwu79gIi0Ufqv5df2+jLsZ9RBKNJZp0
1fVn4aLzdCS3U8RFmL9VH09aQXMTrW7SviBe8+etn6AB6IV4x0jkD5OrLL9Y8fIZ
mzE6fwHcA8vqenv7ewRbb+AZVckFCTra2IZ2sVvBQe1JON/zDru2hKEHNwECbYoV
4X5sy+zcp1j8otiHEt9bpAR/OBr7FGM1T26k3TFtLrVvwbWf11ZL9k7CNPDbOlZq
mIjPEfSmfTYqYOb29GOPSGmeNtxqbpZ7GZ+TldsKJ3oG41zPWhaG7AsUVo36sxxV
iiJMnf+DbiZnG8+8VqdvrVE90uMuOnAPO+cRShthiMLLhHeTa0dPx7dOhtmIdDf2
xydfk/z4xftE0iJnIZdwf1Gu17SOWZGO9OfEyw30hJ94ysfIGcqtSNSZ/JOftvb6
DPLuANuo0yy67ph5pdLpCZA0RTm8VKpBYHdbjdqt5S/aIM7Pg6S2lM+0/W0GuFON
P4k6ELEiS3M9ZWKar3Is2TSRa2xNBVlnABZSq/mGsR1STu8p4b8f6VoqaP3KdP0Z
TnDK2TMqC+0Hawg2nHMcjVgrIjcycYrCDxWl+nO0xq32+/hwiNrWp6Tv1REOogm8
BHsJfvuOA2uHcfK6NI38yvCrtsMGldjZ42TJ/GU6Dr21IlEaAgzQkXbI5cblR4WF
1Qp5EFxrheYJkF/ljLsX8HnW1R88nOCl1+fBFLIFxGZML5KGHdbI7IKr8vk/UGCW
QGliRn/kuZA7pMAJrE0mfHc1iMQt4zozmfBaNljiYfqTksGhsJ2xkc9Pu3MNbPYl
K74eNxOQYPVu8g9zxClErNo1nul9nVl52YbJQAoMucA3E2UsHllPFF5Fm/f/Afe0
PMFyKf2V2xTbSeOVjO/RmmAwd/nRntUVwCKtUVszuDROZkrqT6HI38tINvUNKcBl
E81CJXoBHpVY1CmM2K8yGRWnCOvrqzKdULIO2tXSYK7mc5UiVJ+i3j9dhC4B4XtF
hdsXBFKLiGZsOplu2a2+K3GMwmKXbmRDbU+2YaZqJHpjMYPHpG4Yz7zvCUMIyE/o
+O+bLWeBngwUumMOYgikE70xl7wC3a8+uLjp/wJ4O1PSL9D2PkenJ2+/gmSJfm3i
Qzi+6paLRzoqaWk/BQDoNPDWLgjWwTFmd6dLwRZjzy8BC53aaRYa2bmlS+Kvv8xP
vIB0HKPAQnQrB7k1vOgyMBWHp7DxYJQ81R3y6Awsgh9jo4ajYrHBc2BmWhx1FId5
CkIXdlQfXDlCI+z8zTxVBiFRpIPaLkL1VOznnf0kuduUQRi/CIMibpfeBTzUe4Vr
eLXcRdISp76C8uKsXuuBCZcBqQCbVoUKPVnUlFz2iNEM8YeK3trsXR8dlAtuvbDT
EgZaH/z/5XooLTjar0VYwixlgCuVsbrb3+8S5jm28EEbGOkbBRedOyR68h2mNFfI
hXu+ooJw/UkMyUcchsuutkyg5dof41nS17kgIilcqV/JWUwSkKKWBR+dwTB7jZ9S
jtk2/DRgfcbf6On5dURTlbS6Brcyj2hSaSyG3I//fEBUNQAATZlTOL0hWWhHVZRX
2oPZ7/IfuW0kGTNHGHvcw5ao2xnCEJH+4YW+lxKnHvux0k+NwJnuhS6LWA56g0p1
B69JbLS3AsQmQ3HYY7t0ZD2XidG62GcMbH8bsayBuNffYivydhnohe/LuOE3yJt3
ZuguxLWery7Y2haQpgqFpkNxZzU9VAbyJiXi4uP2qCuEauhs48lGHIXoyB3Eg6mo
N/V7lEnraXgWJ3H9Pjbohm/lzPcbTBkCeDJJoMleYAmAAuVokgdI+A7u7DgmMeDN
cJJ0QBXnh39IsykgpYrSWJ9XMQt9/kkKll7jiwt2dqu7JVmJyASL5oAqnc0xxNsS
VxOErOBosMAO79r8pVBoTmIYQObTDXq7gnIn+KWs8ITcMEmUJd5bvLTEg3CsU2Kj
CtTuVhJA/DNwsiH+qjokGI+yjbabOxFfzBmQoXbbNMjAytYR0A+vNiXBviDJr8MG
rH7bj+rEsLOhcqeS6NzzRlvjkeHNITF3IGohmYG1QjOuj2ydTIz2X/8o+nzwJ4Cb
G9ReECd7+MBjZPBKH/WXwTkFo89JAzQ/dINFC5gs+0f0jVz7fBgfcSO/0LY3N2tO
NS8KmAGzenCMCfnoH+5d218irzwZcaHLtjh0ard43yX5Jxrlg6Q5nllgz9r5YZ7k
EaLko2Zga4mbwMg7rEcCGRj+Th2aqPB1LIFiDVHKLBDN6uUTAOsW9hmRkqlyFHoD
aWNKLh3XFj1PaHs5nbiOvuWG/gu5rVICECbdgszbqM3QbSNNckCD9nhxzidGrkUn
YP/HIe2OADanI0hgURMR3out+ZmgVGlCbkonMX4YwNNih75yXy8Me71zVsAlh9lw
Gq+7Wr5u+fKnYYiKnlz7Vq0PnYaVZLrTVHK/jCtjzZ8+WZhauqc35yX4Y8pXxczd
iTZbxhtykOfgQFVjG/FVtOHGqP5Mc4ysJwfkzp3nhOx8fNfbmX1BzRT6PfNYm95d
rUCaxNTltQJY1lWG3rffyalpPuOz/j4sD51G9R0qVLEGjRWnw1SW+zYqSXFyPTUW
PvQGax568oPaNAXacQLsMrRqu6gcaiFH/I45ZTuCLzVfMphuNXPiteU0fBetZbqi
8SvFRk0Pl8gpsYfq5rg0dmo2sa8p4Uu9DHgV7CSGdVndC2kq76mUXmyVfGHEnAIG
NZ9r7BlwgVhWGz0S12BaCpN3BDfXqgZvzgyugIhqgbd3DrFfFybDSLsGEthflK8j
bX5ZjD7xQbLkadoTBqDALITmw9zzcimATrItdLQIgygRSAIO/v8k36bfBwpppJqt
2MNJ8q9QVywcUf0kA/khlGLnHe0fNSpJ8ezNEXDEEt3O0a+4e+h38T4x34dzJS7B
r1oJ7CuVAMzAql3gBqqfLgtO6fxr4TM84TOdohp1L3YDMqOzcV88wzBm/yDDTuUk
7WmShpljvx+KaCZlYQpE+dbdfJxGyfBF3EYuZZM3uZr505QC7i0NAEvbqsM0NVUj
RqE/JgkgzzWtVu2TSRQCl2rdMcWzcgR/DpijDRXzF1KQBS9E5qfqH/ghByXnb69y
SnRL0zRb3XwnDXF9zzq0CaeYOf4A8u6Rrm9va6MRb9kyj4IH3RQlJo6zMZVzIlFE
/HEvYlKf1+0L9mByuSOOD28A07+LU1BW6imssau6gFi5u16r6qQiOFG0ivuSFCyq
CkNCwi8yxztUOIfTAsQIm+7AzQSw3MpafhfwzNbpyEfE5wYQPbtcNv/tVHZeIsOT
wZG9GznFN4ZUhrn6ls7rp9mU9kY9fS/l9QWCcgFTiIkicAqvhC8++JtPaiYpZcRV
wslIkV60M6dpHc6eWGc5vrefsibBXaONo9zqhyo1HQSDuVB0ILzOelXxRrXOjQCj
m7OKJzbvZd8DW7pSQpTjlhuZlaG3sZYMAwgynTy75/F6meidFVLYq17cmdmR6YEA
9gUK2AB/Oa4WGlavYNauREGJL7ZIDkTjTK5dRbngj/Y9GyK8MDYhpXiD8kSaUxKf
Nq0ggCeMD+8Ijj2ceyRwyIAgctUPKabo2NiZmfq/yOVDrNcMr8kWhudPglQ1s47j
ZmVUEd8369VFBmV0gnXuWUu2SHCXtx05G8ppa1gf97xlVqXddtpKbT0c9r6MB0F/
T8kqOs+OJMcwaxgqqPNj0BonnryGByDKWe75fzUDCRBw4PlB4NAuHKGs5iNI7k9q
3AseMezhPdTexjgM7QLhZkW21CSQWCMoJF7wNx+t/np0icFae/jLVctMd3/UlIPu
nGwpL55IJlmIroiEXZVNVIablkF6km/E4L8I28FpCO8ilQuOvqaQ5PoZG6jxuaJv
DmThakBucRRxHyTLL9T/+R81KdicNmDB3YVfK1/BF6UmBuaWyr3YtsxEHwFAfCxD
h64mab7YOUP5aMXCTz4qwyqEkCpRn9h3Pl0yL/pvFjFK4CK6lgdxidFqbxC/kt4F
eY4fXzfeXmtxO8ydcBzgU+PGpJSBgwpuGqSJnYIO7xj6mV3b9sWoYM4YJJrkDjyH
aa8zXHLMwB8oGsCPtb9DP8BXTP1HtjW5Rm+mi8DwRbAjla5qLnPUlnz+aREf5tqw
3qoLSgc4tJhQ6opOQlA2hdxLnyCmcV3rwYZHCBx5Xh6OdHtGRJqbdxpWBcYU2P3Z
hU5gkePFf7ArlzYB2hua3ZjSjcvXSgOj2MixzgWHH8TqDem3RoHK5ie/1JZc4t5Y
WEX+W3T4DuJ+UcRtU9qPlwT6ndjb5XBf44D/qODrl2S7GrMZkzn1TOB1+bo7yYTl
bZ9Jrp1AHOgsjZH7SdwPGVXO5gnkkub28wv/txZs6HeJIYFt5CHmwBpvq402T7pr
gDq7LWNA0OpSpQgGCC2/GLcR1w/TfQw6i5w4XeoYPJtImAYLFhI/3ZCEa3JTBumN
+2V2EUlVOE5DZfCzYyTi283OlkbgCxZ2HrXevWl/urW9Em17Xb5VMHAN0TPq/FI8
KwryGDnUsqlvYkzF3oHksT6hxIQO4xhOSgQpWVohGOCfAiGrSYuZp9ulyQNwI+rf
zE2Nhrr0BkHDaVRFXldFYF8tF4/19MxmMGreZuoDt2JSk0dhGe4eNcsAq0r8UJSh
5aaEkhA6IVekBzKW+V/ol36V5pt+1UAq5AnEpTl04PA8jpEe/t2otu8X5K+ziZAC
2+DJ6L6cNMjuLZ8qepeFeyuU9X1HWHL3LTxtkiAcyQA5DKRRuWn3sepVkKjbeFsX
fAZwR2OnGcIwux7q3PenTAg5/TI+Lsi45HxURthKOcGjy27FfQ3WCCmZfdhKjrzb
jNLWcdsKvJxva6Qe4C2O0Eyfw35i/zNmt96DJjg5jPDOCnIpZCVqnfIEFzcObO/W
gSareUESsso+bJvlJHfAglPgbymQzFv628s/QQNT2ewqNAHdHdQMAV3lNfdR1qd2
SMo+MFsxOc8Ylj7IhJpJPae/ZDbSt1TMR9mPSxlDeTRnTPpOwfy3nXLrFnKgN6Ly
+bemT6w96TYjZShWR1UmpwxN6YyVHSjtDWxIi5xqgvyJjxGqeE/FdnhnbfN0oSR1
bCaZdaPZ3S2tZEgILxjzv8a6l0DncojJlbttURtKh3mQSB1jQIKkTk1LeZApoRgF
unghLkvy/oW8CuNfo7WJN25PtSd0VSkWdPWLVdwjiVPiP0F10ULNC9ZNIa8d+9AA
+zR4/0XGX8FMQxPWj/wkIhRYMbVRbGVO5q+HONVQoDk69PtVJsFZpKS2yvXaEt7n
rL2yVNvBtYioyewv99E2d8kTUgnw04t6WwAHlHuy8CbML6hbS29FIZlvQ05vTdrR
j8c/eVTUcxRGXElhVC2jB1eTGwjiuCA0B+yjercn6mX4ClsGgvYknpoWX14majeW
Tv/zMhJavvGsri6rqylEGSUeKMCXMeLTilXIdYwW5TF3jgZf1A/NhBS/kEgX1EWr
gQi9e3pEiihALZXCuC2TQK9mZyU8zb84a5iysgPWrPPPDMw2PR009IR54LPU0hSS
rVKw2ppsCERDwIq6fQed2v+P8gzB5Fo4hTc2Im7aTMoZTGsw6nUCHbsWq+AC8bbU
E83H+DPr7xKi2dEWZ4av54sCIntaEbnpo63idygxLcZeRmoEqJMg3FqdJPs5Mzeo
rgZCJ4MFlk3cP7H1HnPWaaDiIllx+3tFzjGso4T6fBgRoHFsr4bzMuFFeGOCZWhI
lxXIpCtymlrlWvCZFgwRfSdgI790Jhhej7P6/voYuEFkzNJf3FlPwswQfgcvzwPe
js8cb5sL0L1q6Wwt+hRO9l02Agnwjpo9kpqLH7q26yPg/tZkEEE1tsKE0IqshTOY
zOfwiGvLobuMCNK2a5Xw3sfKbzXbE+f5WG4KpPv2e6NlwBmK5hn3FHp76TI/0GaT
/NxtOd5Liit+O7t/dv+vF0z4dAN3u+mw5SeoYljLWPThE+Vjo1VwEHM8gxB1WSTy
OV145SNYECTbR3PVtBFzNS7VjuC3tmf57vX8zm9VGpFo6svJeq0Om5SWDK8MfDJN
daZ3GPXKFyz/5sEcW/JUSU3aqP2Jrd/RHlj5NSMolJN6g0PJYoC+VjjJtkG5pYHG
QF+wN/ONs998cyBnCfnukHYaWcl9+dz/GB3kJtlZpxDn/G8HHIU7YGaifFK1RR7L
Ektuo2iTCeJ7WtlmyoRTTLJfTUAXadlTa/RNOc2tomUzjKN9X4lE053JiM0MUhFl
ucAJDlAaxg/MFBbnBBgZ5tpeUxWf1DxfXurIhUeCU03V27Lr0d6fzx1oyG2bqo95
uGmF+Ol0Uho5mZCPyeaF8W4W2ccBw9OMALVjG1S6R2MPgN4QkyIpUp7IQ7p6FHgT
vwRYpP/H7j7pEHvpSJnFsLDSm4OMXnZSGColH+Mr3AvmtTC4efHc5UPSTQRVaDQf
2zazdDHLcy6cgALuetDYn/c4w0T4A0Jr7tOCv0p+pAE4C+7IDDuYe27fSFHS6c/E
IHJRYIGW/LeWJ++QnrCPW4+9QFq/lKjtdkPfJ1kwKIXTVpexkbuAV0W50hvpZj9m
BdtzX/ehmIDE7upLq1Mw2QAG4OVZ2df2MSH7LmJXkiNNEEdczFG94LT2MIvDiddZ
+Fyb1D7AswidslxUO0feASl8gkFMsqrrXOltwaYhTXjFRD4q2wpyC71VmfZRxLdU
tUqn6hEaDWAdF9UujUhr1x/E+b1ByB4wOpq6vqf6be0aQ3pHuF36iPBHy3b0kC3k
nZDtYxq3Nhy4/u+NPIpcvDYaJDqNqkTGM1Mskzz7m1S6T5Cnerg1jw/I5rctEs7L
Df/1ThPTya2YvhHh9Zj2XVBU3CXiNW247DrRRdwp9AElQR4jsGzvpWOhw1WCGuOU
iLtVbwwqoKop/T7vrgNL2SBC4HJpZeDfELm2G54kfoJeMrVpuidx2KN4TwrdEXBZ
WZwdRPLbWfj7C6qu/L9y+aG/m7WZRvmLm1HRdHVLmAZqBNH35tlghgyyHzylDmek
ZAO2QZav53aBhmPiSFolXG8B23p63jUfIrGCNBY1XyC3Uo4IBWQ7pbO31NFnrUit
Yi+6r8NomTS8YbFmHI/HYOrD/VvaaObRtkeWPka/PSHqoaHw9dTNelL1lJqYj1SY
aw5fEUgSf2yb0hwCHJ45GmBFiupwVccKR8mLNx61E4A3DNXPvESKhJqDcoQF1Mb+
XlmgEp+zVK/2w9he6zgxx0Dfrk8ecTy0MIhtt2L3nTyhLC5ScL+rI4Bge+CYMo4l
kP6I0JPTLJy2/2ZKy313JkDY9Tzk8yZfT53Rsq3bPOlQH77BCgDA+1AlJx+Xj7N5
kDwyn2kA2PCZOYAgavkikZzwtXYIb+Vt+6q0pPP9B5ZqjoFzDsCMBEgvBYyZmKQ+
hO6SvDLnVqU/VE1KOTbxIpwPdYMifpR7RNUhBKU/ffesGuykaIF1XqeKAnz/oeW0
Hm5Pb3IZISVAUeI82bvz6FI2FJyTEGvj8BGd7ARmy/SbqJKOrMpKsyXNz6xqjWBN
D0bmVQQsU7HDkWHRFl/iBIRJbEXj5RMjWrZ8+C5EVILb3Uyz04pA3+bK+IWERU8O
sXgaRHrPeAlQ0dEY55mbiY+LxN91hnB6Q3qZo7c7Mj34WMnYkcZTInoMYUOrOK3A
WJG6AnWaVDSL3N6yFBZxg9SXzu170GZ7fb5Likk3v/SqgyiX75j3R5YBr2qetN5G
rNscfGq9qcq5CyDyzEOYvpIm+zZh2tucWAk57pa204y6I5Adst6aXqnAb1rn6TT1
fI5CvnyCupnQ6xUcBtJwRFHrvmXQi+xXTzoaxOS4Uh7A2MlVoASYa12T7FpZpp/U
Oj16bJ03v+ohvWCsZqewHGfx628OSARuptdD3ZnOQwQZPu4n2IlywtjLdhOSp1+k
onGkmYC9Z/94QCE8d9XujhcH+kac9f1vCrzVBV35XRYNlT3ijTSj6jrksr3E9a7o
WfFPB0iP50QzUcIqQGAhOtkPDdXicnwtYBR+mWhSwfqWqHDkfu86A8XqLerCBPgT
Tpw8Etb9Q4qWFI0DzDd1CL8IYbtJCxLqodrbzvPxeUm9wQ2f1rpuwecr3HbuWiGu
JfzWWhhnWx7kUu5Uhn0hYFkVxoQo0tk5TPEKPB0X2Kcxy1pSn7daNiBqsJKjDPqB
0YqBEK+OjCjFo9rjMyHCbhozuo9QwtUgA4CEz3r0ZAEqfXfu77pxyyNhorMNMEln
6Uz9acoBKngbFaxEjLBpMiFuzbDNtwxVZnYd7y3IJsVS8253xPuKfMmFi2JVUL72
3VGMmqeWaTWqjZK2nFzTew1HA6JSWBVWLi0Iwgh8i2Sf2dx9lljkxRcNtZBXEHNZ
iCvgxApT07YXEHH974IivdmTlJbELFnjlsWs8YgRAZVCiAKJMCIRmEQBoEr/SQKy
ymSyc7E8R6QA7kL31uvedQ/ip+VHq3FrvcgaY+vq+qS+cWQOSYZb20E0a1W0MeIw
y4meT1eVaJYtio7bL/9o3bdQi8pQN7aY28gyFAFWb+BL6jfS8WQBaG+tu4IR/LAE
grMcO4l5Q4GOAv1VhBkQdhk7GEQOEW83bkka+TE1q1u7jAmRJw890PdxB6RWntt1
CHKJ7Mq3y7tkmMWRaHqgg/vVdb01DJshOtJav+Qb/S57gQsSRPWZvnGMaYHBa8xs
w14/bB3tAQPY7Oy5KRznVzjezKTUtsbF8OMhUiqaZVKZdD4KDVBKsM2Kr0ZRP3EW
HFJoO7wfMzwMGMjlgkr/kxy4vlGZr55/S3J4EBUmqDdO5GU4ubD5d6UuyRCqoK8V
yJcwLK01jSChak/FxvWyH0KnOSq9kwPXO9D9CI7HFErtjEzME9YqZIymLhpGtJQp
zQJimSaKaFBJzRd59yceyc2qYqiz3KbN3PDVFy04EVHSW6VRaDETEKahB/A+fu2w
QuslQjmTt7crgsljaFor6KvStiGkSdTF0w9t8zU9EV2qLkc0G1/+e3MenXgry8mZ
1p732BsQqlIcbvZoY4InXT5mjLC4nqd+eLd8NG9d/Z4JCxLUQMWsC9R+orPZbhCD
lJOIPPDLD6ssH8qi+Z5YTCphg/jtqi4UX8MsvdGVzgNCfmT+vYHbTKkv8aD9SrJv
9ZRAXt9fC6YEog4tkgm6POnpYGCzIeDMge4RnMJJ3pWNxLxKCvMIP2OITu88vSrG
caDmj7ww7XzQst7bqsEz9HU8DiYdUp9EmhrshmCOTQS51tRpXdmSqeWMAM3Q1+42
XY37SwfpIW5Nc64RQAqvrFbcZsi9RG1vZnUA1x5ZPujTMoHVIbgP3/MomhZB0JM5
2CCARdd0UeOAMfg0S0C30I58xHZgt2m9f1B+wn7Uqv+LuZ5D76OtvshzWlfNFm6c
t4L953xPYfO095GnSpH7xXFIgB6UBpL5FQLHts/Zen0xEnrW0bJjCFOGDhjuc0wd
6baQJG1+h0xYoZlKNA3BsczOrtMKdXtVubX/lA6DUnhSuZoeambfUYDiorzIIpcO
fknj/99tFv2jX0ID1RDlPBostx0+uQwCnuoAenKJR/DiR3ND+6JpclFQ9sqPpG4N
lq3CHETp90VgVt7kqxRWhdCmwhaARnonkJqrLgodKbtSzvbxza5opOz+rrWxpQm6
o4l/7/xqA3LXDJuOMY4UNlLvUY2GVXwaw2v27VzNyOEW/VAwL8tjrg9WTire67oB
rWi/Qd2L0AwTAz7LNf08efS/cDcuD/cjF/mJ51u0V8TREhCQvTHBUGG7jNKbACHm
AXDPo/VSvHH4fb4QgU9CE0A3CrHcx9bF7qc+bMPM1LhfEQTRYNWyTwPn6kk4sCVi
5GeLo3EWCfyMOc1mRM3oINyljxl9YyRdnxVTtuetsqffg2Z8atdKBl2V3cTmmhRC
yaZU+Q63/lP+H7tdAx4kYbV06iiNiH4wcTCoV/VsuSGVcHMZ7blippVJ/CI58xjP
NxdcfjaDUr9S81hl84WB4z8+5bHnV90Kror2fCIgDAZeFh1cFm+kziqHRZP3q7cw
sTzxStMmRaliEdOEUHhDPR3schJsif/aSy0p0acNVkknnQox7ne1DOsCK0JHE/Ra
uYka+3AtobEShjN9W++Zd1YUV5y/+dJJUll8Gsv0gEzOn6JpKuHGc0RR0p3aEbdV
WpwN+AFQyvw5kfkKrGMELYHQYsx9Z1U+0WKtyAtRzI6oCPuuFpoVfBa8fTEjrumb
hPIRcnHwuZMZEOAh/m256GdRFru3Ktgc9EaEgUKdvsrLNtTQpKsZs0NFeYaeU70f
2+1SmGOCDwj/NOqGnH4Sin0d6n/VexZtV+CKmQYQP0Qss+lNwigB+oZYPMTof9GB
NOYH2T9bvZ0nATA0a9Gk6AWJFtlOGt4UlNBbOYKobwsP57+yKCVBpulDDv/01dLF
Fhw5bFqdbPQKIdQVH2ACRDQ9YyR9fhUPLi9Bh3RTAKIXh5qmeWs1Lrt/pCrjrBL/
gFJYtmxoZy8phQpKYrMnfkhq4pojbg8+7IuzFoaRJ6Rq6kHxNKn5JA6VkNnaLphy
Y60PB3qilSHqIlnceaP4AtchF4CJwQiOUmc2faGo3nzB/VxO2oejRJwmPes3BOWu
mFwMD3ermPsE1QkttTYPygAutYQD72+78fkQRKEmGdUN8ZIUkJImyQHmRojhXB14
640IFzbVsx9bCyIUAOuxv9jhVExKhzVJ9y763Hiw9MD5fh6oOhOCPn2ij+/ntanS
xXaaA9hTyy8Tua7H7tKzNy1JSfBzTxo4acKZlS6l4yI0dmQ52PQgNLwU96g+70e0
LSA54JxQe6ubA0hn1Aygb+/ZX7kEIqKHrDVf9uU55VH5G18htZvZIOkb0J/rNNVV
QNcdHVPi8IIDOvY6H3CwaQRaHv4FajKTYTRFQBXaBz7Jm8afqSoewPHCtPny5MjQ
ZIEu84CeuFum/XFKECjx9uUD1JdiaHBl5n8KqzyW/qmUZ/p1eCaOJJHy+CkDfC+K
mkhykx5jDq7imA3+GNNzzQI/pcdNpPuklvpYsvzpHXq1xb2VtkLFr71ivsnmScFf
RkSD5E2+yTgpB0XHUqlypjHKH6mdQXYx5jLgPiYYMeLYyavQxmtdsX/W92gHKHfI
7m8hpL5n72c1GggU4GIKn+BINY8ORVxN6qEDEUg7wY1vdl0adK2tJ+s1IyIswO9P
/tRNYbnKfH7Vkze0DxMIGqnCIpO57WjB7VwXbvxsUGNI079fg4qjad806cvy5H6G
EThOcwBV9YFpeQ1RjPnX7EcQCeCLWSndEP0qfXim2iQx/7R2V+8rVBU31aeBoq+f
ZfNm+HtAY2thi8Od6PcL4Nc5JEegBmBg6yWxK0cYQD2id2UVKOZATS/dp63K+e6a
hc9hiX49URjfAzDAWoGml0Go7AviMC44m6RNeYKd301vEjH1XmR0J6o8S2vzZsh3
UdLBdNayFwTs72tUctg/7dE1BIBRbv3QOXWCm4BOj49YTklbYJQc55aIHwUco0kx
aDi7zczUvDZcMqDZXCM2S96h6YGJo8uBh/KuI9J758/Bad99s+QSf5rJgbW5hLcZ
yZqLZE1w4vi062uYRmBp1s6GIKo4ZNsClRfJpD7CYimhY3/GyNTBu2Hr4KcsIjNk
d4bcI4VC9ln6Ksu9uJv06oqe39RlBI19AHm2SFjOL3Jvz6unAN8w2e0VM6y9k/vJ
b+M6PjFaIbj/7jpxOldxXetYOW3nKFClGUKN2mqKxv6+bLg6JyX6YNpQkzhZd0zA
4LqFrAwTuzGGE8psEh5reBqbk1UB0j2zFketw8tvKmMQYf79+YfPJuArVE1k9dbo
U4AKgzQ3t9epfIF8iqA8XOyYo5jtYQNE/VZ7wRNgCEAoEADeifpFJg19SFDTxZqy
Mx4I9IBzvjrDegjDGTBAKBnzncvHHCC478ehDWWtzB8lkg3dnpLUjL5Y6QSatUTH
bcDueWOTwEFC2/HEXEinAIpd1DNk0K1ex7sY0mM5JHube9D1g7GGkdRJF+MskIOs
BZh5uvDvdgTys/+N7BsPTVK8G8oWSdC8rKAeTN2XOpI0WsIcIywjMcLHGebvTYf6
Zx7ErvoZ5QIxNo20lQx01U9rStkVwHKXYImmzdKHLzJe6By8FJ0FMwH72npXdBAX
OaeV8pPBW/oEsCvmdNqlJCF2wmQrlrJLhvYodjSb4k3883qDRS/s70MwYDqa/UHr
0MgqDwE2ODHx0PkD/KH0bdxzmkxC9mmWAcNApDdJB7szfEAz66S2lSM3R7Ws01T3
Ea1p8rSiVYayiKiydNY60VVS7UdxG8u2/ZZrA6lYk/ycqfcFyidLiAoTC2hbp6da
3iSUE5G4ECnCxMuF0AmKCewqLEHj7q+nOHPMlAmXeSvonoYLqc5Fyz8xgXysZfVK
Ze5a40X1zWYLN/Yx6Bn0ZgvklWJU6s+GwokHIdlFpDEUB8YhPICLLbyKybNt5rED
SwIijaHvdJL/gIMymMBfL1GP3KSPNB1e/STJSlVG7XV4sLilSB1z3jQrrS0dURPF
JLb3WvP7u1K9wE1KlD5AG7v6Y7VRHl9SRj9QJ8NM06yCLeTLhOMtZUHLFaEDlPop
+H4stLn90LMA1X1eGN4niCfXIycW+8h3zRFAmLHot4YC6skzseDWsD+avWXh1gjp
0T8uYsOtCrkHwLkRVs2nY3sNVzdGpI+nCQtb3GH4bXL+VZucPmKwLH/LJrVlbR/z
YmdycSFJNtFwfO/7ZJPE3h7raZv8sQnGjrazMSYpqN3hjTMncM/jghCpwdlO0weW
Ns6t64LbYgcMJ0Wjiskle67gjvjdqgztooO2hCGy9NnMbqsgAC2KVNogrY9mtCbj
bWkGMcQ9s1Mi/qZQklO/DsdCznYDoyK8X8GepBMfRjvYuis8VBoJL6SmQM1bLeZH
ax37nY+Fa4kPtQ14M12D8IPOwRCDaDnkiPjEn2TH6gzwBoyJ04bwqDbseMsu17og
/HopA3Jk42PFTtlDKVXbITgF1b3Ty4l+zT3ZWi4ji9satY62QLAo08766fA8XyRu
v7Th6bhKTjNRkfaPaJoXE7Me+NfTWTAVeUKUQ1N1iW8bXF3Aj5Gq1hAs2BnRaqiu
XdUBYVpi5zkW3E6dbmJuIpY/DAGYDwLNYqcdW7mmN65FR4vSbafifZkH68OVzjWG
wTTwBBifjgajKr/mNvpYT4IlatHsaG5Jvl3XD/+ZCvxHfMIDJisgls8RzANxNMek
0LN3f+meS/g4IO3X4K8966sbu/TpFRPIF41mqbwKbqZZiubMkMnJqSQBW2HZ9C2f
Rgl7NaLYY5r7ds+LOgTIW0ncJWOxPc3oY8oGOoQMmb0Vq9Hae5Epox6eh+7BB995
xlk8HRlbAbFgQvVBIm+N2TZVnjcy6F/YvlkzFBu2jmNBKTr6TZsmbn0V+OyX+3Ah
0WZW0QYPkAeu74aA6IiAfnXk8BNzaYS4OiU83o03Bihv2Jz+FB+yC5+8wYGpg3NI
QJbbbte1KzBDMvUsreGVzy7Th197P2oNQdWzXsRHTKkVIh+aWVN6zheflAcY85nH
ycKVzvJ9zqhoCtf5e5TWD5xB7H5k9yOsJlcJ6FIONucJbho2qgJx9CtEDdYx2cpr
+l6LSU330ZSXMMsoqg2w/HUyrk2n8khoWAQDON6ZQigzo+/K5kYgIM7gF77F2+9w
VxTELHKxERpfly63Jyks0xYpJfDinoPF14/Hy1rxdKidZ+4YM2Ht3XqQIosooCdD
EGHcxKEu/nAW1fDdc7DP3dZHDsUVhkSkH7b7Jh3p5v1EkjC/MbsnA4UXLqYtZ1zu
ExouSvCoL8B9R0Yd/Zsp+/iF9FTbbQchJJ5ZHXE0pmgQkrlnFStbBfzfs6OCvnyo
ytX5uXr4VIf1ZKfgsiNI4EDOQ/Ipe2RfB2nmmzyMum4495P5ZM2DPP0EQ/NPbVnx
bkAnjKtM59WdEm9BC4+sk26PrhuPvcvMcZF+8ZxhlS6b181ZIarcW1SHQIgkg7hr
Ff4i8lhRZHTyAnYB2ItliR0tQ7Sd2MHrXO3AEqlEOWZNZNdLOnvvOANOC9DRaHy1
dHPub1JGh9BVdWAkU01qAb2CmyrU/MRRPXu5yz+CwqcBv6s7zHs9EfCmR3r9fgKv
zGvj+vOup+o+aeAmD2RgsAKuWK3k/2bFosQPaabvpX33B6nLX8QdYWDAXd/tTLL0
WLnkC5w8Pn7I5bqYLUzu5rexCmiEaL8wZJCNX6/XEnQhYz2ocDrdxNCidVAjjbx0
O+5C6eR+Bzc1PsCyXhDVMJpwaoQkHfeNVJ7aOWR+Cg72YUdF47ugPWBIV3mX63qR
hEXUzPP2PL69t4/5ZbdF2MQxFwSy5LQ+sUP/hsq3qmNcMObkVZH7Nc4AmyEtSoq4
ME/wol9i1J2jCwWDd+PJfwvr6eZD0ayHFXHBuTsPzD5vj+JTLkRAPFF5J8nZzjsY
r+OrMB76/q8BVnjXve7Ua1d1JVDFO7eXrnxv1gPmNqrjJSZcN76IBbfAsc32Zahw
7yMQHX6uN4zi7lc3P2I8ENdbOJglHVOIrFEMW9Kfd+JAJ3FCDKs6193rawN1f3Lq
hnndkXA0Xc0cpljw/jkxUcP4XlHGbMy1Q9f9ErHG75z2gIyGXgNldKpwCBEEVF98
+LnJR4NTe24faIQQ+5GfIEreVx7uoNAUtZTcUJRKI3zXZnPWh6pRBGEyZfXHmtbG
iyvleH4YUIi8duMh1mWuCATgua6eON/p6CIvy3M7Yrm3IRwrA1txOouXlCCng+Ke
6RKcKBdiSSsgw1AOW9caU9K1dyB+rVBg7JsQEVuJSYQ35npFx/Im9i5n0QtIPk5Z
csP/7uCPs5mMxU2zWLMXsLXae+06/ClCidldfZRC2cKJ3VOpZdNxFuc3gYVkN3o3
bqDovyCNmHSBQJrgjFnSc8Fy/R3EMTEDQ/NA8wag7xAUr8uLv7BGXx3hLgz+lKRe
Iv7vLLSXIcOOmeJa97zNFeSd9VydR+dMd20OWBT8x3JWZRRQkRk0Z3pgElmoD/Dr
6o96AXobUQftVIXiI+sOI7xfzKfRzZlC2oC20KTWgpZVWtvUspM8jIN0ljNuXHMR
HFEm000lZo6H61qYKoyYJMRxkocZw0lbq/alp5ZpvVUkbLjLIB56OY8NnSrD+uTa
lZZMI5Pk5ZaRhs/ooyBS/busDdrfSi6acDfFYtfHFgHWsg2EniDrtNgcSbV+KEHK
dZENi0AOjEZ6Mtr8UFdkiENuMeKD1buW9xMUrmnM6apcksBH9ltRBdvF3qBE8Ufr
a/4HnSYL3eo4gKsqpjcdbb3yT6btitKqVdEdZFz2qSnlg58EwvlIJPj75GUQovtg
k7qtCjiIjSzQ5TrplRHmGO55UZibdUOc6ATPR3X0ugXV6NECWpbKvZzAAZcAx0gR
+/Y1+mX/sRMd7mYPgvPs/dZFHAW+isuIVBqQ7x43D0t+39j11bQHoJosuMpNzj9u
DAeLNwjCnXTl2iE7PDf+f8jvstSbNExFkJj4KVpwnc7hEIJ/VcV9gcSkmA5K6G41
Fhy3JcU+hK/KdkzhvbJDXjH9oG+hxPHF7nijr7lhQtxx1GFPx8NY/ouST3leWki9
N+Cts4mkIsXaB/DFE5XHw/vLnP38xdmhZVm2g/rqql1XMwLEtaIxDZJebLK+BnGi
U0Wu9bg1m9uYzFukcaksxjjK6XYuEgWQRGZEJyUVdM5K5esMjHBQANNd6tw9JM0a
Idmkjco874OT+kuv+fRDD3kimXLdxUwNmw7msfzzDB1B6WqAnC2pl4o23E4lo5CD
xDYmjk68fpjq3S61tY4wmVEF8IIcefDbRiWLZbIMZpDbclw2t6z0gBKZrfjDEyNr
ew8H/C4IoPZVdrEtREn5tDEFSmoZPTxQGw82PStPgdb8UHGgxJK9gYHZtEobU0g3
3x0qCGPheUwawXrSUp8H0IvP5btGxyTDYvp5O+7xiBqJjBBmhBTiSFmZcKn4aVBx
HJRbJUWmNSl1wWXIi9a03MNU70dUAaShCbkdMuRYdOMOPGzQwBIVNUzBYjAb8uom
vKJsr4mSB8L3N8pQimm4zksbTReIYWJEKlYNYDVbh1IJ3iefwbJhcRFQ5Ygz4Z69
ppsHx7YHaZXyW0GfEvQ7C3+KEHoQWkEv8RlkH6ttpy/TJl0aEksUHsP/YQ5PxsL/
vVdjq+FqDvvTT0Lfh6Kce5kT6+EhD5f2aELE9Igq9AbwlQ7LWyLVk+JuhO2jF3aw
mPSg82P024314PGtdGiYBnWaYaF7j6U6UQMJOnYnJhecy936qNl/seIis5+7DqcG
1/TBMbbRtHRD4JvQJmWIHzFGZ96BnqOw5759ZSIBxNvPXEcUe8T5Nou5X9uc5OYc
epBaAxXzUiCSQTQqexKn2HmeVVpVH1mzUqKbw8rB4o0MzZfneWjyhYRCrGbcQ24V
wkEIis+iDT13q4sELhMO2k5AJvlQ5ldm+pKtNs6QkUT+nk+bT7YcJsArOQf6iM1d
hiBHHDUThrTHrFWDkM0M9vU1BGFO/GWBv7xSNamwbI1ZWLTYsKaBnAl+uTDM/dCV
s+JfdFGluTmzEhxDtJyq+5C6z27KJljnuhD/ujPhO9RNa6AOy1BHfGK71h+hqDY5
ZN9FvDDqEaAXnY690F9VI+GjH8yY/nMLo4OVbK1zBI8OzrmDqdwImsqJ8Tv716tj
IZnz3a/iqHuBUcBj0H69s22WHncn7CF6uENDNFsmg9U3KFlzUibx7sYSzD3f3LSk
YQtAh+t3yY5v8nS7zz7nxlf86vjzm7MHWK5BwOHL2jbLNZxUFIK4pXRu2fkmMGXh
9S89yyGNB6xBrkkeP3y05h4kMtPTr3PvM0qjTl8twQccnd769xwpnF6rxCMyuwFi
UffSIsYdhHHvAZ/XSHgv07FcM6rlpPNo0DocxeHDcZ5EPGU4az4aVaktsxd9GZS2
TVgg/z+TinB0JjepLNumqhRYR7CWWVlx/kwjH1JWI1B9dbD1DfjaMaLlqJo72XK/
IJO5PrdawAWH13rR6tlfalNhGm+j3NBhWPCSM+9q5Dr5DPFk0j/93e6OUgos6xiM
baifMX6neqRJoXy73m9FRMNfwGrnNe8yat02RfmPoy9L4r+et02gpAKFXqwSZ4sl
ylb1WmC8txOy4SzqoqmK7WiWp+7kZIVh0pWEXB+BxAH/Ah6PAXr9rPsFA7ewC89P
jko9tzi60lYDBT1u3kqIdNZb183lN7Vj4+gkL2XdwD3TxWPdPibKrZRAabmf3MUa
TN+KymvgcNSKtFcsQvR1yKhen5trXdq+26vQWgLuUHAOcsRqaGC5AeswxipIT4iD
955wqjakKbZOJDtrb//NVT7CgZxnoYrGA8yj7fmuBmMsPnu+VahbJEybTKLZDQ/f
Owv46utbVCqVwDXM/L4DUstRpJtcujG1ft0yg/LbBNdOi1cZG60kgaDB0ItZ5Yxb
0Pt6y2KACLFH+JImqrA93sSgM1PLg5ydWmYouJPXQevOvJepGSNIn/ts+iGxA5pD
zrFmqbKYceGn9MdtyjLDWDbZkDdbhIWkhruR8dVOytJgs+I4uF/wOlcV1PX6KfTv
qvE3Eim4/6JjjtxSUWQIaajn1KyaiSD/PWBOFW4hWNOlFT3wvgW2M2LBBSW1/Uhe
Fe9pe8FSxAnmwq4KKZGy7J/0oogcAr9mwdjW2X5ZG2yI0d3ha4aiopJJtlIdkJQR
soLspQPiTrMW3OUP4hc+OoL6vm9qdhVguGKosNC2IPN+7c17ZfIdw68ySCBRWoC0
LoZo9Y//v9+HdYH1WysiXwmiRuANRXuRlMuzvS2Xq0Rm8G1qgUUsHXjCch2aWOUU
yhjYnUejbndeldO9bVcQOiKUXgjymjYiKMUQzMXgWLqUe0Uh1+AU6geXvdpzNb03
wRZRefoLaJIoz3pGNDaWjXdSY3+p84x/tHoqqNfSs8R0ZrbT22ZyhwQ3+LvSNoWG
MN7ez3TYBJHOLkV4JXqn533O8+HIKWNClPn1JXpfvDna9SONqeg9J0ZNkVe6Y60T
yyx4QIzJpNmnCW3s5mfTufCYfFNUpehyFFheOWlo/DRwgR3ZH/a60IyLSIcXWnk7
gGkCMIcSzlNud/CQ+B8HRs5I3edfANj/pIfWkBiwm38afa1YF12er0ncI7MSja1H
/IkO2zx4p1WIi3LY1i8KdtASiVyW+4pOd4owLqIVZSqgMaAElBRvLq95ptomh2Tg
xUa7i/LGRnyPY4dRamY4cVj4j1+Q9HaIP3wvTnjOHJgL26wPPfME8rtK6CSltmtX
dIcndkUARrGVudKKdzjllaMD8ytJKoWTviMVhVW/cJZClUF0kzob9s8oypt++eRT
zrhleaGKwFs2iK99YXvOEe6yrXx0LS4o2Uz/pORcHbS4wq9akzGgvMYUbF85qszw
MpMF/pVrb1p46e9TIB6MsuarKIPnuTVLF/15/a3pft/EeM01qNEyzEC3VYpuHLL8
30AYEPfcVyUTIApBlvGwxkyfLlkDGaZbY9mNoHwYpSfqxZjTZe1ZnwUMK4tKpY8X
Q/PpEjLyRsxi+YWTv/Uo0y4xAdrtWGcx4qKeVuM0iMIt9bcSCGIUXGHGcmBpt3lq
D3quYHcY7jz5hBkekLwt0iHVCbtyZEDfI6U/32vlJzYm0gWECakS789pahCQN1+E
2+g6B+6B+c1g23lhqqJE4b4huO6PfVkbBTHTncnlU/Xd+gWcjD/UqzE40Bfnr9zG
2gQXNvZLyvy8MFYfZjUp58o5AXIagK1js/LeniUBaeji7G+UBSIyi5+4mfQW3wVg
7pIhEDFVeU1rGC462EmSfN0EnlAvyXSzV4K4XdNqa/bMrMTmzV/FyDLJk3CiuLjB
kR4CAepMoBvtWJ2y9HLJa9QfUnSFO6bU6wjPZlLtVWnxfJME6wNCNUzld4dcV2mp
/zE22PoZnIYHryX2cP0mJadpHDczDJPNxsjblmjFBfXSDTNwjuxrmGu+MRMCwE3D
bgt6tDhfqG3jAuYs9lLe+LYn0/0zP7SQJpFi54SCnG1R7v2IN1+bJHQzXFB+BgT0
Q/Xa4pmhBUQIYP6FROoKLMwjmfebiijG5NI43tDDkAEWjay55IE0UlpEODWwHrFY
2PQqPppz2A6jX+P6Bb9rlQyE3Jcw1A1+DSexa5h9NkKbkiBctwgXpE71Mwl5tWJw
1ZhVDZLPZz8nRCMcc9S187qmTjEoyScgLXqi5NDva4iP8Z3jJMp+opnzjdJKTk9p
wdrYiw+5Wsk7w/lHpoeDBjnN3XXJOEdkmYh1HWOviQBOxx1fpf6U+iL2v55PbRfy
ziSnB87izjNRDsazixuVQyLGDhVMdJagcYzbsz/4DebxIALOks8fLR/DZneZK9hV
5ZD8IvLjfd8A4abNUBdcgbBg30t9MuyzsNfsTGBjQXbqohCnyCNGhtGEI5ettmJv
o6XM5FI2GeQUap67Rodp7cuhoFCpqNBChq0X0XEHa5AmvzVrDW2S4dqeejSjFHO+
+TnrmzxitJ7NhI8HeRG5cabmr4PH/hufSPETOhLleLDi327JpWKkNgBqd4RP1CI5
5PwDjlceMQHlCV5HVJ9rl14uBevGBw8veI1wEQeQi8NLa30RNxNpE/x6xfbvITqb
2xKhj8M1YiHDnD/hYV5E1uESspctsFitYgf2leuHAAxwbxhEdmbvM6TcURr87BjU
a9rv345EN10SgOP2XCGk2IvMDbH0aWECHcHhoScN3kqI1Y9aYufvQgvLsOFun+Eh
yzIXVOfUi2LKi87dWhCaDgMyS9EQ/CNoVoPBuQC2XDofOiv8b5pgrCWT6Ze1/3KL
Wj3/mgLFlmLH+ocG+VYu8+oRPbABeY1Vap4mB002mBldi1mtfJqu2f7QX79U28o2
FxpGVo1EN62hD9yKlT7opOBSFYSqeSoYrHqee7ACSEkOaT2Y/BMfuscCQT0lN7Bh
eH555/uMLxS851CQH3HlnzZIQeBRIY+4DyO9aYXorSp1h6BDgzvYkyPvD6crHZQP
weuc5m2RzBKPD+BVqGvtrH2ffSqrrAxBpExLCvp0CDBZqtKGN5Go7ZAiFwGnk/hD
9ZIQhRTkFXnZ1Xnw+M8zvElzL2U4cj9wcMmFNTL1pcpASr//cqQr99G63NMJCT3L
28dwD+vEiUuhXUYvZOsppiEE8eStudzOK7HvgcDLLj/wbtKUofohmAnCW2UgNWTZ
qS6bxrKzIrdzS0dSq49GnZjUq7XuE9k4k4LkdhExm1sUXzhuHNn2K65XCkq/B7nq
xnEKJ3Aq5zZeMm02YQ4m0jAiA+JwpQQy26GmNCnRvMi+DEnNKMwzfvZXUpRCOakU
K64jNgxAXq+Uf4FvJf4Nld2D5v8oIl1StrFaWDgUtkcOdGbe3QR56rBk1Q1MdFnM
9XaPQ8IkkdXLBp0HfZ4qc+PFcjMnFu73SpDFtY/SyADuF0yTL529+pB0rXCMs5QP
/dPiFsL43+lidbJYZl8TzWpEUN8+p9xdGSovKpSX438WHsgOJ85ns6rIw3Lp0Ul9
H6/XxWDGCZXz7D+ANW7LbecQukAPPSyblL/npwEhhD66isp0FWaDXoUvD/vSaMX+
XW15tfqpbGtxsNo9X5a1KktfJobGWmLPt0TuUOsf8pt1eCQvEWWs/V91NkdaTD+h
AesWWi7PfLiOrGGwqnTSRtFicPOcZiONWNytfla+3vSvXmV2ND/QEIOQjt0X7Q1T
O/1qBAdOt+w5vClbmPh3u3cKoeGgZnYOxhBRMFxpgxO3Sot5u3/peyelia6yk5CM
iDz0inBr28e8dB8/8IIUNMYaN1aoMr4RkD+m39E+pArj+xN4bpvFtMmCyRUcSmN3
tOYHhUb8f3m7GiXYSfGcsS9Bt6mJESl3dlTvN+d+oqcg1bY93EtP/hjNFkJFhRcn
58THsmMwbwJ6qVaMAC8TTHkXVreW5XeVdu9m0rSsSNPwWG/Q3eHNaj2/H44wYTfj
BYKcUNgMCzg+V9lK3T3zvb+7wF01TDP3FVG7n20VkuhfANCxkJry2KDIGtnrugow
Rr8DChy00IXvyHVpWsHw6Nz5ULFMS/3R6k91KbKbZ2WYyoDQDsD1oVy9mbL3Hv57
taAUmF79+tcuel+OUKATxX7E0gqyt2HiuH1ack8iUF034uDepZhPdisMCC1ydkU3
N6q8gvMNOEFs+tyNORdr1GmBTvqmucS6p7JHaeln5ZW+UzU6TEgNdM8RNjN7yThE
w3TzMn7jMd3xPpmCEG0BEqbIH0ifENyLyvteLJJWQl52/B09Hpy69iRFMNi3+wsk
hpkpNOXszLmNr6K6+hlcEOHAfaHJrs6DAMs12gHW6XsYxuDamWEELHtJjqF3wD+h
ll1tStD0UtM4ApfXsh+YFTvQlPrmHwRpgrX1oHprMySLF3pfz3DKuKGlCb1RE0rw
dp/DWIMOgeADq0Bt9kMooYxfgJEserHj4faorqWQiScp/oWWFVWzq5BE46E5ha8O
T67B51nUa6OTAViJYJq9IyyZBod3Fpl3zhic2MU5nFRLejs8do71pWWwa/po0e+9
iokPzICvMuPOSNDT8EQoFU2lsPW4ER8CxUhKWTKPYkWdK7geQqLDcxJ2xF9F241t
ndAXEKyddp/matsM5PFCYLYm5rM3nQ0zrBaEvKb2OSrsNHVvSFGAT0ysGr5poz1R
km5YMBPU17mHhKPednAPz12ajOfq5+cPN4keyv+Mkh9eZFcTwWlBU7LT87i12pol
PdDbWskAE8RQrO1GX0/mSPt+fPEOUA46KolIBsbhqjrrziCP2pvbOTYEx16Cyqv4
3V+/BRDpFADf4eo7qtvPM5soJA6gw5I0RboRiJ+F78uy6FLzZNmlFIOjXdtT/Q4Q
2/3hS0iGnoDSNt3+1vpM6uBZdRSkUj7dvUgCjZIflDwMes5BhStF6RHDmcvQS7Qb
evN7AgpsJh8PXmx+6W/L6F3FLYEbrJW+mQRE3RlGTYWbn5OmmdKqeM4jM/FjgkK6
uG8dB0AlFyJS5MtAo63w+AjakyCPj8CAOjd1yGF1+BWjmuhKN1mQbOXWXbtAytXE
qLVTD44rnpS1WOuH5MLYQk/X/EUl2CgNNPGLSh48PqL+Cg/cxRFWnDXupeKBaVBi
bXqUzqdW/KIbvgKBpZMmDjcIkXlGw5aTtaovaToK+xASnusJySqVk+APPGO8gYRh
PydP2MjnGzDlHH2pGSXZm8sbn2qfMiJ0bgPs+tfEeYYuobEb656ETYDCnl88r/Ut
62WDahN/J7pFsu7daEVsS1cbv2RVfdeJtrREJsTZCUoY+q4zRZjdRRJIST1iXh7X
RERlEoo5NVFl9X98ThI7nLY66gTt9n9H2WeXgoPN/dpZpg+suPGorTq8tk37sj8d
9C+Zwm8H5JJb83W27VEZ14kozhUpKrxIYzN/hkUi9BwDC7h5EkFuuV23JtTktFEA
tEf3BKOlSeVJ59tOI0IHCjOrB/a2QLTPV2E7oLjHJjHJPkbnnXeinVPuCZPEZRde
OkkpK5Con7VkpWxEthJDj9Yg4B01GvOmj47MHdBVdferP7Cq30E532+E/Y54uhxf
e9rQsuroEYpx2HASzMOZ0uBdCFEM9wW2LZjpazuuZcgNw5/DUb3tFmnVZ2ckgbhe
0qVU1Z7x+9G/T66D9M5dsg+n1rP6jB505gxqCM/trqCwmXAQmCPqJvGy49/XzJeP
1nprPkvZ4VVxciKxcuy0/wc9wD+R2wleHsn92o+GWODBL9OsHu1HmZPgrJxrD2tO
rC0iF9cHkay6ESmDaKYOgJmAgz9rfLioenx7qY83IG/tENIB5zLPyfmcbtng3KRx
JOJBRh4a+sdV9AgW7lyh4XoWKlA50cjQb0wA8EaMtUOOv1nPavO2qn4ob/pT9CdA
ef+S3pkxemRY+UP1rr0iERInRhtopTIwoiwDB98IO+WeUrpPXANcN9mFbWcTyYOL
9a4V/Qm2LdOeC5O5wZNbL7f3ReKFCWe7TTR4n+dI2h5GbqIMkbyoQMj38vbS+Rd+
+moarIpWvuzZA6Ord/+/WE6nqMGJ6kdcQLQv8VsyD8FVc6sxZuTsv7B3ztPSHiS2
nekX+M/sANY5d0/YmUeyaWS0xXnxA+2AsqoEj0m8CRfBPsGD71em+S0pOJGuVYQo
3UDy5FbDBDLGEWIz88JCKgEwyYJWgKcrt7fA4gAFaO8SEhuvstPz/Wp43UhfUPjA
GJ3pMfMsFViXLsDENKij6hksiNIgA14E7zmSXCjvH6WIc+cxs44jHx+92KDjHOEQ
hgeFEdn0ZAeKoUmkOKdex5yLOilqmAn7o58rpuJ6Ejqhq9t2ziWLtEHeoWHZ/KPf
ABvrxIH3nS42qTpYtbxEbTRNLg3DeO3QKTEH/ocyJ0E8Z8kcT+e62jOG+77OzhJz
RQUHOpjY+Ihg3ICGH76YsAYtAZv0/ZYcNxLYJjjbkPKnrb+sQM7UAZPryPiawXO+
cRO9c2JLq79AZJszJLk8viOdF72Uxd6n1CcKtFBStDphM6J3I0tQQcHPrnfDYu9x
/zpZGWgJumtEH+0tp3Xud9RU0ZEQ1VQ/T6zsjr9NCs2eRQgYROVNp43gu+D1jcf8
yImtbE7I5i3U1Db7BROrgjRqIfyswZ3vvkBTcHS01ctNqmtyhSlMnbCYV+dKz/q4
u1k4K5rTnHcaTdji3S6NIpuUS2EL3f/wSrN4G9K47+UOn24kpNWT1ZgyFIM5f4K9
Hsye49CxnPAQU6kbjpV0tTSxC7PqMo6ppbBrQoJdv6jjNcBigfpZCjibbxfiKTvs
q39UyPZFW/VUhJhzktTAY1NLvU30GZaEVkvQleDMOIOCVTT5LnHHQTVI4xWE6KvH
KV3v3mV5deXrGIZtPZbei12FBigtDKOIrPCsjb2rkRaaOubxId8tfBXqr3R6I2BR
2bG/T1jjDgTx8rtDDmjW5uFGi3ebmQPQH01W7/dtT6kzyjZY9SXI/chCjJ+Ous7O
wnkWJJ9cczWdex7i0FRfzAGF0WleFUcv3KZOg5qUkpR92J95rIhVcE/IoD2DCvKu
XU1xhI3bULge+aTVG2eGJMlP7wn09B0xsKB/uIiSy99uHw5liAqYMkHEyiJ8I15d
w+J3Y58QOFtjppImSA1uWav4+fxlAr2L8JWD30bG2cWfbOF4NdocuP8mOaDMvQL/
A6sf24wHzwb27j6l/T2VpXjbrl30ymP+EXkBayiE4Ztpvy0DOKG1nMV92r+z9pOo
42zCD7f1zidMr8Jht1TRAH/JZT16Xxd6iCRj1RbR/q52Pr6G/mIY9lXjywYfAYHB
rxy9K1VutjrIRZmJoekX4B0EUY62Ef5m4rWnUyF1dKMadVwJPUBNUDoOMGfW/gGR
Qv/N19PaKHB/7hrTWlXJ32k3BJS7ho3BcbQxfDAEUEaN+cDhzFMWqGBJF748l7QP
/Q6O47Vi6Ql5elZhcCGJ2flCLJXxaWEAQvARM5FVpB9DtQW2OD8JIo3GE5AP/3gR
5ZE4zVZMGr209hHSVSb+CB7cIAAUqdTZ5h1nWSKBkK5BYmktKCXRhyQrZsHwXmk0
rdaCrcUidyKnyVvmd3QbGKPNHISauduYtg0N2HhRt0CPOzWldrDiasnugZ7rc0TM
NFzrEuwuM4vjO3TxpHUeUTqcSNsOSqiwbDnO1QnhiG6J3vozX2X6ORfxiQetWu2I
iTaERNWq68xNZb/qc1j0VXPIOuTna6pa8honkX14FB2EPNTFjNipSL8r2CGSB+c/
gB4dPNzTscRwkAbyOHOGKwJxGBxZTLhv1l7zS+9Eg0y6WLod5OvelSL/JlTptrUl
SPyHF4haKk66GZzrgiGDjNxzFkBZSKAnkefO1y84E7dnJ8qMIsaifsZKYoqfFSMu
Evlt4M/cgLJqedQuYquUOjhTPLtizPy75FL9P+2w1hCCZ20N0+vywYPaVa0OzhWx
WDJePzdwbxv3eQ3HcCNFUaO1rJGZcBevoO14jPRfw7IUceieyar7jfTk2LJMxey3
u13+D1VzgZfcog7kLAwECgGQq82p1JFknoY5gztsCppLJsNRJgpEnU2VCvRCdIXI
O6JGA4MYHoCChwmDjA5WVvJu+Xb3h/ijRxnxaoy17y+sCfbvURPXLTQsOeidIn8K
VaUye8UuPhJnnDdXOYJN94stH10jQvuAteZ4IQO82rcRiBXmTs2lWykoNeqDOuwy
H89B96gR9SGAXO31T5fKtIyoL9VO6851u9vBoOk/VqL4JUZxlf8ZciqLpvGM40b1
9iILHQj7EZaoQL981jE6kcy+oaHvgUa5PAHA9ewbZPl3YwAKBdKSA4SCbUVfKL8B
+u+Olefe3ZTBNAWq41s6hAReSWdupmqx9K3f0Ja1N8sGWxXUDJXllG6d3EYpXexJ
iKP/4+g6JmC6eYJIPluUd/iCF6YzxkJmhjYdhTHrTLRo2uNDu+gqRocEKPSYb1Tg
dltLM7DhhjYxq4u7p4AM+itB23QaxaqDPIzLDE/iE/MsXhLFRPrCa7nFlG50FLS9
OVIiViFTU/8Bzzlx5q4tH6wgzPzBNj0YHJn7ydrn+8YoJx0yfcMGgBmKXE4zx5ky
uI7/BXkK9UBYa8pi8o1L2jkVRzzhFj04wfHeLtIsbjA0PU0gk0LAUpHU/zrnlU5X
yyDBOBIgrje11mwm4uS01jeMN5HonHN534yNB6vanWZU/Yiwlagy+8O+XvFVGxI3
hR25VuVhqCgHPsw8gLsSDNwpNGVEcE6WKOw0CTqCw/H2DxltR25ILGCL7HSfRlI8
Ay2s3gNMx6cDVI8tcY42X5fGwb7NheLzaaxQiaTAiphGgHnb9+DkrX+BG68Oi11x
+8RCFqeB9KmTqyMV9h0AW+1EGpxL8TjkpnESoUo6Dsu/tkhkkoL1o+LADbWNzJi/
P55Cx4h0ZS/SuLpSF5Ms2KKlMCM2tqcPwjq/cmJXc7j8Tk1dSxQE6rw8Hx1LG97h
2JbF4/05l3CRjmtzwP+HzJ87axDeeRDmQLMGZ51sjz86qz/8YHbFQ449sKtoohmQ
xvchGT8Ecc64sOinriDiV3MDXJDu4+Xg6Gh0whZlhmFyVxXM6FK4pLkYtKiZkiKW
Dn0RO7insIXAhqj81+GuwxpZq1cuYWW4DM39BNROtfU7ANHM36t67CFXbHVAiCAf
0IEJuyuvL06rTtEQ9isDy6yV7tg5Z31jenubSKOCEq4ucCkDDx4BedxpIUlTTlrl
iIp1kteD4Nvhu9sxnEd8jMCr6I6fUy9iEksOZGhVYgEtIxoU9Y2+Iot6P4K9tohq
JyAK8c/R8D6y4BONLCRLf17vCaBiq5DN8Cia0KTTnlb5bwPJE4tYZHzHmEPrlb7N
r8UCG8L029WApU4lwPiJNATddrujE22U1yPUn5FyI9hoH2aCTX1EeBnsLk3Q4o+a
fkxaqdlRTKX7028nP1X5Q2CWJoYYWGxvx3iCbvuX3qL5qZ7oQ0OZPg7arm7pemMA
qKdMScYJMjffzc5CII4QVyj6xGKmdxqt27n/IGh7clvDnK/JQEu2ZCXjHNZOdzvE
Z9fGwGGIWSN6dGmcmtpIPASp+qCPNtU+QFgS2PTFyiVqa+XrDsXKEk15DD4t+EAp
A8Ej0ebSPKoRH96EIK6IkHEfpwDN1HsmUDAtEEluVvlwiwNa7WhUP8Eds4CFmtuv
8N54Hsx4TlbKCECBtLdD1lesUTSG4QhQDfhvwVwp3mw0Wi7Zbwvf/EI93GDVryZn
IIaS3UmU0mEFvgSU3hU7SH7nooSxYMLPjwZ6I8deFGqZ0UyLzLiK4RhTdEk37uUU
uu1krJI8sWdUjexnPgEsbuMHJFLNMZJ4eLtxuA5zDeIdNIlvATetwR5jbZPJRgj0
PogbbIU1ZglH2CzMwdmbr1Jrq89C4xMKlBQ7jJKIAw2+gM2vpZ6D/O6ueIQSH4xY
4ss77nkmBpiFhFW1LAGK1dlT3Q41vgEM+AJZ8LpM7Re/3bf8uqI9W86hFW9zUZBt
TD74SGQNuJcMaEww3ayim1KgIjWce6YoojXl76d/CZepw+q1uDo23yoLvVXG/6OC
E+SpWd9UBah94PulNbqqOP3LOeXHqLKfE9AisayJ0+rfNDNqnHgXTzPoWg+4T9l/
lMVB0Lpky5xqKL9lPOqH0EajWA+jCV6ywyulfFz7RDPMV/Kr1iDIl8E4RhCsOHOM
dGxwNuPcYtPNio4CBy/c7NCHVxhta5yy9np+0KWRgaWB4TrACD26idfmZGSIlvr+
/yXL6mDn1/qWnBI14cguWgtPeYvy3+EKZqhRlw44ysDdmeITz5IfK8Bo6IfYXLxC
T436jep3HL+bDP79XAzXnL3rLabujICkJIMO/xt9H9E7wuFipja1gA5C2TKamJvY
8igHEU9V0qQpa/+S06WhW93qTbvgKf1MEtsy5mOCaqf0fTHalbZ4tBR8OnPZIgy7
wiPRLAkB3l9ivZIb0za3naWj+/XJ3dyYOuBQe774xfB4VD1ZziGBQpKGVr0y4Al2
0Z7B61kRA0gM4upY7iVyQrLY7IEnR9Jl0rX8I6q8HWlsHZrJQ+r7ry4I1wQhVO8P
xY4iGWXFPc1VA+9uXy+QL/L//XEkVvz12/VDyCRfnx3YPKeKZdq0ZymzMDXW1Goj
VOdWTdATQMPagUf/bFzbppzjOCUfGFPb8p1Xla+rPDuDACVLfAzEfprqndn3RepK
4BJhCNUkFi/TPKmBH2dm0VwJwanqDuL3CkNVQHFZE6i6D7RtFQ0jPEWdJv0vFTu+
zK5kDiqWoQsLabx+C4QOlOe8YfQSJRFWdNUhGfzjK7lpR1+5h9IWGCB9gR3aQ276
nG5YgIpzs8bhXmT8H8wbXZ+mBX/FTurExqLvUMB3hh5DNEkCE7Kc9alP9PhYeoib
N4V1xxMilotjbOCMmcn1zxMi/kQkEgDg6InPDojgDIxZCfUrZ1S6DI9l6vrhIiQ+
0Su5crFcwEjSiclFshLrxy1GUGdhPKFHZ0sPs8qFBNySSnv6p5uYL96MagFWGtw0
4xvosfS1dgLwsyG8KorlgLZMLE15ihDEyVboYUrfbP5hfs/noU7Bvm52uJILBdIe
Uk1Zb+7QQwVseeDNy/+om2UHkPOX0OOOBzlgDRYMmAvu1iUGRF2ADESDyXyoUTjo
kKm4QZJjScPLBCp9b54km7VeCIVu2Yhvv9ODf2VYD5sLnZEDd3J+nSE7a/bQOLu8
ISvNUg+s+uvZJ/67N+Psgb0nL4AXWnyl2h5aHst0E0W5fC5Ut/NhYE1cELGFPzBj
fh4+ELI1UWWnOJaMIaHYbmDjjRhsOhJ21WmCNJCvFfhy6Ue5gKDqYX0HagyBPAsn
MyOJ3C+H3AhyOwf5wJwpo/doIrLYq8AbqLyGzwa22vSHpFlIX2+hIe+gv5C3GBKi
KQEmm2hDrzwUKC5Y0b05sUyXRTlzp4pBt4NnVoJbzUqVM40a8oUyWMHjRv8XWH/I
PQfqK0SqSbd4raLXNsc+jiGh9LgQUJLqzfOv28QGPunVtJovElsKegeqoKPR14aA
vPB5VrhTHewcam/gQwJ9SHY6G19ul+lg4Kmawn0b9MFhL/0fgqDyFNTM4L6ceQDx
Gtry3cNU1Ph7ndSOoQqPBc2LIHFZe5lPGpAqE7xs7o5FIozw1Mb7VLyfiGtrFYr+
B6hHpt96iaQAhFRq04iDVPq6yRzdpoKYTYGm4oawF9jY3zYhq6qP/FO9cXm/nfsW
I7OUWyvudLJOAeEvwaHYgYz+0smPNaGVCCTk9ZKDDxnjZVzlfBDvWiB18NDC4qaS
brRUQ1wnOxaCevlx8tEaeb+N0vXmuQr1MYqJtwu33NhuLAC3Wx6AAGz2c8cI84m4
8ZjQ0ya/5qyuoz3cyStufs14GfzMb1dqZCe/OLlngiwQKjsbLIXSMSMWWtIvOxa2
DmiiHdOoC/pgVx3tSeiBYkRi8qDrsdxVUHN2MEmKGkizXe2/yXPYf9DEBRhnKZZU
J7nJ6WrS1KjWAlTMs3bO5/xJwqi6Em3a8uoRIp0oJXaUDcqbBlpzBwJ+tWqbCvMs
Arto1fngPsCfxJtHfH3yeiBbsINX+nfo0gqn8ACPjIqXoXRjU3iJDcD8Vzc21VpY
gx+PEnPoJp3TLQqcBUnltaQas0VvT4/TylNxyI2UeFPSP4y+JPnNcBu7wqg/as+p
LFi8HBDZhbqtTG2ibjcSgMC3KDagB93apT+C5uRg0j0RxQMM69rgNp4bo3bFOfQP
hyMgz3Nio/+XSPlIMOiJXr3msja7qXobIa1RJScvZj4sjdppQ1Lp6DSXnjfm0Uem
0s8dPshTLi1TaSDxPQAR7jarPje9klB4EvQWncyfux2w75NoSIgjdVmVgqkYbjUI
5XKE4o2s6TzufaX+AtUb7P98QHj9OMX/hf2nvjCYmQ8KcIrLMc4azOaQcpuIw0KI
4C6mTkZRHDM7x5HQj2/KTEnVq2jCcieARt2/NmxD/siO+bmjA5grK+9VP8vTC5Vc
gnKgGTkPpoRrAoMTykpaMvvqAg3DGseb9gNctz4VknGvGkurxxB40FLHc98EdiQw
BIHwZRzAyN17fcq+2VG0OWrl8Hhe+BZo9yFCFosZjW+8oEb7OOLmtoWgDCHveSTW
mxbttXLofEd2TKiaW3th/Fb0Y798cpq6WUX/w8EhruDXfjW2vdYqhyhBTgIPF7Bt
JlGxxoVrEQKRqf+csbfQ9eojlyBZyPrHAYvf9YTyRL+k9RMt2VG2Q0yXdzAyMHik
QO8X+xa2CISbsSpCkZsWMfp0Y32GdGsCptbycdaNF1vqdy40MOw4tNM4C8kme1C7
WSGzyT4pX11SVGJs92J9TYXxTsOi9aM1iWWOcNjuGpsq48JfClAnUc6yX+gJVy3u
8QUyGZetkJYbQQpRkBu3+N3UrSHooTHNHqGyIT9UlCNT99UF9wgGl/yFnMWdAJ3d
iQ8CsrSeW4QFRSx2QBOc5Ax11wPt/IMrxW1Vx7PrxLf04Ye38jCLpwvQIPlYeUmq
qGeWGnVHKSywR0CVZ5wM4iJldqehrcmMboRm9sR5w1qhYKA4ktJ5L1MxgaJ84+SK
JatwMAtWjybWPcTdXqZ3jMGONLI9dYMZK+UGT9x66XoRFxgOaPpazWvpBLvexS+i
KDAX+HE9OAUt2NaWmUn5WN9eQ5DXj1WeWG44M3qUw7JsPyBAxq6qn29VLlk6fB73
3uxNPkJtYlPAoLJzNiqfspamjcj/tLwRt+LuAUylMXS+QPzqp0nIoKmeqj1uXha/
uE063AjdMueWkgvs1MyEWmhTZFgiZCiZBcVQbWSnwMy/gHHhwhZJRdPafE/qF/mp
R/wpL4NfBhUNWaHSflqFv7f3pIR2XnpeXah+ERCiHr+OrNayYhicQVfMsPW7hQxs
rg5O4tSHzp5xvo/5WAYG+IgKBiPhSV4dDULXAz8m2tNpLcg1naI4PtOF08pXa/4t
a+5LRHN+kfSwniFw35Z/20hd6MTPp+B7uHNQ24WYmpT31K6k/SxpKnipQ6jordQU
+WY8TQcUTZsEqxz7PDwUXfnuROrPs5VIhGLeiHzSunpOyH+YotmMWQQKd9oPnODA
FPUUQix2nfA7oVMtl9KzUjB3xGplWT+78Fw5IfCaD2XbnlD+4DeDo9HQ61KQaKV0
sY6fYxc7tR16ckHERSvfMzLMUs2VOwkgnVlGCTOYMvsD6jwqkFHsrCJ7BWed7MPk
88lDLuvVugrGL+SuFJlYqEjF8RLASfDMvP4tkFByWLTD+79YAHWfcli3Aqo0iRwT
gzBeVcXABOhZGElmyV+wl9xDhD0KQQIKCYYchLLqmHR+TzGp/oYglZHR+t/sSXtM
ARTDsX2dl60G2Z7fwNFgZLSfoNzNjt56FvO9HqBrbD4v742tveI9fCLOmpC9/YCB
nBcZ4/1hQG770Sw9JWn2eG2zIlxsNYT+lJq/wC5uqbvNQfcKB8Bpy0wujEzskhrZ
mwm4mtYq1uufREpxRtSl2x1y30jvZFpMwbTgUWxNPSfBApLDf/u2fcOxU7xJ7Y6E
iRdLM48LlQEkbn+6znE+12jgyDZ5A1EazYA4bRjV+Mph+xoRx/JLAer515S7E/6S
LfC3JAwjHH4buBPcpW4UFE6HQWoXEJcAO/mvovFPDEsjGQ6YW+PRAPNojZ5/3Rj8
m3jPc0TZVoIfBhxnXYkITIDH5HQpTOXzSIGdrRGUdW8xjdYWywOevXNkQm4i7kH3
d73eo/N0UlzCX1Rprl/gAbIN77hR/CqZDejZ2qevPSPssWj+KJYl1JmAQEtPcDwf
tzp5G8T6l6kqvY+hgNlnlj59Ik59+S9YYmLFbKwqzx4cmNDH5o4eTz+8qXpyPfUC
6iRpPmv8Ws8R1WkmNtd1vlVeL997vbU48cDmJOvOXKLzHtlPJW3tYqfZXZ7IVCUK
aVUlX6Ov9EHvSk++LPxvZbZs1aNuxKU3qznAklqGw+2BLBkiSMTNMRBLg8n6EROE
mI9BRE7mxQEvnfLypsmRDO4utj/MFpfalgNaOz0a6ZgXp+Zpg7fBFxxNxSMzsPMR
nsMUgBnWLNb7fOhUI+zFfteI4z4wqDSHG0Prwtcu4WFzUlCKJftvj7X5wQ7si7JR
atn2rMpLMCNkRcbRyue4Afwgapid7pe6kYBIWN8jz/xtFk5hrqvQZEePUbEC89ae
R4KFTKdHOtrGQlGhxnl0GV76A2NZ91r5ReiRPDCg5Ja1svLXllQehFtP6E5i4Fa1
hk8uMJclOf+kEtxOPVkmAfOU9WWDDZkxhU/uvRrETvImT0Od79ohGesirILdwSXu
lHlQjW0fa6yTH+cjFmiy5KdkQvbshDL4ygAwd5Nrm1iNtuhYGWyB3GmhOJqqhy6w
Ag/gIabjHgIWg0+8Nq4ln5Pgt5FjB/nerH15KebUFqOICjObMRH7cf0KeV+eyGI8
ewCrm0dK94Gyl/3rM26Ec/4yEdYakIumC9re5wjWedEeyQ91vceYuv7x2p+kIxsf
GGAFFFCQ6SPkp6qNglt/7amMhMC7nt++PmYjNHW3obTLN5FC7EBo8GMHRSCkV6nn
nwTlVTSw5C8QJSztMR59lgKobSmUU7W8ddaJRLaoJkaoiqbXS1/1xwChodaS13RL
GcmfoguN00P/DP3hnN98J/Y4CMU4YG6+4/dl7Jqf2voacyI31rGX5E6a50hEgl0z
LfpXWRQbVYK9kDr1cV/TCIqxymMn6hv2g57fOsAgsJLydPCxP5mPRCp5cQVFzG52
n5FkND/8zRbYtXJOVTJUEsO45+4XiwDA05XBx8mroXchhf4I9LDGF/gKzev3oPBF
H+VaOtMxI2fhqHKe3evOHMbUKJQxd1IBJuH5bnJtWWJnuDSiAyX53uH2Eb1QZoxM
fUVAPwoTh1nEjuL6/haB6UkSztuzi4SvbbGeozoyso7nHBXYCd7oGSG1k+Bll1ve
R0aQ4JtpBYnY6fWRZTdq/aK5rIGDtV0zDXEjYxW16mDJILu703TqBtNbAlIUaWwW
Djl6gpBPcoFvOE26ywOq93Wv46u1anfY04No7by/4Usz+gO+7TeypXCY10Uz5yH1
1QvYaNawrGDU5ZnCaVjpqiDmfUFvF7kKDNTmZmnjm8LHcL4FeN9G6RYTATGLPPZ5
Ri/R/BTKZoqlWBdm869K6loetp7ZmrILbxHyqGfM81a4gtMPaDxcmeLPG1yIlsug
HiElajPFkid6sT3ng/+NUpRyBNFHKrxB0KUHYcWd/CYR1f090QNj+SBnIegaR4T3
9zEtKGCWYOV8ImwnJ/LrmFboK3m9YKdGueir3B6IWg1yb3FLcNEiKMaCG4lJ999C
Khff+c6wIUUTTyed9rV/bGEem8qeE7lPVQAFSLl0WDOx1OVuW/UPN03OGqDd+14q
D3adTCb+1uoCwCaztAA7gIQE7+10cmidlVr3pMeVnl20aWzovlEOybs12SKrJ37q
lZErXwiR7x4xzTZMkSfmC5gj0E2F2Fb9BN2ITNMd+KZJer5CMLr67t8ooJEBQKpA
153nI1GKY79TP7q+VvKZ/4SUnflCo+31MZJ/We/ESLtXlVWjQmGD1LF/2GTRn+p2
NrvXBl2GRt2v6ZcGSc/B26qb+5HqBdF2HPHgbjVAn8udqpdRQde1t71vMGAAbdl+
TecP4hyXngvs/r89Hw8XehFdM3MO3UrHYp0i8M6OV9V6mMyTyzIPbWNzLy27Kl1H
4/uFlkSRvihCV4WahYzvvBU5VJfNPIQLICmUqk3rTktyIc37AMWtFl0yq+zwjzCu
uytjxTPAf0GQ04tgyInfQuyjrTRLD7aaSi34qReeEbSWJzS7f6LTClOsLF3A25od
FbfWdyfEC2XUtZ4Twwkg6yl9mKDKk7GeMk3toxriRhugtncj8/nxmPRRCQ7bu31V
lQyxeI/BWIoU6fjpccaSmQg0F7SAeLlRP4wXBxO1vLOWw7SA5SY+KxtO341nlOL3
91wSLFbhEy7jrWqQ4F1SG4xJXWXJiGLCvIobPWe93QzhxgGJ347RnGwWOyaAXW4l
KFUxEUcYfy/LnBsf03up14CET6Orp3RYzZdh3daOWiGHxSQbOPy8GVTzdOuKyytm
90qyCrz60mBYa+niIokTHlcUHgRWb20N7jcEVnU5Q7/P8g2zp1x2zLttZS5Iw1nM
y9YwDLFICNxI3KQDt1pBJf0FN7NWJNHfr8ajVwHFaD4DNw6omqOTcTaZUOwqWMz3
zKvR1Igj1n42nmhWXRjpJAcjwEOBkCArgoocr3kkZMfV3wI6YGh9hg2IPIcciv6L
BCVhSLIuux/e81XCb7S1ue46ANqMxNJymLdporIp7FbarTDte9fZk7VDaBVj3SQK
2+nto08lFoKU0lq95t4KWrOsaPSDh/m5WoS1FFI/0n2Rwoa7rQA1TQXO4+3rRu41
mi49UbSth8hzY/IAfcpwlBwxxvUyPiRh3ycr9DMNs9l3KY0Co1Yz/+oqx1dfgkqM
5UjtIjsZ2dM3pLLr4XqJmgsC963jOfs9O8pFHpJS6mWjNybE551l3sgWUKfg9w03
WjyApwJLykCpqZUcUAW665U0PtuiEUUe5bSG80yXbqUu9C293W2fDcDmJrE0XD+z
txASyzKJ1qCd9q3NjqEBdwmuosC9k8E8a9fov1KuLJ+1cAXSo3GDzBLU7EkN51GJ
vASQOiBO5hrbOXrjj/S0h+cEpNJf5c2Cs1Fcme5QvDn/pO2bYv608kxPCuKmdLgf
Qh2DJ+ix+RX+nvXOjjUBfolGd9DIicZCyShmXmEdBttrzSDNNECMBGPmRkZT4V0+
dptm4w7yNc+gC6cBDpswi8x/VrAe/haOYb3m6xXGGE9cqJ64JS9xqt8VeiIMU3I9
ONruT+FzeZ/1VrwoIlFi5rSivSIEv4QjKgjK+gvtoQvBvPdXCxnZJ/hfiTh00ixy
uyxYby12n69jjoMfDHuK29ALBjWMPnBvwrb9t8LPzx75VhTmw0ZtpbjiCnjthpl2
kW1+AgQCc9vlKiI41z19JDcyP0VzV6xBpMAmpdt+lBoemvy02GE4XZNszoS+4u1n
9Vq41U2V1pEH+tiKwSUOSRuf+mMhBV+a+keEsiv4slwNFA8eMK3qMS3uvj8+624a
I7dVdzrfIYzDHNqjAnOt0hVGTUsXyFUNn3UXhIA0NNooddpXBRl9anhv9lSHc692
qMHjpkIbMUcIwzJPW59aoH68slfePQV0xd4bnSh6GWkGjk1F0XaNg6I0ifeqXmdx
OXypCkAqtjQHsd2hXO4mwx+BZTcf1cqviqerhhzxc4dnVfdhzfMaKc6goGOena4h
4vgX6mSNmmcEcik8EGeCGGP8XbwNgBGNjU9grv2rEns3VDsqvuXrvnWprYSkfH59
bJUXcIgRRG8ogBxJImEhd/iULRi6rPWFj3TkQ2Mt3cxJ1Ky851Rp/Ok4lA5Y7Do4
yKb09xasbrYby71tC/A6uhjVcI5ddBoN1AXjMHzXLhQZ56jVtzphZmPBtcxVvWGS
ZMJLagu7/K1Z21Wyw/pP/pgg7T5f9Qyuv2FLTHujj5KY/dKrC0w5pg9ucuEwAcxV
MJBHFSoX2NTTacCoPV3ID9rOxKY976dKoNHRAVL52o7vRr+unGX1LdR2/k34uyXd
zzghAlilbV+En7SwrCPMplTTQxvi91k8QdOaeUjHgdPZRTPbDW1wE/wKyjj8y6hH
mPCUtPSjKOlQds/5zXHABzz++fq06SZ8a4/DIP1J2Zvg2xxnl7xujKjW6X9ARd7s
hE6p6LjElGSVc1zBlxVg6T4lU7zYxffLrNU5aYjj3TfywamATUB1QYqW3tujiwen
HXEEgzyCEZ/F6cimoz7ixPuEzW8b+AimXIZEKUHgWrcY9oyRnZSId86SPdPGIQgh
t4mI9orOt2c06ZVZWfTaqxsr4zWum1fh/X5Jh+kPRcaMda0SzqOwt1PO1bfnPQdG
GvYZeAnNNrKxX9YYk9b/cz2OmbapXt+HIZju+tLc8lG5fUnheLhk1H5T0TaNfJYr
mWNFm/Q9G3GcHJDe1uq+1wghBexnbpRdnAuS87BzEyzK34f/s0EiIP7Lip0/QQtI
g7ZqvCNrwXjhRwGsb1u+wxRgNUDy90lrYdgy9EUpz2DZQS/iwNfeaheopzIjRwhD
S0e0HpsFbpg0RgpC4ttK64PG4ZPIOmVmFM9PSm3aq0WlIu8ilGz/y0l2JGAr92FI
rJo2HEqhHVe9JOm0QKsTB/XG4oM5ob0+C2hvkdtMQHk/Om0oAPXw+nxGIrNuAp6k
3p2bByeI/GPjrGK4DA8YsM5KoVbfsi1NwngzgHDLw9Tlu4/hryiIlZXOdgVoyzQJ
Vd44BSnLh2r5/PDbB6P9Sc+D/gqtYRVY/v2qy71aJiQAvxc2idoRhQxeVSLO8jGg
/6Bv7k7oxC3fCZXFb2bHdTTvDCDx94CaaUab+gjN8/vuyIdr8OmeBj97nW/Jmo/q
TW5f/Z19E8Kawgqom4hTxn8n5dlinSL8sUP9FYyFVkAh0/DK0HoIIdQDthGVT9hu
eRaWkZDO1dr9x405Hl+yCSYhZ9MVSwBNPq60UAq5+k+eSam/94lwvgn63Xhr4CKg
iQvI2G2b0lIvrKfkjEDYouoM43ZjEF3TzN+ASYeBleLizGzkUzt/MsMlOy9bhoUd
8o2IsAif2rWPm/9/XzF7Xzo3tWUTTs/EuUYgkVwX0sFh9YS1AsUa/CBQyO1fpA2w
tIMQvb2VFbgevhKQx4qFAFcG2elmPyjd0ij5Vs7ZBaDNJ5O9w1CwS2r9Bq+QhTjp
CHnvq8TO8E9mDe0AXkWe1C/kdUYyhhZ2WVEJ4DK3G1JvUxeiJ1UBRqXev+0sN0F4
OCyOCkpQkqU9ROb30xs1Mbfcod+zn+LhYgCa4DYtGyurFi/x3+mI5KghaFT10xZP
GJU0aZ1I1vpPTQWWXtu5/MOP0DEtMlqmlXTuiCFHdR8ZaA/Gh53O1Q2Y7l4a/xCq
vf2bgxoiVF4xSMRnUZenALhlh274Ii0p6F2M1rX76N6P0u2YAqZ60EZk7C9zcoKJ
8Ov1P7YX8z2W4FKhAre3WdLoc15Q0BIDHfmjjwLwErsWEMUOyD2YmIm4e6nw3MNR
eOuYicI2TbTf1I0Hx1xtzg5YF8kYNWuOdW1XY5HTDlFmO1yquvHeEpcvBqY4mqna
dW/dr3wxEYVVPK0k9/eoFnwFuHJnPJeWR2tWouA+ujMGniVJg9QMzd6QJdYhq4Zf
g+xMOn5XotBeCtW/LcLOVeahLPtb9NgWTZHJPCOt/qvvnn9NO+OmryJBd4jgbxsm
3SUzeGXZyXjHIW7h02DcRQZIbI5yv4h2wlTGd/91XXWhBSipC5cPhA8Y1pAFZNOL
h8oLG2WEsZWQmNX21ronYTxWdZ6PO6DUTWYbcAZOyKuRS2GWte83eKJHHJRrVHxi
e5Qe52yh3illoHRbcE+AtsQaMM4I0K+2tgYrFfsalylVaSkKjKuT1aXHXunBDMay
hZNdTnVQpa+iR/z0NG5EzEW9xkaOqRoHTqu8j5DYLZWxsmgYEsHH7B7jiLewS2HS
S4zPUW7WUKLyU0KMAw7+DLAr7140amTA62ITUhc1gb4chzKoiQ4TtHqafvkOX4e0
Wme2CqZ1WVeBRdoFUA631wbgtU6Sw5fTtAY2u/y2BCkjJqJP4UmXiHxLb6eoB1Ze
tR9yN5cTS5mLk+tytnzGmdGtqGUj4OOkNqDw18NR3MxaObB/EGnULpt1N0i1D+RS
ikjYoys2uHvBWHphmy5MRZwJxX7u1oSk8pAMs2+xgITf5uww1MIHTRq2BS/jVHfm
RLKR8IZSz7gkDY5LBzAN9gCyZ4U0yMAA1+wxKqGNGH0JYzSIzpZqGRqCfkVIDouZ
i82peNzO0kRvnx65gj5af69dBkPkeQXp2e97rawB/q4A9sfn9hJQflu9SKY6ORas
S/JundDGeWIrnr5PaLZIXvTKZL58eeMuB6PLKDlOLrUP0psFpl4WW4E61jLQ5JtW
cWK0sO9wvXp3OEgldqkrrXUUM3MEde5t24GBlYBnH2F76jJct8oSriD9aJwy0R9U
Abds8ZVbB/fGImEpYeMVvdRBbgMCdULGSXFdO0XJ1yxQBIbxlAhDCRIj62yGwsrD
+J/RdOTD4CFXnALnw1cbPGDQGx3odaN4KrarYPv45eVqONcPk6Qi8uEOCJAWUSu/
gR1wxCaXghgV82DBK3WuumGeVJw82o5lLAgd2bDzWWTCRH5GaV8DpxFcWXCe/Zfi
ud4TBTLpxDTxJ0uP2QL6zbv/m1o/d1Ds9/+Pj12Ie5KLB4xJrAU1ombM832JUtkw
hkWOtCA/JT0wJuUEYOvMwhSOAX3xkHFSkFWHrSr39k3NCgDj8KB2pI/PFpVF7dTA
S7+r9Eze8ec1Zuvn8Q5xF1I3S7lKeugS3RRPXd+Lm6dIH28TBx/s3TBXIvqGHwel
544Lh/ezbrowk49JWqV6xY5OD8iLP2VP9znaTLQldVd1gN1lUS8tiQlUMMIk0BBi
1qU9+BHrWj9Ij6UwMWGdJcoYcYRbUPXIZ1JuN0j8mceLI6QbiQItYxPRU+UdsD2S
mKVVV1H7ExsJqMSFbPucrb98waYDH/S0ybcPuNx/T4MLHpViB2Tpso6ef+59rK7K
9gVlMV5abKty56DriqJsHLbgT9t0Gr6ArjdqnhQN8ftqWZXueMqM3sjqkqmT0sx6
sJ29MZXznbd1gacJuAuLLuTmyBQdVyS2kR+aQMKMO1h7k0Y+Bh4kpxKgScnu5IZh
flMdOQvU2xRicBElQAvzjTNKC+V+vwjKc1vvQDt0uzZlT/+vJoMfAzbrzqeydyTB
w0vE77+82SEOc5U01gOzm2tsHTN+dH6GTUgl+GZdl6KqDWsvL0QXUtjxYIDYNqeU
E+qKAXyRWvGHowMusSQvCvqqwRN5dBNpHrkWuSGGhCBqMS64+oilFPSe7P/fPQGt
2L69JqClyjwoMR5NHWDvcdTBTfXyJRfZ45t7AcASfymYCOg7FECxT1GtATiNMuh0
3J3TnfY4jFOI/2x/AkVht2jJy6QW/WTff2ehdFC7gP2X3N3uYs6eVxtDxCdV9Q6v
zXLFiaNOe1AzLUxZm0ELu+O1oz3KNOo1pngnntdH21BNW5GnQXB8s9qBn0EpMWEk
Zle+l9qjM+wPuB1cEaACWv04Fw4MdoA2msmi9FNz9vfYLupgvjodCzSylbenDgKx
EY2O7yjtNoQoV9fLN5trHv3k2Yf7xqVCfXNQXDx35v/GMakZ+J4VrC4G2+6iQCne
P2+CgFtXKhSYrkWN/G/550IJEur5gI+08fGGSYcBBXRkTX1BxE31czstT7zgWddq
pU/qYk7qhi3VqS832lJkRRpy7vwOzexk9RL3MUZFB2G4ewmlctAnfCGNXEAxIuap
57l/9dC9ehcJ91HmT3aujw4bgDDt3gs3wfcmgnHdJl6sjKu5UN2/qVFuNoDRh6yB
fXAiGfxL/YW8BJPDYPEh7xlrqYJrgHxzW0X6Rij8Y5wwP40PDgqGhm2EMgTmxGBC
aXSoj+esy2CXQ1cWIeyNovUvvAUApF9OIUmJXp5WSQvGRLvq9iE6Vv9/9USl3Ytr
GvMDwee9jcF+gA5gYzyiw7WrMlWSvpR3Q6Lr9VrIClNt9omyR1b6EhiZaXBFE/1D
+d/YCpbFiPKO6N4v5KpIQdDniV0C+CbSBG1HRPnJ5ZwHTb3dZq+U3WQ+RqEqPsrX
PePIc+e3M0mh9e4CZctRpYzEi2psFHIPrAa5d1kvKhViF59NzfbOHhzMHv2fzwY2
US3/4NPstbbgFB354oSm6EiniRPHZLHBD/kOzgSVADDNUDBXAZaxKvJNJTqKRHAm
01YIdB1bJPj44laHAqFiphhgngUX12IIFvwGCzlZQM09aptSla26mlUReMVjl9pN
+rSO8uBEijHCIl8FLmaeF04uEuoZ90BkApp7yLHWuopq0X/5yrEwlVBI6rHAyo5k
aGkThDirFcC2heLYExT43IHrX6og+5A+p3pKQA2mBAKucO4AVM85zhWGF7aPRDEK
iP/xvbjliODv/ugfS8Z5pQjy2i8/GC2+wFOVCNBRzBxOsZcriLDfup/ySpeFgVkD
SmZt5Cl0fQcWpLz4hDMJ4H7s46XpeVKkfTL88BNQGvKg80etxP7ejDk/H8uDI01W
2imIrDmooqWfbugC1ojyUIyZIhJFgEK4bMMZuc2HLxNJaK1EWGLloMniwlquFc1d
96Pfrr24o/Hzbo/saD10p9ZvBI/9h7EC6hgnDVXLjOZhdnwnd+9KA+KlRfaG2nax
Exr3dnFOggDKEZqDsXA33Sv5jI4IzmnSfmgIFBJkWtcBWiYNhn3hOTVbWqCE9SXH
iZ2cTGKSjt/BMdrAxouUD/paGVStKoOWjDDX1ZzN9i1ReKaiUkcYX2v94xvbI1QE
cttqP1I85MajtGNYGwRfG1nNaZr/vncTXN2/NmTCK90CJ1VTKjneCycDOP0d66OG
zcxff32CYyvRxIGzJHC1ty7hlf/tDHJvaYQE8Msy+yqzLxVOh14qdAql4vm3rSwF
YdgHdMFLb7Q0StDajeCpfWTw+uQ1EqbDvogXrR6cxSatArbUOq3D4xDxJd92T4pU
2XQh0xKskKg5MaW5LVYDwJkG69qqA3xpR+/53jsfjYA3/sBLZy2naY1NinwgZR+t
J6N6DGwdkaNJI13mVB+HHxHMgg8o/RiFP3tNHjVdtTPDgq89lwKBNW30mGpELx+D
jXChzQPOB946TuKOdlwxI+M15hEKVdbZKe8zomJca4W4KWeQUrGME5KU4jX7h0GA
jpxL4IbGz61plwVW2p1a3cRlPy7MHWFbH6910TxcCrB0Cl9bm4Up/pHN8AhFGhS4
vfcAxROy2HXMxQ1wBaeYtf9ihXVsFHSm9Cdad4O6W667r/3MWnMuBOrQvdci3ixV
NBUw9ewFV1UOniRSiO0KfXPPGBTyrbXtWv/Uv35c29/LaGe85cGfBpPNkZanIQLl
zLRoESeJynjdIOn/1A/pKyaLqMtu2rD4c0H421wayI+Cjeuzf99q3apxshu1EPa8
6vSvu3mI3DDApMpV5wHSYPYwp6/gPhEqRN4qK/oXHXbK7O+TIaZJ4rHS8OrVjWeM
hVy9vT+P5bBgOAm9oYgQ3ajF9HF12afOjUPv8G4v+ZbmcgB+pOVljKMLnUdutrJM
NdOack5iIe0eDQXU1byXSS2b0sdpiRXjJTy9nnU96KBsoDf5x1xf642NVQniJZgd
axjteyeQpVPn8wZi+l+p91oF5wm2cNixi/asJwYQmnDt2JW67xfuyZFOGye5eO3P
+W7TYWCloM9IiJCLmtxqZVjaT/HBEXr4FkFck3W6p5/KTqK5Dad3Qk3yaDEFNndo
/B+NZeOWF4C43/zFXBhCoeWsahsGDrMu/NNkpSpXTvhu702l7miJSECJ3p7AvCVZ
83Pgs7PWsqC3i9/DAt/5mPGo5A0nbzSZrbCK0CrVB07QUZV0V7QKAK8g+ktPGttd
yxvRa/GoJa1fXcPG8+UDUK/mXoHeyfWtcwKxVaWPjNRmWvkysdRq5kHJOiYYCf20
zJfrh+4seIf3iPWhPaRDtr3o8JgEaZGHOks5o2ubnzH78wV1XPc7iwaoS9nwyl1Z
RQTxxf5ryyQwjeq2KHIFng01tvAC8kFkRBA0Wlx3P8TKTafKP+iPTChIocnFX0Va
wHmvW3jaC/9pVkk+EN5QprqtCxRbVb4ZxZMYoqlR8NPVnKwO2EzCnw7g2YzdmY3Q
0jWUfVzC15u4aDKhDHkQORPr1ri/JrZrSV0oRG9HD3ZmiYZdtNFiOtibocP7gmdE
iLeXD35vJypPOcw+rhlR1U/6zm/cKG0ols3dNmIqOB10RyYFNLnU1/luyB4Dfykg
PtuyTKf49qG+Lv4qhjifBTd4crQ5kpZuF73+dek22S993APv/gpgKxeY/r50fUHW
bZVfsCQlej9YigW4+tY8/mEdmveeazPtQqSrdyU4A27Mg/QD2pP1euvdrZ2VPXGG
5DO9Uk+8leEb0EzL1O6VMENPgNGeQNCuGabi/u2gFg63B4Ywgu54nGZThSorEKA9
oRpzzQjoKSzQL+q8q58pN8u8LEIta86f3kpa1BLEVcZeOigroPfGhdH69iGBLR88
ShpFgDbbEKt8rikVTq9xdsMKWB9UF5X/v/nZdHNpuWEWC+YuZnjWmDwjeW5p4WzX
/VrhCfonoiTxZKK1akKG2oAmHmzRkegqTn82RbE7E0a6QLQBe2aJ2chisE7t6Q6E
WdXI/5CiLafJP3YTmvkuDnkdGAJYw7zTYETWl45ygcQMo8reAeYFDo2wOxdNEq/T
xQz3o0uSKrjfTyDCsHM48c9Ea8VfS6EKqhuqoQl1LN4I5ZhGaDvU39ZjiwsiAA/d
t/PGa1Y5OEDY7ijnH3g24lBrHThRXyVeSjYeT5zstfACsG8Qpkzl0sQb5kt37pun
S+I2CRqTg4hPHT7s9eprczbaBvs5iQ/tboaYqWtC8BhqEBjwiG1xL7de+0SX/aLS
+syBcNua/BAkdYhSa46Ba8CuhvsN7azfaHaJLxzTXxsPohiXcrcBifXiFFULPizz
ZBSSQIX59fIoeTSXz46vWuAxJWdmGIFn5hy8fEvpEvfibcc1/7WkoQq7jaxb2rc/
KAUAuDwnq30a/M4dHZijKE3AAN7lhQCcCatRtV/YqBnh9XKrSXLQd0iUfGYG2AHn
BtECfPfraB88RiQYbq+EEVbHJX60uHY3QmmGeM0sX2g9Sv7lbLgkIkJYBbaE0ECr
zCa+wE0t6PAwB1O1FBNzR96Y7sWnpLk0+ToeD1SkoTCnFKc0ySKex6MPu10wzCBj
sU8iummMHO/l+gXlaRjSBTdLgc+reg4ju1nFUl9hj0C/7VX8Gk8YcbgrNGCn0ght
KEGf+sLf3cu9yefKzYrP0n8u16kHNfCv76O0bmJK1UjU2Sg/Lqlbrgjgnwo/C77w
mH+W9KaO6Sv9xBbt8rWkwMeGyHK2oGPV1TbkhTlOl14+UTHAT/6PurlgrIpiRYQ2
3boGoQbqzXdV1/nIVkAlmIOlFfoOw6bs/0yloedkjIXANsI5bRL3NWaQv5OGFGZ+
hjauDq2NvQPfGs6sDGTMzJ17aSKOfrqJYyoK7FdAZDjHtQ6jxPwWa/P1BrzwZgxN
N1yF5ToiLRdbLMM2aIJ07Es0M/BtyM9eJn/I2p3VITRQ+VN9XR5DJv1ArFI2l+Mo
01YeLQRNg8yjWfnhohwiX581L8NPcRUWmfzcKdXOMoTZmu4GeB0O4THrQX1hAy01
o4SBgbc+T3zKB2UMt5eWxtjQ+Z6JKriEZuGAJ19U5rZ5neLYYH9GvJ9sqQEW6BE1
10A/P3V7Je4e+0OxBFmP3UHEOFzq7eisBMNLxmmTEAbLbisVmLrZJisrC79EBsHY
9tRMtR24pB5m7Hc80OL4eD/EEPH9pIOiT6phTpTfAWFqF83yfMeZ0BX/xOpBnvYh
JO1xzM60q40kX3eU5VbREaGbw5OnSYZdRmjeg5u/JfXGN/gxPn97ild4nWMbBNgU
HzOEy3UisXnV/961LZisuYBrZk3+zrmHpdZBPxXsrJwsQ4Wj+vDP9RImAke1YWc3
u+Wv4Jqh3yGby+KSzQzD2AeFVSMuM5twGxo9yKvRTWVMP7Qn6Wbsnsv3RB5AZNOF
uEpauIJrBTyxG0IoXW11xw0ShXh4X2asvtCiZw0Gzf7Bsoq8uI2IKANyZPLfvPPk
ANYp1cb+Tu0fgah3Y4Ak18b4YfhTQl4FAmruwUr9FkUSOl4/Ebbgnk73qSW7kyZA
KTLETWwVvgj/lwVq6v0xOxZOJVda3ozzljmDY9rLY1Xl3OA5s2LD/EBZHpAHZDlo
6CX6sXLr+NWl4/kmEmskFParbOjna4RzwSL1zSsFJUrANcVsV+FFim4uRnB+jgsO
TY/MUw3qNcN6/hkINNazUnE80M5y/J4+YxkkS+tPRv6xfOCabvvTdE326XGybHkd
IPfiDeBgq+lRWSucKtEPq5oPimh3wPY1u6vhlvm7ekn06OHlyBKQPjSwG6tPuNKu
Ahjr4KkYepAscoXChgakGGx1SG/EaBQnzPzQL1u5Qb3mgSvb9klAytIL1qyutGi4
n2P3vSPqKbVPhxuyyDInh8Z7vGoBaYPMTNqH9TvXf3O+OnP5RQMPLnDH4Jj/YBxZ
c3Q11lsESThnblAaODVPIOO0ENMMfywKijdBv3PESEMYtFnGTsm2ovIfVwejcScF
aOQvcQcG9clb0hUSvrscsjn7vQdpaHGRmRC2xrN0mQCn93rtb8/cw0gNJEDWnXn3
mKKgQ68R96VdKyOn5CJLrmBcJXzE+HCsA9LR6AkQcl9pMsPz9JLdiapGRfLAFDaN
SiJaPA9ECmsCmlRoiQY13Jx6zZAluA8MPKKa/DrN57MjO5wleksAcbreNdUnig9k
ZeyGfpQQlJrHs6jvrNfCMc+CXUSe9IEeUcB9UxjeSMPCyvMxrw2M7Kd2J3vH8Qfs
YiVVjYjw67RNWLc/ZXzXWoj2I/tClu2+vUIlQdkpi7PJi88iIyclX4zaEfJSfeSn
8j/c22eDLLtk/l78YTRKxrlsmH+C/JW0lMY1QZXbscxGuV4p9URmjGaroGuRk0wZ
Mf9DxJ3gonFpDudI7XIxizDUnUX9xTnETcPJltpKDjAKAMCwg4USIHSZ908+tuWd
voX8t/Ea80PH1HB4PXrNC+zigVmvdXT6rm3OuSZevQB+AnOzbFne3761OKc30UX2
JKP3CHSg/gb3RXQcXPw1CNDSqgb+QQ8cRccm3cf7qowrL0uygvb4vnI716XmNp/7
DQm7jhNeRGKG2gBrG9i8+JkqSc/mS/Sc1QkiVr0cDoRgKno7Sp5+ouuTroYKW9ud
3T+5ElOTQEai0SISfCe4QKoLzVtCMK+vK5VZAbqreYjy/GhOAPIFrs+s7DmKBlKb
ZHsSr1p08j55zzbET+jWGLXAZvQnnMd8N9F8S4jAIGLfd12NF8KrgLo3xsY/dSuS
bIb4Hu9hhSei6Fxf/831M4XQxlntVQWhkqUtqN/uFktcPpMGifHVV4CrszWtbXYs
/0Y0Pc/uTOQmEemHicaEKMD4uaSkp21nMxlbJgCRDTQFKSwnLLdu1eEP5UXPNbbf
walQFohxa/ZPEgNxp94PVTIUCQV2Di4Xc88AhsjXB00nTorPEy1ait1hWFTJkZqU
yOrw2PjfEI75WMkJO/l5XoRb/n0Tn88q7TjOICOeXD0NCBBgqA/PQ95/G83xpvq2
F35GYralnYTyCtEplipcIjWuW4VtlrqORwdlVCZL/tHEq1ZpvpFNC1IYnGj+QZs3
+3ssyv8FTgtFm0RolWt4wr8lDtf1MzHaOPsx3PcYFqH6PykGmHYVmlwGnKSg7mTO
oooEoYOQ7YsikzLXr8d+H3LKWkfAzpSxMCQgG5oDO372NeUr9iilPKgQSDJlI8dQ
Ht6mGGLwWUBQuLmTOZEsRvvBT2fqXLzjMMJN/OHFFzvj1s4atn35pRhB+RQkCtnF
gf78Dg2ezrjY5HFkBmOlIqbFV27SRPgtNMhRdSe2Qs7WbhGoCWxGMaqClyrxFMOj
LSnaOrcLfOR45alRcOqk2PC56UbuA+i5lyBsccmrYmebrdjixJlrwXXX8bOJyEEw
Ox569mB1cYweKlfd2SJ6YtFxVKjvHjCfZM4UYrIHRaDoU2zlsLwmaYNWluQ753wm
m3lod0qeunzYGmll4yJwCjzIaeIARZ1Kb0/f3a02bbOfowXb/kBiK0xDY3E1Q5js
xVQUZUcvJex9isxEo9pHO6uFpHyxJWvJCF/7YBaZoVvcoLVILWSZDLH25onDtXpo
J3Bj+GH1vZyWOU6ZpFzNT7pB2zsvFFNwv9+d+XoWt+2qAYN7m2g60QnQJXzWvesC
FHD8VqIU8fKfgDPHdWCdXYsaUsdqmUHAyYjOIqNZ3ZaNaQzGUWfeddNMKVTQlJ3u
nhUz8/a0enEF2nt1oAmLQyX2fMATMO81Ib7UJWQJQq9DJwuVY0aEUglW2TW+1O+S
w3VBFeV8svQX78VMawIBnU4ejvpQ0weAgji9c0mrnloyyYpJZ6+RUyWuRh/iFDsS
GV82WrDybVYz1qN7LZYS1QuOXSagPOXjIPUPs/jUKJTFlP7kpfv7GRbOaPbScjKo
QZEjrM1GBtGwl6iXLNa5dNevVMMhXblCFBQl0zeIfOTnrWJZEJlcSyezpER2eO1b
C7ir2TaZz1IchH1jAlyMUfGP3dV9zU9pbaKSxmOTA5PFO7gh0NSX/SvePDsTdTGa
HoKh3HDQ0raq5UcDw8lKrQUCm/EveGQ9TBIWbzrzM1WI6te6JXe8yw1TJXagz/lE
vK8XNwzOv4F4uH8EFU0H9IEf7XAERI8mgsEKW1km9tQSmXenPvMy7eYWbjzpjgHn
bfSaN2DVJ1HWLr4yi1VvhYk8LCm4yZFdGCoLzkxOg6CrmZoRzOHJoWvQCef9087h
NvgKJI8WGlFSalL40tbOPjum3V/8ywjzuq9U5KYvSap++rzzq1EZfrdDeViAXKeC
rPnm2K/MjpN0htfyv/dfquWCNRKyw8MCu1lUpVgfHXm1CZg1BeObwb8aBzdXgxQI
lBHW43R4Q4+BXVgcAcdOqcj07Rc0bXmjmu1HBo7DTT78ewXMKmLh+mZaJSWuEQvU
OJoNq+vSSfIuacwbd7UM0WtJmS4KS8RNPfwJ5acgq248CHJUTdKRgZ5/iFTdLcV9
ey1C/vkrE7puJSYNkVnWFqvyb0KlY8CzN+3biP190ZFTEPIX6llNo6UiumZBy43R
sW3wpbVcGY1/Hctm+uIC3ob/InCynxu0nCgZVeKAIN7sXrejVL6dRF4aLpp+2B9o
5CbTnfbJhQ7OsoyfIuiAfjRZ4s4MoX8y6YJZ6q6ss3DQqj/cYljlPRCT7khp0lRe
u/XsrGhPXlQHhvy0R4RSt4NjFOUCtUdiBqwhGOZgrRmNMoVmNMBnuEHmUsSeZzZU
r8wvfwEuleWXt9nFE4oA8SUlXmhGuKdcuCaU7eRPyHcm+TMFSHTP4eGX59ArSkEs
hPi8rFZzjcdVdMMOsaTgc0GPl1352oyO+Jj0aLEo2iBTPZcHkmEvvEX+FgnOcxX+
TYQIIBISqlxPlEpiOtVU4ixkdTT9L7d36GuZ3hbESkdwYdf/YtD1g4t0lLnUKjE6
k9cpASnTWJXqtqBqRkakK0BT1nrjtzQzpZI8AoV3b7uR59Lf4ykpyQKZs1YUIeoG
xwipTwBplkqrI1mAtafhG6rLAzTwDPMqHgz5e4nlUuLCotxRKt24hZ0kv6TU2++6
O7tqZb7nJdtZMrWhD35ooLaCACexdUEK69Y+DtJry59mvZbfCZ/Gu8D7YoOohH5D
0/4VoZgh+rHUS2VzLa6ls6DkqN+BXh33sABOuizBhdNE+7KMbDycuukeiYI27ZwP
d/vYeTN1t8tYwvLUUyGddUgg3WSO2Wzanlof2L0pF5xavPmmOLBwit/uW6EWVX1S
kHpWdkEbb1+O+qoAqkj9BejqR+wcQoARLwuZjBxNdq0Q5ACQglpC+V3coRSRQOCY
oVUDU/cUz6q4tiZqB8kPUgHKG1ZaeUPLJf/lplOus6lw1aaU9rAdnzp6+OUJ5kIC
GyYEIm1mad9d8wqMIfJUsRKa5rohTqW76+QU92B+a8MOtyWe20wBaLDRQF2FzTNE
9SZxlCWWISsNF6AiIzPFj4QlDDcT50h61I5mce3OBLlCwBF1MLqmE84FhsBHaPXk
FXYRscqslkKEweWee2Yekz4Qxd1ZUgl36+xCy/zf/x9W4YAZ9KnxCvT/1S5QVc36
jr6DUIJh++1gwarBOJGlGvXTbhTSuXtwzccl1RXr+govbmC96xa94MKCtfUpkCh1
V3G8NYDEQ96nFxHWUAI7I5h0duvfbZxbBPY5cbGvdYlHmX7to61yruIqJyzkBlCU
Xg3GHF58zHSnWd33QvYXtrWfieq1/Wee8++21jp7qR+fLXNA3siZjCwhNL2XIpZc
IHw/8KvwaXxpWRKUsTXNAEgimgiTfPil1pM6De54TaAJ8X+FEXYLp9aF1oV06xe8
0t0YcAk6/sjgQrSqr1uK8SFiS4svt0gLLAs6AHwnMD2Yp0A4dQNOQbEhvJJLsMGI
9CvU21fWtXBfVLtZ+v7AkQx8i6Z5K4rQnbOlWPBY7YkmCMk1sn5MInFaovgdDMvq
JNZfgtTURYmvHUlmMQR+6alYKFlmOHAxpoIHc3pQlAoO6OFzJGY5QN3KJUahSZHM
m2hZaeb/0w3/EEL/uHbtHbPN/8w5Y/jkL64Y9iQ2bOpF4bPBpYsWkmbW/eXm57QP
1tZN6g1Mgnqu910dv8SgpkKuupUg9WjLr9r+sF5teh2HzEOTaIQFehvp2Lb219xR
g95k5Pt9MJtfdosrcT6bWVGa/dNzMWuy0fHO+Xw9VP9NZCXOqPTASxwsA8DNbnGE
6s7muwPrc3TS2ynF2I0JZNXNVzwYAGKVHTvoAqutMKPx7XrBpGAiS+6Bb73wqRNV
TR5cpOpc+7pcK0ZaWBMiinrfnaeeNXo/cDUOO1hlak6bDLlkIXuQqYjJ+JSoJIwo
k4TCMtqdOAMBwpjVmiJ87/5mcp+8OJ003egkxtQh3bU0TnrrI9T/eF1Bk9Ejq0p4
l7iAkXn0LW1Ukv4lazjQ5xRXWPiavtcsJhtDP+t1dBzG1sx9L+T7Dk5BLmWAG67o
5gIoivoe2IYROI5Hsy3f1qVW/mCwMGd+Zozs7u33/mjCQW4UzqaH2Qf06ced8Ve6
HU7XSTAuZQgBVmabSy5PoyRvEV4YAghih8FrQUXZ17E5taqkyn8jaJW6IToPnp8x
xvMqO7iLrQazu2yU/4+l9HjQDhy9b+ojifb2jBqEZNwdD0mOrtt8UYqXkOqI3Lt9
KZ1/bAH+RpsVfpeRRDy1MDaJrvWxB6RP6TQPbLx5LN41Cvh2BmMbBJ1AIFsCgv5N
ZtN5yTvF1boNp3vnv0M9EPFy0mHItXkSOJ5i3TuN2eBzIMuhfcguaxRLFf2Y6lY0
6OoOFgNPB03+CeihcI7sjK1vRHnTr5ikixWwu/fZd+tTYVuVoO/jsgVsZOS+A/zw
rgW8U1mYD/Kx4NSRsEJ0TPT9TL7jd9at5tdqY2MUy4DZbJBr6MntyN7PItm9TLUr
5g5RJQMf46snyHuo2vwaKL1G+JpUTC2blEKnNVmX5UL9GDwXQZOe2VH0+AY0UbCV
nc6xCDBZiLrgFQqxLMz2a3r8oNiIVXwK+QA0tOx7JyH4cr0swGl8jhcOo/jLLRcK
unOJGFYsMCKc8tdud2ShkqSozwCexbUggYCRFmL51aDHe5P0n/quaA8ttkBPdH0t
9llYLGygmPbOQgEHRpvQRTB84cBQHMPOy1Ps74R+Xn2q0Xt1MqKc6B9S/SPwpP8C
+9+DXf2LDVjSPu6ThLJlvKVXAZxRETLvqSoLRXfFysgjarfFRfEgVONNpIJNrj/B
9u9g0xtsb/UztS+79BmAh8qdP7OiyAAI4q4Bu7m4VqY5hY2RXIeWO1LBLhWeip/u
X1LicP082af3TRAHRhP49gusaX+Gux2I9wgpNAYNEMYdtmyAskz5Ixe4HznXDL6U
DeRF59Arec8DhBm8kf4HG9SFV5d26v46i2aTZWI6ajlS+2Q9heoZ5oBKVITw+wjO
YD0xmFhjo5srdcb/uNgGyw8KTpmU9BsVE0SduZWT4Ct3AxzsmKb7BtghqHCmWTnw
QSPyg0UXEMqAAbu692xgCSc1ixY+195/6gdl9Yc86aeIAi9uJmnQe+nn6WVeSHSo
/KGCf1kXDdc/Vhw8YQBr8B1622Z0gGO1jdRkw8zGFtjmYbvJJsio84j/tIDMk2XK
PDDpdTn0Z7ERz7pMClXlImi4IVRLvSmnWCmv93+mDzO0ldBylf0S7UE6WfI5F+x7
3BwD28xaZklUKOCb9rLECy7d4NEl3ONP/fnLK2uoqrsRnxf/P46XxEyaumO5qt/l
PRcjwwH+OHDjyIx8FEOHMDN9f1zgl4IpbdqNoNl+CAZPWruqj8yoC9rnJEqzFW+d
PpW6q8aWqhjEI8XgT7raJw9fFwKVtID0whCAU1te4Oyv9FNs1F5Rgz8MvQGFUP7T
dw7Gmc0hojOhC33KO7UsvwX1m2X4dX0jggyOLWcEsDau5/LmAbFwXZRHmHvA0mGF
HK0dbh3ra9hPgwTNLZSwBH0QF+uAZvyQbtXQdPR2lQ9xxzBW+NyN+f1gvgQ5reO5
fK5GN4OXM1GCK6dpdkI42ShGpCajchlzUFgY5MdSATlx4WrkDBN1c/0USOq+7ccW
CGQsqXMd9eUu6IZX5ttUkqAhbcuqzz3sI1PC0leRMJwYRrnJkpeY5+O2D/DR181S
11RfTcmAJuFqwYtsJv0UYSqjbmkcr+NwG9VIQXlJun5plBVFkLNrMFFVBS6ws5/j
3QALGfoBovGMgnsJmTeVmONsvThKx1TDeRUkzdyjWZQr5+kHpWcxxQay7FEI5Cqz
YivLHanIH0ZK/l84P9sBKa/Revewld999lVSCr5GvUkyRV65/MtWi2YgXbPh4Qa3
c0j/A4PoAmEwq7QWY7gUfGiLSeKNQbg+mwvIQf2YAZh8Zl+7JjM3ynlApicgBfdi
UiTHpig05Z7x02mnGqyxjQWCMWRqOJsuF2o1iMZvYqHi8bKwjXHuju9g12HdisOt
EFJvFEcWcjFYu8sAp/WiJKwVU9tFzLzoBbS6IL+SBhHAzafETbO1g2SM7Md6H12a
kkcapcxikORJRjNIhvpJiEwaDoejfhzDnxxnoe8aKaKMF3PTokI3+3il+3XB165s
AHHf/mR17kotzjXPlSk9yUaiCyNHC2k0u7i0h4XNKV4reahxasVTtWHV8y/tfh6i
KKN3g2XAAOtSIGLjMRzhVveZWAqNCLKyb4Fi0bM9NaoNVgoKevY3RjaWbes03Lu6
FOyXgHAhBMz4OsWAUoqOXTPQsBT8ow73mrMH8xNm9fQtSxVbvoCm3/sjXovum4H+
NNL25/yt5B2zqzKuHm6Q90M7TY5uPIil0VitgOtJwyv8dGHk2dp3YybZRSLjVjC8
LFtOxh9SnT4In7tNPAbI8ABZ91HI19EAoc5beXyqfr866B0APeL6m+fubzj5JWt6
/NeUAPGi+W0eNErSArMmYbc+Kh4vjtw8wJG82zFD/Qb4fi0r72UaZkOcwflR7c/H
i25vxne7j3D9rZ/FL/6fUkXpcrSTFDBd/PYjWq0+RP9ax7iS3dxP0cwXP9zEl8+B
By8Red354LihW845Z+POwMWk2CrvaoofUaCbQBhGJBvzM6CDTc8YkoGmynxDQGN0
SO9K3l7y5htsCmCOJDyx82JW3aR0DQ/fBWG8rJCaeCei3ITiuKwUKGNwFX7w+qew
7UOzPC6cJymJ7x99pfjghnGQpyy8jOuv3/Hpx/chmz/wbcKzzejriKVY486WzKT6
UOGSMv2VfFl/XnKnsf34xNDA2MheAvqTWHd9IupX0oeqIwsHjcwAEDf7rJCE4ekC
qw6ce5QGrGtbPHOSpKvOQzXBkm5m29Nu0rs9YCBmJOQ47hjWJgvo2ctYdSqBzyhl
yaSabxnsupBNpx0hDiZGqO1rpG2AQ3RZml12YN1U7psNJxhPqyP2X4BaOA6qH0YV
dEu6SjkSl3H8Dd4OvkExWIhy9QIfokoK9yH65bC+OrZpYNXXv6KGAr7jwk8x4HcD
n0WtE5/q+hGCWXAx4BS4xYnRwO/jfSr9l/9mYM1DmtCBkjjhHZQj9OEgow5+ZCla
8MCRpMOr33AbV2jdm3WfaKil4/XpID8TtCr2/28qg9kQX9m73DiyPfP2QnoRV3Wk
fLn+z2aNn9l0cY2im5m138ChjjA7i75DUVwJM7HZ3tRy0TR/Uy5PC5AejgaBl4CI
gaxt62Tz6BFXk8IY2xAFOmvnvk+9kiuxuqPrONXXOEcM+gbZ0tJtwQkmmNIr9Ade
4ivZPsEF/b5dm39HEOGqUH5+2xmZetYyEbVjUFtCAGRqbOSb+V16Qc3P95+wEYrj
g0UhckEixkFTXGilkMW31yNRHYRSJrVP5NTIaYsDVWdfKTO59LvOwGZQ3dkTvIcU
zorN/ijuhcByqESQCktkz26fuJaDibuaDJ/BsAHKVUeHz7DE7xs0tR7+oR9KCNgO
udBpLcEWV+t2Grm8Ir+43eWjCnHXIdYnRoClD0dPf7+r5Qh/kopnTKFovYbLq+Q/
o9mZss7Cb8YhDPwe52RVSyUqqrCnETnhb2K4ncyOT+6mBV6zPnUQ2LBJ8rkh3a4D
jPcMGcx3WTF6mLz53iDxU/QbjUZ0ifUg7cILUQvQTpmRL8cjQ5WtUFpYFtEV0cVc
wnaP9fSg+0UQMyt9GhcMQkKo7FAZsiDxZhshvkr5HUWama1ILvbeXG2y4NulRFPA
6iFyhkVcygJ48dJjRpgIeFB0qk5tqInqP6DdAFJrEQYU6bJUY94neklVuiN3TpPu
ByyjGffedgnS3FhJH+Zo6svuVRTZ1lJoEZ98YLdoxFKJjoEK2JXsb8+Fap3YzQth
YEwZcXRrmNnGYzALI3nm/2exHFb8uRME9eAB7V5nS1WAFnaMY27dbyt4igWhVZAT
PGgSRIALu2IB5/URUmTCbpagfBV3SZ5pDVdqsIz66QfVGlPhChMqECUFXchBvftg
rkzJUY+AL0AsPxaRhOdw5SxIOVyT0wZ+TcYJjBfSbaxFtK9RwVhYUJKxRkdqJDJY
hIFjhvOhjyB3PKfkB1rbQO1a3QQrPX0jrAPUA8ygHDXnIUsho10tKqeUjTaw09ir
cYbxWfuOBbwzO5hSbq7je/ASQVgy72Q+jfVo+aWEUi1zBWQI/eQqTNmA/pKiFTXb
gKFCRG2fOdmdCxMYm57uDqjhjgtUJw6TQ5G4kgkbUHqsBy0IwpTUeaRLYSvELSx+
fYyb3bDm1eTQvYylFWvTWRxz7NF6DPOF66FdSpsDcBNktYiboiQ3wG7jeFn6ZobB
si+cU9HdrWFQ+l81d21KaC9wdl3ZEtVHC38VLnfJXAdFgeAsP4Lvv1Sg6aazXBs1
4x2t4Ms/m1uayVaVn/NBI27st8YUXfQgavjUpxFa4SUaeBaPsEhmvg2QDiW0KgmN
g5dYMOFXGR4u7tGZlddpIIuuXltRuGqQZSedGWZNwHmQ6nf+sSr7MeJl7hEG0e3Q
0e821qiiFrlbHlXf0j83ZtSTrQ++P2QMCsr6tsu1JqG+cjKqiHN9JPlBVCjhQeFU
gsua9riK50PjcnT5Taw/Yh2GzwZBLhiNMcUXTWSWQllFJ9NHRvIHm0S1XY3tQhNR
4AQFn1NAcct/upCeaCreIhckOKam8pmm/Ks/ghg++bfN6yn1o+1zUoJQS+ky0T6k
qHeH1rrrushrYJfKDN7uvhbrWFSJXD228c0wO3pA9lRDk/oQ6Vr8ZKou5J+0mg+K
0cuYm9mqqZ1JT70OWTI2GItrVV2GpHnwzV4arpi9baJPdurZF01kWxVSKRwWUI2/
wJNieJXNzy+K7PG3YZc5eOVJvCECk8keyne9mjakl06X+h/r3IntAwQjXfftqi2i
PizgSWNqK3Wg7OG212/yaCvbqnydRK2M0FC/P6ojM7py2re1YmB+CvXe1kszfJpS
lv7M0DtUiv+1iKwRlv/2x/QCXTwxvOrOUo3v45GbSeX2EoIbX/bimY5siV94aCMt
2dJR2VIucmmvRM5i+/0vJH+l9lbkv/5lyxl/lUNThrpyHNzqOyBS/ByfDe0zOC3S
xjGH66qyVQN3jtO68O/gJVpH9bjthNt33ernliT4+85eL3FNo2QqBp63mv0E5T7f
LdCdMlagHZ9FD7j6v92xkgrWjt5uldy6r0U3qAkY9HznhHyFqoiyXi3i4Bba8n8A
ve5U36WF6JI33yANAQ0jVL5tomyi5ngPUqT4MgTidB1ZWB+rvdWDTQ5uGN54/84n
/oyo2D+BCt7vBi9nNPBNIr5KzYdhAztVv2c72Wu7Ld/u+ASvBimskVyGenZ5tdW/
mylLuheGsKX6x8ZhYosxc85Fz4EAphtjpdQXJXy+8PgKN/oQYd35xDe0nVK8H+YD
U1kbxjxxGRVVfVXwIiCqdVhlo1p8uawZaGzppoK0Lk1Wr2xdxXwFrVjF6YHs3NTs
NMG/h9jvuwlDq7hkEqMG96FkwVTltMNOz3kQnqM3Rbeks6vvyAWkgHQ9PV5LH008
zJurNzh2lKaFpLa4/6Mecz0WC5S0Y2M+3sji8xk9C52nLRaPqaTnK1lR89Xgnehp
uXo3LUAqROIiZd49sra7OxA1148vc1SdtO9vPeKy1/I0lA98Phk3Ea7Dhike/bty
SUJ4lY4dgDMrN4GvCoAEX2gOsy5DFfzOrz9XOc6EHR80r8hH4j+OexXREO2+7H1m
W87iUH/sWkmZwrtWu5I+MKQO/1ZxFlfiNPrVq5BiQi8DJZHGYsxL2o7VVHfKOrOp
5Gvg4ieWJZcmbeDYEzLaAHQPVqIBGAgJSBpidC+HplbYl3nW8/VTlViOgL/vryEx
dIGrGAUN0f7aRp63czuGfLZOzQ/xzHhx2ChOrEorlrKPS5LKK2X61yf8NAcJnL4P
yggiOLD6D9fUUWeqB8Vrx/rqAyHvUXOVsTBqp/NYR4kmdRszgDtDGr50byXY2AqF
VAzXyBXmj9VQz4REYy5+rw9cKwUxX8pbRikQhgsWhNOEz24d2p3V9ZusCaymb2B3
hUf23SgTvAcXvOiTVQya3cv2MgW3vJGOn8GED9lazhgU/o7DjCIfQWH7e+4ZXFPg
do62MnvogtB1uWNmNOcHdsD67jd1hfhhMMTj68/nnIyjy/0yTIIOe7m94VkGjAQs
25vc0cO+4Y47u31/pjicIRHkjWuUA5pQQqmMFhJxuNPpakHlXxgzdLqcgiJh3Pc9
vSWLk/35m/P5IJSnGr+ANkMXBTIdx9dd/CDEeS6109VV9EV5pRKOEKkEOoYTiJ86
2IJZky59HbwlXrGO1opXpucqAIBgbiJcA0tUSje5cXKwUnLIIM4KwaV2Lu/f/tDa
diGo5b0VOc//Mqf1cEdMw1WKDR2p7sA4+ffJB+VpOyZ1e1bHLn16V5Cks7u54BIk
amUFO/lcQFS/SgVqCBjyZJV1Sm7MQXFa3lLvXa6qGDDiwQo+aNPZpaRj9h7QfiCh
n2wgIqTsDFxJ6iykMF4dScer39LjSZVD7z/vTfMxbVizrpk+bvhMofOxZ8amTSgj
OifGAmGmYAx0JBThgNhNt5Lmy2DdbF2VmkbAj6Nc97SVBnMfFFSYqBOIobr2L1ot
r00od1dFQ53uQpEkhvMz0U2/81X8YhfyyQYRBpBKnNzRsCHEpWVzlDCpJ5oQR28a
tSVvS5rQJpoq/QfoM4vhvMGt8eFIFidAAJZdUbfJxnfP7r0NblZvxEIHBsX6msuG
5oGnqxR57sh4ogtt7nqZhNaRHAbEojFU5Mbwy60IbFzzID3v76j//jkMxqq16eLe
5+dnc+TjNFTv+kgsfBwjS6skstolJ4ahGy8jSfxKkngVpKxk8BsHPIwDrwZmpSjn
/9kZC2mFnOtHSXxB2hcMOrLFQihbL/c9C+MhEG8dJHaEBuPFhDNtv1VWYiKMLE0h
cDdpr+Zt2XAn8dO6gQFHfF07Biu4hofcLzNiPmqKfGQe+0gk9udSrNKsmwZjHQ+n
ZYGXBVIanQFowQBtFEUjiBBDMgv/5xM2J4O17kSICm6ctSUT85xAipoOLCGlyepi
e3IP/nQwOmXcoGKcZ6Xb5m01wApAEsBlbjsnARAzY55GivxDFC8QHRLn4oDllwTy
24hrs2E4Lq9uYAnNVCTV/+q3e5zO8zRhTGtV17Jyz3YxItmQL4bfKV08VXJkPTHb
ELUQecxas0lwWWH+tAiyHtYqIAMUkpCGz5O1UK+fH6CpArQ3awbiZydUqQQwTwH6
LZwxuVUJxNqPwm9oTQscoMyosj6mXw2sW67WBFvScQSJ2JqfriglHZZeG3rxwll+
Fj6gA4LcEkylTKpGd1dHZPK6M4vRCvEijTEueykVkVdfSvkvUri4KMuLko6S5tcL
Ld6FKs8zUcvOGBMKyp4gazH13I07Q2nwinwQ+uNOxDQEbQYiUtmcVtzJ8lNBd4jz
4UV3CJBlyd3t1vdAMp+I69Rp0QdCvd7Z2Omft3mf3uJJEJML+bKDeUQendYngYe0
xGNCbhF8tKaNXT82b6P+74NHHtlR8lTPNaI7utYzmimITJtiNlelU6IUcORiNwpu
TrhOVjWsHL+TLTU+KM/P41v4JrEIqgDzBkwQ+iMMIVTycGI/Z2cZkvEo2ObSKFcn
LxTAzhHTij1F5JgkVqij+24Q+zpoyVVgA9l1/+VPfIP8YiWLNzOHqd2DmyYoaCtb
+GFQkod6haSDOtJdZn05ULxtTfLHf7gmqRSLAUp8ZRzl7b+7NyQne/Bdyn264+b8
FA/IrIvDQ2nTeyrELcUnZTpG8m+OGob6dhG9FcCqJxyzqUOBXuDsLh9VisdM8rT4
77MaMqjgpJespLYhGJ0W760jgLTHCuaxshBaRKYo5lLYx3d5hS+LMAgpK6e5bAbJ
LFXq6La6o1RnElAvNmJtghVCUTn9sy7uXF/8l43YQF/XDIaX7NydMDVeNcPJ9P5L
ph1bDlQnUN1OX1pbYcdOyCDkm7MWdiXmAQyTS4LS+T2DHY0wtu44f6f3L5oQPHny
0WUfcsl1LHd4Mu/4IBDhnl3DwIpKhPy0zU7q4e9Rsha10SrIW2lOu7K0PxeWjh9k
ciEGuICIWN0nEXFJAiToTIiEViYH2npHRh7rmqSwbMK20HvyMFjkVW3st3kkwh6L
hvEebJuC2vyb41+wQOFoyWdn9Z//vQXXCeK9wTkcq63e6jr/ADK9WeVNuMcsJ/jz
rrs/9xix6wvsiTWaT/nlHULGKM3gt4FqSlQF3c8R76Flgg4GMiBMogAb35wM5ilQ
7vGOs6jjsKuGoAHE4oTfCI9iT1L1E0BMGb9PMQcJL4cTF5BYKfgWFnjPknvd4Q+1
D2VLOCGiFu3zRchJCOenjTsQdq/e4VGTT/S1bKkM5iZK/eIZX1Y2dYeYnssMR9P5
JROfyIs3kanPsPcPC/Hui7VCAHLRmWbbRSTIPO17X16Bofq0Qz3mTxu/8Jt062f6
NVTegoPkSMZCya3K5hbsjkb1hEJG6P2QSAS4dVR6n3VyVHPZCvghywAR+qXcpNFa
8i03cDspPST5QCfbRNXxXJBMQLh21ZRpOoeiwM+oGvQYHSteNjtsxCkppvpY3mQh
u0Hznk8fLE/qdspbNBLr8bMfrTRC3ARfvDD0V2vq0sBOJ5sKnAVd53wcrJ1Ykmek
HOwCeDCXqx/l48LQkOGW5JgC/E5KN8XWq3fi+D3eLxERQM9MVouY3Xn1Y+ynsClH
q/5hTwIZMjhQ14oCpHpIJKjcCQnPx5C4EIJug3t4QkEYlVpd/qLFlNKyyRYVerdK
pMFHdSF96+bGrWearZoEnNZlTZGZ0EM2YdaJP8U/UqHDgbFBF5QH0dH6KmheVbkB
bvV4K8sTOlU4RhdUWr465KEsu6/MEneEAGYLiLjyQYWuHV6gx48mhQABSg8HjVRo
dsFws0Sj8fzO2W65hLeU0uJALGQ+s4O+8Mp7Ne4lW3pJaBOHwoL/wKc6D22G+2fW
wJsB38oWnxtB71u5pGm/GNFzV+FB1Shdfdrl33k1aCsRkpGB0Is6XCHVk6ItXc1a
MBdQpqen5Yi3UTrOe1cKe/m/M39eXoPn/XhsRsxXMSOeglgdtWZutHQk+tGWnWoF
XX9JQrpAoENUmFLY20oj/3kdZUI6Cb9/SZDX4E7lHdhXKS/HB6vmvCx1kUO7rlAe
SYivbTajb3Cf4O7Ssi6f52esXqXqLGhWaYe4EWgokMczUyiENIcvF0St7xN+jgG2
+duvdnEMrqKIV3k4a6i898rH2MyhzIg0b451SdhX/F312IpqTJa9tIJPhzJcUgQO
WTY/ix0mtUU1XFf34gZpmc5B7iZzW6rdNyq7ImDZQsEG7ITATWtBY0TD6HIYsauu
aar6zQUHqGE1y9Was4nvVWKLB97GwJAEwshl7cbjdAeIx+bs0nzOxxo7aVplaTBS
AOD/nMSqqPVJwcxTSmsfvgaKLsNJCyc1Rk4AimzK6iJ+LJaasUE9FwDMzbwqmkoI
Q+wtAQ1fIGUuletGOnhInQCbGcGonFZ92MOnTT6zbpAbfjc1bh5Yatkj8a99lGCS
g+8m5rawammPYseVRATlDIXiFt6tVGf3ARAnYOTqhF9w8feSAjC2ddPYavt73AZW
Ig/0OhHx91aXBnKn6HFgoznDbx1yL+XOqJ+XeHf0JLS4OfuspNMSMIU6FD5SRgGQ
PhiSy2k7PyynqUUS8vDwWT+tCl9JLTYTij34nVkEG8zR07amOf5CW3oTd2nBoA6u
clVwgyoIqv5GIXzH+ZxMLXDmCFGwVyjI9RT7dXw3jgNS4vwW1e/E2DAh7Uk3N7DG
/48N1UtQb7QGAaWfb32988QsXSlxZ/3kkT/HQ/WWjoeoWHhs+NuReufun4Jfn3LM
v7VZTs1UziuwIC8ipZFtTsn4TLsUryI45nofKvpxC3z+rSRKrLN2fkdJMsS1PA/j
zM/vF4qULUbg5SMelWHLhyXVrk6p42dmPJ7Y4RYkI0SyzziU+em80ZFKKoKzgYhJ
yLgsdJOHRCqx9YvQGk/2esnS9Yiu9KbjNGSlDZSk4/IYvaBuNoTVEKPIWAJt9l4S
Bn6jGeXSUlzaDSRa4PiC23DTutcGXfYsQ0q6VY99rHIWeuFowH8OtmH4RNJZWGrd
QFZuR0cQXEs3NF0veJgdlP9azcZCOLIYQTQ8JLkehQi9T+CU62tObxMy+dUzopxU
OYHQc3JPXB14zpdX3d/Qz1+jWzQtNJ9cU2/W319ZtLH/nfihg8ogQp4tOOL9IMHw
01QpLyZ87plwUHvRfYWl82m3UE8MHxq656llHo/PtDWWzIjz8Drph4cs9mEQJkg/
PfnsiPGlwz+XG3ME4mzaiiapB6oTMvIGx38xVpLWV0bV0ABVC5OQUas03n8bcvDf
CmBNeQWrhuf7g7p6HKbCx2S4yv67SsdfJHOfOgpYlw6j+RX4dZRW+/Y05xJL4bT7
hOsUI7C/PNFTSsMDdym4W9VUPx2sqwuKbo/p0q2ddwptdjMCWGIA/4ioA1CS1Jdq
g6AKQ8TXcf6X6xq916r3VLaYZ1/Uq0JTi5rA4dyJgCaUcT8YBq76sTrPlsq+cX7D
pp3vjJod+bvBxrKFi1oreF8sQcnLTlQuSjFPnS7M1FuRqjN12OOCfI5FS6mzWfzG
JWRLTzim9DpKj8rzYBK5wOwJ/r4GpKXubCu3MKI75fDEWGzRVkRY07ribgbp7eab
ACSF8QHva4GD75XYBrUtCzDI3jiPaYRTeSR4602jcvHQJIeo+IhCHClTJ4gCAdTf
RMLDb8t7ZBDBcQcHQXYGAYYGXVEjEsjWBN863hMuw8w6/qGgsptN7oX/Yc5Ojv/D
u0Q2Mkk+FqolTgQGGs1QNME417QGlLL7Tf7neqK3fBRkcmZzJvTXGjqofOOR/QU2
Ef3jyMpZd9Adm+kMR9T0H30Oj65ZLKSv2mY1eyBUHuaGaijOvaNCP7HjOUkM8J8L
MHpmVC5JfSj1bh3JAI5y8fRICUMfI7xxKaTYScYIUCWtGRDK2vUhywW6bf5Ty3w7
d6IWnnu4BQz7XC7l6PRYN7hlFuKm+stB9GFs0tyu8C217bnaCecca3yDAL/HqCLg
Xuz5h56R0k195nRUWWzNVwQV72GzhuPMzUo//pZxCqNEPBiX1RcPXabszqan1gud
+GQoZ2xXtmcV6yrTVtZUUVyNgrtKVQK1WMgUsMGYdkwwxsNSSSXaNfSdKdJYCR8x
3+3ncDJWq/IKwJOms3FChBriJ6Mu88aVRCTG7/cGh7lpm441tky/WtxM1AFRdXZy
V9KU8k8skSw0bBq5IqUaXy1wqX2kHq+WTj0ud8/lYKXHmizR5tHeC9zdma0e/XmZ
2k+OCbP9HTuQQMPRq1B3doZ19O78HCf1x/xTudH/Yyyf0sm3QPpZakL3yvRBfIb9
sskIGwRssNk/Z21n6g2zLGdRhhLZQ0HaJVwSQDS96qroYhOArnpJ8bsHwRk6Ed95
9kybPJtAZipwmMKPybmkCqMIJTORByILeZcu5EWgJUK1IjbbRdPCFnjMrfH4fIe7
fJy3mxcCXJZnimiGJyufHtZXTRuITbraRVTrxyODJhf5sP5+U+fTKvW+Iu+MmI2C
GjL1nCa9FrBwGkpR80KuA53LY9xB8ql8SVPmm5ayQyYUa4nfgAAWO+ifnvD6vDUf
gT6f0lk3SqwNmoMUx1YyvG19LlNh/hiMVSDh8zsopDF6uZ8l5KN2nWy4leF8dAvK
DgDrFQLv9H8Kty85VBFmpqUWOd7JkEWBkSpbwMxMUTfmQ93247HOJcyVz51l46u+
iBDqWTvuLGUwzEJUi5yP47V8/tAnbtj6ZS9Zk8OwnXUgepSSlQ2CBgUbzbe8nlIe
fjfqeb+ZmeKVU7U29s8Zqp/hhtZsg7QBLhcZRsocsI6XiIme+xIflIGtLXG0xb03
QIX4OCuRQzFIixBgdgniaF3c6HLX1XYvtngifQUycRCZj9qA1AGjh8na2vl54Rfi
WFIxrXeEq1W54Q6NeN2Y6T1FeGW3j2DNipScmOsUsOCn+7jjCYZypXTPnwONnI3p
QTyQkNd0saXXwpvb2v86LeX5bwJKY+qKkqTsebgrF+ygRarxJgbF/4z8KHFWyLlm
0Cdy0mt2zyS+vTjR3q3+iNlE+cdDm2TTeuQ2dDej+qL8Xoc5pxuhsXzw/1a/zuBd
dzKveYcTVR1/wgakBdB0UDZ4pj/zJuuXEk7+eSgQivqsIZrXAdGPhNu+/YExz29C
BCvgXeCZ+2tmPa+71QCjiQ3eVldIp/ADmAxsN4YOmLnz9YcCnpAEl9Cmzi0RKdN+
8ogu07Z4eu9zByRLf+DNE4wfgCn+wK6KtWyBTpMuaP7i984J9k5KzcK4LPDBP37f
m0sfMqhWpBi71oNwEj37o1g1Q7GEc5tCf91vzPGAY9hxmG6TM3Fzv28Tnt5Ai1e9
jXVCJIpsLYTVTOcxySi0IWHO3yszqFqlXq7otO2z0DTaju+JvmsFCQ3YIXZUyy04
9zoL6o4Fo2pYObMnVGN323GHwI8/2GDmqZ2pxVJzJ23lGGtHysm8wFqSI6w8iqkD
KPdxU76/7xkjM7qZljmUNSltr9qOhHDpq3jyNpbHbmxeAV3J5O/hzoVa79N/Q2cO
hN/5XUJIEuA8mAsvAOd+VBxplpSWjAPmG3pvV/x4Sj5nY0hBoYH7enbYWlTVEVRh
Ttk+VyG2GWcQ3zmW4BezAGHkbElTugnZZ0NNxVC5kjP2e+l0z9zJ6aCztaXQRCWc
7vCa7yyaRPvMXQsiV185jXTiXOaPpYsbBczpDO6+IUh9biwPcAC6Mxj5YCD8ah3G
97+H9j6M4oukV9yhlvdOgx1+bcH3YiUdYaAtv5qP9IQgbcCL9GVcTDdEnOC6WUHu
wWYtNW0CEe4xnXwI8ESUr1qKSxFjCoMwOnjWGlE+8enEQ273ZSTPwdy3Jw7y9KYY
PGG7gmOlCnRwdBbDSz8f38AaDasvDTp6soiiLkf34IaM81/blDRjwvEWGWLjuO34
8HyUOMgtgcZHCDgPrv+mKscQ9Oe+plWwh6ZojO52Twv7PbdufqN5ZWWVduBwezZ7
gwAAzfygQlC11nESxj4q+HfySicHWbPg/O5WdFjruqKwZwTA6LHYpTR0vRndVNu4
ZOkjAX1buNuXWf34zBxMWAaYoytP7Ic3RLJ45jipKP66LGRkwQxZdgoeecqQO3/U
CC9Hh++/hFFaRZwuvAmOLc24ZBr75azwwvWZXr9tAG3NcKnBe873l2BxmCyYA3O+
o4QylsGTAXcpGFq5SSBz4epIIhQ8K4c1BSM5R+60TktjQWsDJKkVrZu+6zMcvKci
U1nbc/riBKhJzlxYVAY3NKnTJX9sYObxnyZCeFpfsUwnIZOwVky4onrPPOQ55sEL
rOsvrpqXaRdbwx8mFaB/1xCjBolpyGXvb+5b823KaG+tgEq2MXwIV1hsQO3OUCF/
BFPLZ76LdvdH7T6AUsm3bRegmqAfW1LChwYLQtlSZQooiwVT7TaVdr8XLJTCpNY+
iqfhbjiWk1YlOMsR4BTWAJ0dy9imqc9gL85Pp29u/cxRheCp0f9U+rRBywWM3pLP
XemS2A2nLZn1p7hARQ/5cMyPW9YPtjsjky7WFONVLWt/qRzVuODjYLD9Soz6IAP1
9WF30384qcJwfwtX5z3PBxNU6kMmFbWVI3n7b2dImRhGB8TN/SMCKTBizpWyro5a
upcDiIus1OGpUJMoWe/4UyXwRVF9za/Z2TD/xv+W4mLJ9p9kTnJh4zsME6ln0QVY
pWuvVPJdfWU21YL/NonoxiieNP0qj871+G+JnpCpMfC/fbxC2GMc95T8LGw9qan2
Uds/TLGSTn4gqUJ+dfotvyjgn3ar7L54NFTYprVTZQ7qban1n0Rwxa7NyDctrdtK
WqWBxsEJZQ3xFxx7VEY0k6gegpELNAD1WRO3BxaUJg+ttLAVRALnkXK0AT5KKaUA
eXkg3s6P6BkOn85/oGpToyVpZJBCGQEhGrNSmhye1/+14VTK4dJXoVIb3erF8y38
wvxLx3vx5WCT4sav7jZu9ogXG6PgzQA2zkkaMgV9zBd7qks9Ru3I6qel3nrw3Uz6
oFDqgjL/8iNtj+f/+DI2J7P7DdTE7WZ/EKGPPhZKr15PnP94lGbVGn9tpy+u4gQ9
kTEBZ5pDMAv6+uNAUt9zyEfRf4miXOkYRDbBgHUy2LJyUrOyqTR/fHc4ADz9387I
FQz7oB4SHqUV26+YZE9wz/AkCVqVjzuTuK6HcpFfT7I6Npe9zGNpRitN/w2jrU5o
iDRclakgR+wBGjfiILNmm3E0lyhEnThUgsHAM6qTUhBebJmfIbvSJNVrg258vVgm
YU/N2rvl1qUJAzMTOHgjSzc60jVOApPyDDk+iPaOyih/z+6THsE9cRSQGOfV1HFz
A1WfQWSg7gsIR1qzV4pZ3GCU/f0G1TrTagBSKqobrqQxqrOc8ARVPvyfVy0VYUnJ
RSM1bCvCIAQ/UtkTz41/lNO6rGyZRApO7mKsBkGDImc4DZ5q13rIaNupplSVkQpG
koq5f2V3ETEYoWTO4zqgnKRzsd8ZpFZrjMmiJzqhctli28f2dA7hm+NeM2vDrraU
4FBWtxoEIb5dpeaC/RSq7cO0a2sbFweblmG6JSeAuDO/vwD+8T+HDb3R9FFf5vsn
Ed4M+JvlkUErO7GK+fvRFIpysH3dI7GdmojoH5C3ExiJR6C65fQ8qgaeNWoM60J9
U5nV8xeYHKUj+divv+Pc/lySCaxXhHRxs/9d8U2CWdC0Q3Z0/EotFA98DPmnH344
YbH4dqbSS997mBB2+USFiJ1DhQnJHxGeGfBKmFd4xu3eFf2N1ZcbegvckBxmcb6j
TD/VP34uMTfuin9OBYI1YezEcQEebSYZYPlqO5KyCgQ4UDrUhiq7skgXCz5yBs5R
WCKfEoX1pAp2Soifec92J5FluJyiy0HDP5foLYTyDWO1EECgnKHeBhSbdYYo3iVT
tZojVmfWQHwJJ94rZsK/axpqxr+L6Z5O9421amYnxdVXAzZDRSrKdwVHIIZBBJf0
YK1yOmfxx7O2jodIApjF7wJphyOW1c+fB2j2NCQmcrl6j14/MwDWNAWIeUDk5hNV
KWvvkQXTOvQ0K6E/0+l515pSlg3CT1+vbyC1i8CJ6f2SWUjxbnLNKVyh2VVT88Nr
/jmfYVgFvumR2vZP5BInKkLlpAuRnDvDEYKSY++NCMwtPplnOcJjX0S6td5Xua4r
9Ah1+IxIvEY5hVoqna6Kbv/0WnCKBpP0/XU+WYJ4s6GlU/+onTbrg3laVfSJ3EQ7
nwZ5ufcmaRCOw6OX+2ImH6+6odBpPM3iMVHpd79srF+SVUQcFClL11PHoHO/Gq+H
ZyaZB0v81EhbtnYPZ/H7VnHDyvYc1wKzdNTupYtv+b0xRdXvwTFRJsCPhN+2x6Jv
nSXKdxNrm52Fgt4GZTflRXGt5a68KX7YBPwHOjBtAb7/coELoe6oaM/J9pkPWkZm
n9dFwd1Vd52ouu5AFgR4vnglG1W3Qs0r17vqkWA3ePt6Brw7Y/NIYF7W7KGlZkQo
TzfWslynMkwcNmOUxFKMOj7UW6nz/i8lrMrd1hCTh4RYadbaVFQV3HrdovPpykZP
HGyFaC/8xZPnsRa3tv/EIjV55lpmnvUXAAcN0fLg25l+u7ttnXfizzYryx1jv3sU
TcE6c5eA1ng/kigqoiLWcA2dvUvJ0rvfJYOmklBKxY1wcZMPYJum0EujHOYYvYT4
dy1xlEWouPx2L/8Wq30rN52xlqy8IsIOoHa8lfRefkWAFrjYtgD1kI/VIe08VWuo
uifqoiC2XOojJabNKv9qBEbHBa5L3pG8P4j4Pxx5i9ROU+RYxL5Uas9r78EiQiiE
mBlZHYM4iJURjSrd3VuNUb3UrcsdDZvynsPz4sfnbjs61r5RV6zCXdnPYwlwsKlI
mGaDF8wJQwaM2v6rFJqtmBpV5DmL1nF98cG4k/hwrtj9+BP17mas6Yd76K6Ju+qM
3Vh43XgY68lmNFs2xwwBwNDwi27qrG7coW4v84WZV4iwfJ847WAIiQPoMsGfHugv
lGWUuw+2ZK9l1i8aXXREg2si56g+ZhIJXzEo+F3LtD4pKJ4ISonZa7ABuqGABgBF
NjGVNsXHgTSyi1MzX2GqyrVraWtweGAPQgQo1MPviXo9+3Dy/PIiOp9SHryqewOb
G6tT+Gv92Fk4C6O9gvI2/plCj6UKnxTevBU4EimO6F2FgkInbwy02aJo+KuLHRjl
h+MZK/XzR37+CpbXvznqHpY8IOGilP88Rqn/vW1C8W1pdJi+IYxwQqC8a08pKMkv
eacgOJltWjHOH5aRvQruTquBmgtY4H6l5PKnq9tTcisZnhl78HLRjBXVvULz1ZhW
kD1yTSX0rbJ/aDeS/++y4T0ntplNP036KdNjbUl8F0Hwe5nxFMcQs4VmQ1IDR1Sp
2sOIRYHOBb5EquWsLS/niyIQBYiarxjn/RXJ90o3xAOFErOxwndiUBNJVzFerPUo
qsmq3eOUQ9ML0I4GN8+grWN6v9SJU/K1+r/rDt453JhVP0FFtEqNSghCT1Ru5dMz
cjCBH5ULyoXGsGvjW+7UqYYShVn/edKE8fIJSS+fHCHUyZ97zSi6OLdcCxOPR0YU
+fRo0vpU5iw4d/QZPx1fCnf8C4sSFfEbNpGtW5lieWAEh1jp16ig0Ck82KDeCo8h
P/DdM0388YwSCXLGDkmc1tXqFKYRRwiF98zFoCbj2Jstq2GnQiY5gKXPd2D4NjG1
GgsGau1EsQZJQlF07dZrocX0bcKIAEtgFYxwxIiBYGhlXUeL5YVBkmiuIPioEKD/
8SVG4D8aXthUfnmlsesOIIlC8+lUCmUocFAD5Uqmgo4VdRkVaZWwoZcykm2z1HSm
9QKHRrHQ9GkKlh47RwB2GvHka3VBNBoRjWF4vsqlCCsTqDy1M6CsRb3TpvWMihio
eOXyLcj9EKYBxCDgH9R/lExQgvvRlB7EwccwUUyuqTjPtE8KYzHByhIurfWYjCge
D707LSN7JEK6ShBSWyZ3wGGDjpQe15VoK+iWtFgVbmsPwvU9SEmGvX8Haxo6rUSx
PiPpfv71M0YnFs3gbA/Exxy2XVAYBS44tQzV7Xdz84kdkSElfX1ZxX/oBMipRUlx
PxXYXpZ4b2Jg2i2SQgrhIaH3nZWS+qShtPUkBMKt2FNSSAGvPGW98NxOapla0YI+
OiUKfsYSkVuVrmWOHWGMs7rMBYGPcmZCTXMkpbAePKtZ4xFay0OmgRX8WzvXcIjD
csXf0pp3nyV2QcmLNJLRqekdUvKxnEdjlsABPTO8OgiTrZfCGLNBZJFUwV5Uk0g8
RnOxEhiOK7wGVCsZuVvspnwrq7iM15un7L6PSK+loi9FxjcnoxO3uHrasL9QVKUA
+s/rUBw4dQAINhOM7TCM87QvuTyD76Yz1YvxJYdd/kkrAr3iwKKTS8RvrgGOFy4T
btJ+lG+o3YoYkSPHBzGcuNv5fJ0TuwJyigwfYSG7X2TtmvzfLV5BkiHrTYRuh0VF
F89vP6pRgOI3FCLLAJxACklN4DfHI9YrHzsrVWVrpNPGmrNnOx+A40HFYEoTYGf0
9MRr48MqgU7l7xDG64CRZZ2w1EHLJlZJQ0QsB9MDpeOc/bFDBj3bKA6cffiNn82Z
m9gsAn9xNtTaAv1yBTFRCgF9BScd7u2w2rSwCpu/JepSwoD6fVAq4qAR08UDkRDK
35TJU/qnERirjXOUCqwlKgjd2BLwxu6ixdIkoLIYcblgJnSW85yL9QIIOU0TMswx
yBv+vLbOSHEIpVRlkiLz1tQfa1IBv//aQ639rQ4wYx1yAkJfgkdyaYlsZx54ybuc
og2iTxW55TtFFtwESu1k7NW/UF3uZUxi1yZbmY07e7HA7wxNVmaRB2OnOsO2dCDL
S5AbbsJNaAV8j8lDD6gLeZdEYgiOiBDR9G6lyJN29j03sRmptlba0E7erLDUinm7
RLIFop1iV23S5JM0WuUrRb6c9PB6d+YDSiyFu3AOIM8ZcCilt3+Wt/la0qFiZJfe
Kjhes36RIiV/SgYvH5G4ygSFl8cRgkZxHvaBRuCIfvlvRHvKo27/fZoRb85fvfRu
E7NU9KcLXywsi3H/s/CUi99CMotiZmbyHGTkItH0vOLhsVfrGS0o/7IB+wped/gL
HNC6/+elMPEixEDMHFiY32dHByCmddCnwoLKWKZoq57OS4RkOwjEp/LHRtthB2QC
028BR8wxvmv5jP82R5FacOe5a3CmStLCfv22M+yVEvwBB6eOh/hRJDuwK01AUW4X
eDXeEhvlyWL+LLrNuQnyY4v6ZDZ/Azknsg0fRfqVqQcsNWZSNE1f9f9hIu30Q5vQ
Vpk+DjmBEc9dZIT4Ma3KXhg5wlMXUVFMRl1VduneR5z0pIlfbj31dwJYmqWBn2xh
RnCB1WIIo0J4t1kl9BPDR5XL7Og3xWpts6IKOyo0fKqgEx+l3RN/6E+78rxaC3nr
4Sw7dVZMOBuYd/9B3OER1GtW6PuX3yn4zDPouTB75CargERabbQ8pUkNVUATMjim
DYPI+VfnmlI9JQfVU1hBS2ietRB1jkuJB+Uwj12CT+8RzZw+Ze3PEBc4NMxpfZOh
xliDHn70G4R/Fg29UeRm1yCqWGUFyJj30o8r8KDKviY+3SNJ4f6goD0IJFZNUaxC
j7nH1Ao2xPyUryJvAzNCbTcP8hKy7e03QthFT2EG5ZYCAMWMj1WikKL0MNFCapRv
wRpZ1r6BnyvK30cGrK9hL7DbkmcKOKJOcsPmgOZC6Q6O25x9gaA4icdkpBO7oYCq
NemXgiOtRkV7u4ffVGwF2H/aWkdq73Mg3Wx42rFElH825YoI/lG9p2gVOIKqYgaD
JZb6VhjTad5AzKAT6qytAGSCYbHWrVCGaqantbrvCJSOpHNmAEuKJPWHI/T4pKtC
fLra3SzfzKJixER4i9UCn0YNh2qntq5/PU4mHPsTiHgI2Gn3UoQon60l2wzR3R2O
gfCcMe6G2TSStovVCKxx1SEalpNyRr9xKGuZVG0ooixbojxcBcB7N2S3qBgxRSBv
2NgNLXS4FkSMypwv5gX3c/0alIWpu+y3jtjkWeWuBKC6tGMHl/u2zXTKzsMs1kpQ
VUr6/cf25H22BS5hwUYxT7pr+ILNzvJzTLSqprmkrjpwoUWLOvDVIJbx7g/Nx3UD
k8L5aOCg7Y3SbNlHwRVwheTOH/OwOVRvcp7BfEP7t+dOl2/SZbINmCRPT+yrZgrg
R06P9nQsFR68/dfLMuBIlsGgwrritFriHX7ymekbO8hvzd49ZiIPXVjLdQxmAWnp
TkLjq+uzJ44mRKVYLGbWKFJKEbLjVy8OQqF5fCZENgItewHooL6YXVdg+xpFGqGv
nbLiPZSWScP5Oik8p+JZYMMg0Izb3EJ3mzf1cq/j4KAVX3nOerNpo8Fj2G1gDHhI
UpaD5fURxl3K5/cQetE8lUcxYUf26b9p7z/qbwFyX6rBS/D236MDpkMT/DW9kAfe
cxjtM2nIsAFV/DMCZHBEmHXYFmqDl4Csnvv1w+hUUj8ZBfW9lFpnZkBSRwlzwlLR
w68oyCvNftZe7HW38Yitl+oxfVUI5ZksCznNhwToxb+kDtQK1EslcolJXmUNeFCW
guTd/SnMjv5kJoAVGbysjQhuPdo03zEfPn5PuGXQbLORdb3Yt83G2Vd7xmFqymOR
vy9itnlI8X9bhQyQ82tiI7cTbxFf/rVA/aXE3Vy+Kxth6wvvJYc6OURCVOd0HTR9
wr695XtFvYhZmjcmF21y2W2vsVvjY0ddiQ/WLIiT0XDnWnLTFu5L3fxqBrC5+IUQ
PmK3hfyN0frKoINVxUv36buTGiqZNaYMXFhdsBDUhz5XJkK5HVnDSpHV8vk94ZFH
3QANgOHMJEgl3Fm2Ls8oUg7bLTpUNM6/QK9Gy5AXdarJSbQ5G/++qOgpD43l3TrV
exhAXaT/0ntIaufodBRng9Uh/DLLUEMjR627bhuOyF6sgxhoi4lMEqci1qhira6P
6tIq3If3BE2ci2RJ5XPjbWc5SbWmVefp7gSzjeYR9DGkloeF0WaC+2iTEPx8he6O
VNFQnRe7bIUv1wjvlA2fPpUReG7GhBGmkUAgp8wm8wBa5zqopW/c7YU8llquoJQW
VyZIztSLrIjWKwTz7X8YRcCp67KKa4hftF49ypiWrsLDn4gXDMOXOLwGCsRhbF3k
rQY1MsEZADWq7KnCarkEUbBixowEWLhG4FlhwVd7c/sQ7MJ/U9Hfa7dyYoPH2qAM
DTNosUkIjOoJH/Ibh0EPuNFp7T6hcMhyacnc9IAcOCQ056h7tcGMpiQuDLYNObNe
JswnuZRsPbA65FJixhBnthmcvrFY07bJFsJaWHG27hivjd3GQwSPXlsJYrCKKkUu
d56lHmyq9AGgOlk8sxljzvMQhoZahX0OlET1MXnuQE86oYz4ulJrYTVB2WID+wAT
8+sUr2Jq4wa0YOlCrosxwFkweWkcelsWoSgVOSIuBRCKQ8k0w6J1w5Ec0mCSwTk+
vvMNTTSo3TRKJUIAQjXUPkWxwScwyQjNsFrUVS9MFINnrNvqFY2ru3xXYY2MypN/
+uvcf05uu6QqTarzrRSgo4Gbg4PUlMEvihgwyKBYamtDzynT00NXEv+lajxy13VG
tjQOZCzH6lvjBMpmE5TXdxxK++YaXoDnfrmjXgalmpyItXXGqEwNf9lRCPRTvmFQ
L7MoKhBZp7Z0nh1BNvcJnqeCfvcfm9+3+4W4pwnmOKLLVztc0lmO0niFEwjfWb4u
Hi3lPj4dCJTSwyeACED4l11hCxGweJkIdEwo2RnuyUwQLDmKrFjrZB4LptqWTgrM
LsabRo+6CqiHWWLaF9ShQGs7E8MReGFlV77dgq01GEu8s8MYNquzrDGC9h8eXmmJ
D7+aCesZLJg07/kwhrgDVwD6g7UVc70w9sO9F9yS1wJmXPxZoD3aeOlh6kojPL8w
7bEjNKvSrMT0iLgHQhymx+uL8y1BqigTUV0pctqsZJc5FDI2vez6/l3XX2fMjE1k
l5Pt6PNOEtsnmdYNW54s7jWQbnQSpd/9to4kc2N9pUK0UvalV79dDAyPEmas+LIO
LtuuWYYO79vj0fvlxoW3DU22369AQd65LF4gj3/1ESOdB6hdLMy6tZRToYNcC13C
rppPAUNSytj4YEMOZFdbcJcYMpMlUgdzwtr02zehnxOqBcgdaRtE1B9eIBire1A8
juJxs+BehaoOoeKAGO24ADay94Q5YG9tZ1t7w4XzcaoXEACkoK4sd/ENV+lDdhml
lzlGn1wzCrN/4qT5yqfkZKOrRZkZP56yxnyvxVJt8BbQmP+zpAoItRzs9MAX/psN
7ixlpZT+YpJP+4BVLiuXYW+/Fk58pTeniimMsXeySMVF38W2Ruh84wI2HhnY9BZm
Ekkbn0ZxZS3GX9PIFy416VZLpBfduDdTAtk7jWbgsU0SqFAMOHmy7VaAfCfwh6RX
S3yOEYHUWROjdw9ObwWgDWM3rGroYakErZzfzgd+poOh41abhXx2u5hy4L5yYGNy
7vvOBCRgwCPxseUbM6Uwiy5YfsulnA4KXMdari/5YWMXnBTg1lyb1KUKP+/M5ppY
3eyaW3L1BaKr2eJpDGFE5rlJl1K3T08/RzaXCfpwHdwl7ZB68zaUyAoW2U/vG11b
D0Y0dfd4NsZcTtS/hgQ0hDbdRHImDHkeXJ0ZjuuRloQZe6pkDULKuEsvKHyqLNrq
8w8hy275S9MIcytN1wiWMayPVrtS+5Sboat9+wCtbBck154yR6MPMyfLRfogJKim
8RJ2ILUUm47UXQBRdqkozcumfSKK/5Zklmo0Ijtauz4k1K3XFFGnnJSKJ0arzQ61
HEyYYUPjAfXR67b1QwIBlafvyiGzv+2qkXAelx3Inq6v+8zMjNLI3eyUViPkC+6M
0cPYhdyxg8Gsjk9ShdgiMbzfrrPNvF9GuJIHVfnVDVxwA6wX8cHtEwkhbQPNaYe8
eVmpkkw4MJOBG8IpV//TlNwr5yrCtccuXrPpI7Gx1vJ0iErvaZEiufx0pgRpRcmR
HLdsKoBnXHl6RpgGU2YaTJsg+6iWkZM/B3zg4wphrjffHTkktNzgy47t/UuB3KiS
UICl32J5tXkCqDyiBgvEsFyv1Jm22U7dJttuwwYuxJsnjGaOPNdTJ+DC5rL0IgUw
gHt5e5+mz9il67qRP2wzp3Pj+jE1vdL6xYLCwzLCHQYYc9y8G1KPl7Th1kE+ejga
I+OtjogOOO0MWBFGh0NuU2wOCT/85tGX1aSjUUW9dlkyUPuiB/GqbJdgn21/TSSj
hwxzF489f2ak4Y5nZISlbMUWHjdbtN5Cdrp1002FlZu58gH3l14Zwlr65DUwzTPs
kQP7GvPBGlKAd4wbKd+5S1b9jUqAWEg1LhAA+2dVhuXJkpMwbGTxcjXoQf+C8Vtf
ORys174yJ9jViOzxMJyiENh4TYZFukOyfvrxPdOsBPIAFTV2TR6G1NZUmej4/kor
NlG4kE9LOEGBAHnISw0EzqIt+a94CjzxVSEDvUZiqmSdgGNY8Gnc6b1H26fqt9HE
01f+XOL2OF0S6MRJKgsFRK0oNipL4fLy/LOFHTHXPYjHRCXTiXFZAdcErrT5OJ3I
AVfKDU4Bec8dQtSNn58bFnFYU6FQ+Se4/Sb18ggh0UOqU/ZvrSmYWraZWisoIhnE
ZdaGnCPO9Avpde1C6ffRHk0f7fIILZeXnu4cePvqhAsb8ZoqPOt9UQYY72EpFt3v
iOdo2rZD8dyOuagqxTz6LFT4UWqfMzqh3ADe8LmNbvfPcG/ODJcqFVEBe5HarM5C
1PpUnnZCrhOhQUXEnWtvtC55ioPwUYgdyuVRAGSRVDmsuo4HeN0jjva2Bpxed/5E
HvVfmOi3jxlQJQbOCWOm2hnJddbC6yIsbsUPej1sf9ENMhDvyyN7Acp1+dzFQKkT
Z8bA8ZVobKiw369eNEo6bdLXmaTdVa+ITD4H7hi3j/s7fjReTE4M7RNvuVDPRW0e
vCO3FGjhrdGfQ+K9Ed3nE6IPKH18Kt7ykxC8DXH3m6c85b+Bc81l+A4MDl/ewxeH
PC7hAU/gTEiZ7GpYXe6BSW7nqdYJ7HkvC7D+qgsIPntdkW9P/QRu0fpQkbOK9LE3
QgUdRsltcFYegenclzq5avwKIdaSAQIyrxRx8auXAV7XHzVc8Fj+gBFuxahoWQD5
us3CjOtZ714xd+nkzLM/TofkMd2+pFRJpFoE05f/svq7qgLEzZaIf7ORx/u8s7kV
OPaRYwZZHAzQ4iBptfX0ZcGtfXkLrQF8Zjw+07KVzM+v1JFsfvNJAJSk2extB2EI
gy3bbsT3A+gxVqQpcNkHRs8wdWg5mV2NIL6dixf6eBhuysuL/rhLQ2na0A3M4CJI
kEvUAf9tJmi6KUFIbYj/7MVI7BU1C5h/xug4bwNjZftk3MVGU5KSdCEf9PNDWdcC
95Wfc6PBaDEr6bhF/PXYg8DzDRDCvsIJn4hqOSq9pukgEVhL3purPMBC2ni0jFZZ
1V00Ze6d5C9/SbnTOcvDWO1BMRVGlunEdMNgeBzwfZpjgeXqp++VMOfDB4Lg9sHN
+buCws2LFXWg5EkkQKZN3Trp1Ik5RGlBXVUFOG0jmIdb+y/jD+s03QC0sATpLaU8
kDj+oOp/Q+HY631r8LIFJjBruY+j2an+H1UUkTviPt4Ux/mHjYIAHtrBsn5fS9oV
mRGLmomM6BdxPOOGD0xyE+W+iC5e9zEDgcwbyLTEnI0GZengHBpOPx3h6TP83Agc
+bFljwayNmKWGEDQHt/QlDszPbUqkY24jsnsAm+IWtnePSCzwiDZfYfpGOAuqfz3
y32QRn4nCAETyCVNnpGBDuXMs6BTsy/pb2jksee9VXSMtGA7RAmI0gJz10w5qnXE
HvJ4lIpUsmTjRI8g8Vks2RZTndYvX54Z9vRfqzvffh7xCETOtkkIX6a82fzdEwFI
KLBPCNm70xFPrhfbcF4OJwFUlD7890bkNPM6lZ0PwlKvNhQ5H3j+tlGc2Xq4PsRf
76u/tPKNrbKZx5eNaJLciMj1lzg895tGwrFVUHDCc2whw/6abwZ6gVPvssklErkA
75Skihi03flDRCsOxQmHOCHX0y4rnpT8bwAU2mMfGCdjrJEFQCsb1OLZvajegoIV
ABh6MhulW/0bc17vmsSDDWXppEWMpr/L60D0RSNbTtDYzC7Er7XecdmCLy5+TuZX
tUFuujnH4dwQtg6MbpPUsZ1mIN2Dki54RQ2GaJ51BaRIXEBjJQ4OHKNf9gLBGQog
LpyeM1cbqOnFsH0Y9dH3sXteVCS93XbM2U5gNXOYTtlHjE/QMJkdrHXRd88IvKsO
4ehwsnDbMzUZBK8U9XHuN/FtQYa4OuOQkoO9TG36l+GA8whvDgDPxNuiv1pX2Jp+
/zPo3OGgbPXnmSN52tqWB+L8c4KHz6Jw3DXYfZbiURV1oHupEd+u+DpwWygtnE/e
OIjZVEujm0eLp8LtX97QhYMb1pcbPGG/7E7K8jQumzfNStNkYl/K9fwr65fGFuMF
D1DVprhjjay7rgJ8uL+DhMjmwT2QFisrZhL+tkaIj5C1MAOUACAMs1j02tSSIIw0
fC5hFErgAnLI8wEnO6aPaB+ButF4zaVndKbsMHl6U04N9GyCbsigX2EAvv99940K
Ku5jwMD3Q2hsKr6F+vDfsjcP5paJaYDNft6aeFW2VF7hxSr0Foy3pS6z95bCtTKh
mBh1JaLhvv51mwvevytIReVI1XIfjpzehsHqlf4xG3Dm0jCCarIXoEX71jksTrXH
1xgntZ8XBrYEKRdwVfun6wnDVpjy3SV7vxHjSjRjycyx+xdrE6NhPqvr0Hk5xFHg
5XSqt/T5OY/RpbcCxoa+UR/BQ+tdqVZtUnhIX2xAmPLz8MRjc2jz3OELT9T77G+q
bi3wAIUzxOpLBlqSeIR+Ma6FwxfCw8UpdMqp0Aa70z4C1ziqNLJuSX7+mmdG3oqm
vBHzEwBKt9O0n3nLIp3n6fpaW3i7TB/twapK1e8G0F4Oiv4L7qVJ91z7AF0t18gC
dhmdOxpGFl8HLwmCVSzDpxvf3j/Jp3NJL2iSlsQkG5cRHzD9+2fr9s+eU5R9X7C1
pGJ7Y6SKbJQenscpGDN+RKDZcvPQPPVjpz8XuhDh4g2Tix6AXD791Sq6EUeYosWy
TmA2kVt5ImOzg8fRR01T56Iaz13qhJ0Gu4cKvCQ9byjAK0QBCXv1pRVyMvUiBN08
kftpPfpHO6k5zjqny8cIP3mejb2LOBHjksZM/eMbBzQp2BJMOVQczbxCBGWYyxWB
p1NdGBZsYS/BJezITbq5ngesUjFYrYDGGxIvZXGrXyFITuZk7+zg9JFi6Xd7Mrfm
xgPMOuLjQ+i1PwDcrTCe99dvKpvmkshtOnGs/qQDsCXctBQGdLWf0vd9/k7nHf95
r3vs038F4T6WVNtR54NILRRrVcifQqQWlzVgufOVPTl54fjxdrIV6FXF1c2PMICp
g+sM3mwnDl/n8Sw9USeYaxe1JUgl9bfzLo0fYAC5uIFvqFh2uh1WNgS9dD0YGzSb
nnl/ktZu7a9E78GVUlAwmrgIylW8FYRgw6WzzdOhPtxDOyFJkTel/88NelQ0giMP
AMRqlMjqjd5sTUFKtsyAbkOXf/4imB94wzhJggyUCLGTLAAmqlRbAi2wP4ztf9PT
S4kGQCOXS2R9M8JFICT0KnQ43kluq167VQezLyZPGH0PgeDyrjxwjq7LRylWqMP5
om1FbfNfq66QOm9jhVrTajIKHMtQPqQCKSexEu2x+nWnr29JCOVT9cpEi6C3IaTO
0iqjt+bp6usI/kl99tDC6BqF1pavXC8Do9Aa2Y3Ug9nik6JtpfQbmRLrn2M82wth
+6Q6s6uJHaZ5JEmEHR5gklTh0qnHjJ6grAPn5+NSZB64Nw3wJ+950y5032ISMIY8
3u6bsPuLf1c8F1dakKukWU/4tczTyZ596EwzRfsH6rVxD2h+fFBY8YNI9WJ2+AaX
6TJ4b/Lwez+KwhU65zp6SfNefc+tbUZeTfTWzTGuZX67y0tFQBnswPU1522iF6WC
5I6IrrTXb2v/Pnzdjw+UqmV+8rugO9xbjFDEKwLNkVZtb51s5cw1NLbX3qy22lPk
jRX1u0WH74blw5pXEKX41gEAkv2DnnHp340SuqhHdZNHbC4VtjY/Q0sYXcrKueZp
ORB6IIVsSg3Kzgs6BnRXZqHMX2W+AaVHo+5MGv4nEWiBd14TTw75yE9l7E+rleJ3
G9j4XZTmS/dksnubdhXA/nMaLxqxcIAZD2gI+FvXCljVqBRdgg86SV1YAw0GP41G
17hJ8OwNRbdDP5ziaPKI9mOW0xk9Z+hi+CuPKosOPH3f8/8W9mePJPBxgz7vUplX
tp8BuOcuTd8Kt8x95/qXThQOzwVUBCkWTt2WLBsx4Qykyld5YYRE0Sj1UlmPLGDI
FVWh2cQzFA2JKk75/x/qDjDulAKgXRGX7FxG3cnfv4TeNIzBQtCNkjBrFTxWpEOf
uS2p2zH9L1HXaoRiMoJIJaEvLuFlCUOVH+5xfdlyUiDSGpOHr1rOLLoIqE6pMMXn
Io+Sv60Hhu8097NmZl7F+KnKEiuCmlP5kEjz4FVVO+333czHiTFDB3gy1GPlmtGF
u+Qtdm5Q2s8LHgKvM0u0Qf3eaVc7j2IZKwERhu1aQPfVa8PnrfMVhz/e6JEH4RwQ
Y95U/E/EkW6hEE6KGrblg4YkaKzsdAOClPYHWrJxaqdNdK7sf6+3WhzWOBlXYnUH
euEIju09Jfa9sFPVB/Rv3/z315m8Phuh9npMmuX7U7yx938E/RfdiJCMqFYBkyv4
wYVbyfsSWpX3kBrTs4JHNFEfPkHCjMAzZAdnU85noZcxIkw0nf4zPmrZghMqbEvJ
OLPkIj9KApOVc65OXJ8rmRIeXbWGR8UbHcAzn+zBmKKidV9jI43iIV/Li2OwEpmh
5oPkpFVJq6obPq0p1IJoAiXQmChhPTrzRcm3ozUMvKtQsZTh7TvQBtzlAhD1HLet
vNwq11z+aChtOqzXo8bEatRyp2OMbveBfKLnHwnRiv48LVNiKgJTVpo2u1vx0C4v
GfIEVRJUse/vA3EIKA9IsrgWpzkKkfCZJQgPrrnZ9KITR/4R8ziFDG+2athhZ8Tm
1K8rytT1Sdv0LpNxaMy/G9plOtjRt0yR4UcweJilJ9DBcZpeGBJ1uy3hLXSkoOVn
EFyxw8OXefz/vLzVufiwfTzKkguR1TMN4F6r13PnqqUVCNtTTl6jUpVJZ7krJrSM
+PLTSTMG7VHRpOGy5/saHYy2wZGRqRoWNJiX0+MplTkHyiAFpvDB97vb4VFWoGn/
BFN96uCg3twn/SUJ7Los1hRS9oQ1ylPoxTINTjr53a35ZqtRG/Qg7BzLC3zuV2RK
i+UIJh3j1CjVNieQ7ILvJsYV491sfYeWoF+sqHTOWZHM1juLVD2Rqie/AQEwY+Oe
QBis0jmHQsLStTSdT0AjVEu0aA6EtlAYjMLFIDdCGHhDPjRIRSwG9GyE75ctRMAM
0lRSGJzixQkjTrJAfT4X1YkWnuojttz6Tue3kQZwSBJ6/+3Qpjpqa9j8HIgv/U9m
79yWnbAcQna8CPO3xOgliK2f2a6mrLttM32IAbYPhICkOesfjnU2JqGQhZf8iWWr
eouAHE43qxvLC8+OD7r6GK8oxyQSqxylBKULNtw3bMnGOjW2TfTA+RvaDu2TbiGw
Xfyr03BMlmnRdA3UlJIUkKCaRaKnbP3CEP1Cjso4iWpeJuo3t/O5KId7w3jb6ke6
Q1HHKoYfJWUNsJtr1b3n4I4SuaWxUOyuijphwuZwFvdnJaz9LxlxN4mFamDGCY4L
LqjtTfgha5SjnvEbq78vq8Rlv0hsIpGOtbZub1gLGUzXozrdcHQ1OfAmXLM2sWTK
uz/bxrTsJy1U1MMQOUQUf/h/eknb92OWEw95mAEKeUy9mJ+gD4w3XYW0tdqSu6bk
Cg7TVzWTcdev9k64fRtvtQZcuPDfNg0A3UaIbT5POy5knnLZUlVsV66rfIZmbO3P
ecFKSsOBDtK/F1o9wvGiBzlXVtxSJgLrnWhIJr1wa3e+Y6lPObctEEMMhkWAqA8u
/REzJYbZkN1Q+XazH5z0TGNuoYETcRbabljvAGWgmgHLt6eFUblTR1g18Kx1ztE/
vJF8hnkc0jV24k30c6ptSJBWZtUUMjupPwN1KrQow8OEpUXuOBqoFhpC+1uYhOfM
IqBgC7HYc61F3sReBY81MJivXgm6o/c5uHDApHrYmZFaiBdNrN1BTKfF2cqMVfO6
wzcl3ojzcPwnjwg6AZ9LvbJC2UpStq+rdC7zM6BlY+2JqBMw3Xl8E14S265q5DKd
N0Bak8JADVm2UtIUJtbmv7g5hrTSUNhQi3aDNE/Tocn1Pa7COSOoyuEJ/Bec/aui
JrSiwCIJidAfGrTwsh+i59FIYecarzTm6YHjXGG5AGqSv0BtkeNvNjOZILXYsJR5
+bOhzGisiFAxtstiz29ECQ4Ma40TAvkqK4Jok+jltgtVvBC5bqD6XPpTvjvWTsTz
szqEWfczpXIkckzIUAAGyUFYtX3DV9RiBegXm3TomtDql05gkiXXXk4brv09KLd/
u/FJyb/Sf/e+veAna4J+S1gNj2KvZBCOe1/B56VyHK5qdoO6xk78o8R4vZVzLg2+
plP5zzIPMPgCQg2K4ntUL5bnh9GtHrRGPQ2hy+6xBdFlRfFe3bDcKoQCfb0dGeQy
L6kDe3JuCSXqZ40r/lDD1XjPRozcxrS7evO86UAAmQUKZq4aOFdyvMwAoagjuuDP
7+D1v7dJ3ZJBl49iqRhJizOTHxu5L9dSVtEbT8NAsfWuVklVLQ3z06QSCGMzf1hr
MdoMouJVp8s313of+lGZbVOCTRuJKaK6qJ/obJFgws5rmvcY52NxhAgcTXP1UP4E
304ofm4Nd1wWIIQQTtMyUUUbAprTDjlgOmEC5aeyDPh4BKdPfoGNAGATUKMOJSNT
tORV3DV/dT8hyOLosxUQa71/DqBXaeEZ4Ecur6IgIbRlZxQDGnbTYaku6Xp8p/cD
M3mPMptKAJGtti7UR4AnnadVQ5FzOCjpxqVQj3ZKEDGQU1QOSeL/IYqNZIIHUEby
jnOFkqytGQF9RBbMqvhXJJbuOmnUzIiQgS0YkXHlnvDBG9sjI5Qzi7TYhJgqGToB
YtqKVT1RmQ0eyqgN+m71ns5GEl7f8nPutFRPWwvcxjZIjw11u/EPXoaVuzGwF68A
UDCnqqGz6QCwDKpUZrEU8OA116GaphzPh/cWG0zf+5K6nx5l+mLcwQQC3ebI5/KS
GaTx+crGN1hP+fwYtKUmpmw9UQVsM+HXwxlEVqXpJjYnaoC6uaA6em3mq9vtl5ox
bfGeApp6WYb8T1g1HtdEcPHG5T6YGb7n0PwrUUReQDf4AyuocLmz4ljskYqB7crd
0pU7xAeB1MsFomlGymf/qz8WezUytzv39t6iUnSZnjdVUEBdQAD9PQHgASDAMSN1
nyUlQMpRQRDX3h2pDoCly5cEMNZLac4Ua7zLrHcrkYsngA8xmdijJmaRbd461+Tt
xaNCjDKal4gH0WFNRHJ8AZlnxaMxL9chJMXJP7cHq/PRpWlZ5mbooC6MLvbk9tiT
qZnbde5rDwD1h58BeM5z1r7nQXSIxzTL4MmDJKul5ZFRrWhu8nvYrdLnkNu3EiLI
NBWi3874jjg9b9TmICSzFVICL0NUHYpo0HsITrXguHxAOcGUNargdN9SbhmNTsiA
SWpMiaiKGy65kNGbNMR+Vkwbf0YBsx7cRSDZ4eYmPueAvymEE5rqgXbgPLt3uYvT
ibMzq1v987CkuQnKBHPoxubKCEjEKR8pxBFMKq3wETuMcAEMVaw6R1RZ5pni5/mp
gCC2GzjUinMI6/ym4uHmO4bs/UyU6kqC5jV44q8ARdrjJwaBle4yrdj9RXJ81J75
d7dQBr2s7pQ9MHi5St58f25Nx40bzskNnPSRMZ3b8E+xjn6FK7GshPBnkzZ4JhPD
KIiEPd4UNpEVwV0VCo0JjzCu/3ylz0GO5GZvMmPvtYbGdn6ROZLWjOn6Rnl3KUd8
OgRRecr+MiCOlpV5ZKeqVNjGRC5HZUwC+dIlRKJHzbMfQehdrABk7VRNg730rVnx
th07PbcPMCr+O+oxicxWF5Y/5aq22s6maxpVFtAW7R0ZsCmDW7if885L+oDXsaOb
LW0APTs5QVGhMmKprkmJlGEad8jpfs0RtjxAKF0ZMiJrVqzvcXJM8oqLQHV/+EQ9
4edfaNCuMDsARde2U76xOrvYGjwflJ4eUVcUvOms4wHFZOx8MivCB733J5zD79F4
EGuSOLUD5W9vXfNOwbUxcMy+V8W46JYdGPc692lj8eB1Wmp3YHLqniNR55f208bF
2ipcWooSLdynUCDDr+tt0NXj+UYT6UwNpt4OUMFIVywI+5KpW7RnixPwK+KXOiY3
0s45J0RWw9rN2f2SiwGI2t6QzJxoJYOv6ZqhzXxdRBDM+iHx4vJar+d+tt+KYvEO
lbf4nBkflGcZ3wXApQUbGoqGVNdl+R5eKZuqDexGZfkqDTqLeX7H3KvPG2p4+3Pi
n1CDUP43+rbWwQHnulvMoyu3g6g1Ch1uHkHcD7YSmIwZ2jqi9o+1z0FUnpPZo2Sm
WrdQqDGDfxqz0pa8zJ0bUJz9h95zQN1Yui4ApvC8D7sPBGBcWnYsWoJR2LgsKAbS
hKN1KYoHqcek+fEpdymbdv32v2gCNZfd260XlHyyWtEqe2q+aN/DBmmyTnj/h/XB
k5R1Atgell+uLvq/QXX8wIMLDMyh3lPoduEmr8LgHFXa3617rgjBSyr8tqowOTqg
F7T49hqgnCws1c0Sd0Rzn4mcn0VievYe2rE6FA5reNRLjp5NfroaMH4/9YCnLnX3
7lkGer8IbmUK3i5juYFjeZ7zdG8deOts2knF1jgfXtVZXmIsARTnQXnRFRhP9KJI
gETkVyfQ3HNqCyiKbFYssiii0BQFImM9F8kJjSZtm5CHJLqGoeOt0qVgOSDqcgMe
brTsdPSRd/gaDIzyx56G9/CKAkNcjAThQ8TLJGn+RCFU39JGW1YM2kCTgRAYtPWZ
M1hQqUdZGpCkER4u0Vp3dJwia4EBr9OZXxIfAOZFYwtWPWzM9QL8ro5b9jbx5nwh
eGx+0xL0nh6t4gqFDouDg4dWK0n+b0FoXRiwFFj3UYRb2NwC5rBUCTS1xiT0mroO
B4cu4qPcfLnhpwcfc+De4xpcWZMFIs4qNHMjaUL5YK4rwDQCPaLLUugPLk69j/6t
ndNa+t+WLKvRqMzkRTzpgusxmZsNDRIGHxDyntnbXJLu/wBrUVa07fNhAh3acpOV
P6lhbVGfN080/rGhyasOiDb4uvznOj5VfBSRnUaX5hQ+UdPTTV1ukM6D+wndbULa
5VW/HiugyHs5CTdAlbrQ2mmIxZiJN42AFDMHdyNfDopPOBQ2gCjM/8vtbO0wRdO4
CDCApRrxaU3zcOiipeYXoIqaPF5XsCFJYS7uqSAieIWhupwesYgceuVXL6C08C32
lFQGFGWmPEVs1e7JU4FVK0w9DUzCiyzL3OLlAn5nTpunC11pC673CMKpYiSZ/J2e
3dViHGNTlDGH2ynbSqglKGw9jT1H4NXWdOfed8PvIEOgQukaIsJgX7P/FWOPpT5T
4RzGlsGjJb0k4TQAxPX7k3MLHIRGd7yk6g+vTXm4d3XulQFT/PS5Lh113AAjXITq
EEzS9I9LoI8AMuGr/m7k2gXOIPxjFG81oLNIUjwQvlQXGSHQroKaCvIweR/mlaKl
SgV4PVmxSGOxa0vOAu6pZcr0jkal13qMyogz7LP1itnsRXUX/N8tiLzC156I8Ne3
Xvk5uwxOOQv7EcTp4kkxoFpdYjTlN147iOrlCKrzELHmO+VOiSxFO/bPvutafbFd
Jfc0bhAaJ7QBrVAEXScL6uzBZ/MoYQYdXwOFivaF8ZbZASa2KW9xd5Nh2aa8rLUO
oGoreaj/ebKTU/mgoslC/QFaMFdvm11XMgyW3gqL7tB11CO8J2TUADQT+qrJQLwx
f7cBFzlwUhf3Ksht1ypZsz22xfBoKND7qZJYwgC+QibwTGMYDPTH6mS1Whmya9Lz
rMtBCSVbu/Etvu2PKNXSG3aWs0YTrk2EIjttxlBuYipq3N/AK4HyI3BymQ2c1Axp
FHuSmFY/NetCZAwPE307WZPIrpOS918sBnSSUqysltqV+WvHQ21+S6dXjxNwqATj
cIV8OOI/MZj/KV5FTNhF7MNKnL9Zwvmg3uv5t4dv8BvwiSY9hjTqttfnvHck5eQw
kY66A/zIx/diC2zjoIGSOAryNojU3zE/r5NoaCkvXnNboX8V1uWflRIlERN0bYGN
YPqKKmUjua6585dVbttvEkQa9/dbCf66roDGckMfxleXugLg01cHqFSLnMYoqHLU
KcdoFCVdRZFjrvL8DLx5ltupKLq4spb5Ol/X9tyxhwbVXJmIdDVpm5s/cWrXHwIY
nf9HA1apxJlkDV4qa8UzrII+t0GNmH8XJluQYlNU1EAcgNQKwCMf9mRdgVMziSB1
BGvWsePq/uGDGm35Utu//IvSz+JIxSZGIcL5u36lIZx0Oy6RTSJ8+YOvzV5iwAgX
/7CB65COBJuQaqkKaJeq37lLMw00XOGkv2i+6M2bqRgI2Kjiwbno4OYqYEfkxD3V
rctaa0d2mWb8hGtjUIF1riAc/2LMk43GBJEtpKXik9aYOsD6kIwk3e7c3Sfs8lPs
TB/9g8+QUiF1YXC6ZhF9sNWAmU+LLb73+dUMkZT2fGFRoP/Mr6ckxZ5+Oc5Tr6Oo
LKShlXmnKGMhp2S6TXBoSCaNgqsG/HB/5d7EdvA41h0tC6lOLlhlAg+ASY1dUE3E
serY/V0siJck6Gc3RyWZbbfNHaqxBbh00zU9dxcUqUftvVXPRtvhU5Zs6N/lPdgI
N2MBLC/rxpoMZmeqUGLyxbilPb9i1N3Gdf3A29kBN0wic1r+QSqkOppXWlm3kScS
thKv8IhBXiW0s5uPsV1JlpDfMTFGikP7SbEDTlmVHmm63jNO9Iotbc8Ch3V7G1xd
Tx9O/5MmxI8zy4ckwsy14N2FQm3qqU57PlJsTO8VZjkUePZ9JTH1yqULF2sQDdf1
xwpgPv9R1cflo+YMiRlyazb9EpDsSB1w1jlDDtZrFlPnk+y4VVZ8Gt50fRCBXwsD
WWxL8VYNGgbQOtd9rXBowQ2sTuZNnSkw9exUiRP+2zj0xYCxQWpx5L1ZTdZW9s7n
1I/RjPGFQCUTg+sHH4ZClVJe9V2Zw5na7mBZAq6IlemEWf3+/uZtqSz5uvfAY54F
vA8/P+u2fUTmySJv2w9bjCrzmA+/ST9wgxaQrleqWLWg7TxB4RQ4yTCTwM7vl7f3
2PYtOaRkyuthPBMExpij8CUR3sCpJ13F5gjiXuwqj2t1+MGxfXINzo87RFZFq87r
Y3BMQnTiGnmToXZgF2y1A2PnJ79GYCiSBMxKyawi61RXpMxTf0eLUrFF9tec4sVi
VMRJ+as8V6pocjzfyU94QeWlaFlToKymuKAgZ7Hp3hQ99rwG5MGhVDFncENx6ij6
qk9S3z8o6dQO+UOoW39PZ3PRf4hV2C99OCiXI8tVhxCI8WG6HxAmleli/FOfytCP
pt+jS0Q+9VOkZZkdMubDqOcuJeh7eCOz15SCUumrcjoVQsXSkECmW4jvmyC4SVQh
xjjb5GGzwLrtzTsoKizc4RFksqxMk9AYNipngR+PmKCNog+VbfqQPAibZSJwnUtz
wgBTFxtq5F+W+eiN+0oTYZFKzw6qwVRT/gXzRKMiRAcZsrZhQE6OYutZ+uAnZBFX
YKmaE1w93fCFW2QhW65aDmimDQ7vwPBQfZDKe0dT1WB4yRkj6gEoos5VoklAtlAy
aLslyIfja2taJXLGhz5LkNuXKTtnlT5rJBRzUFNkfwwuS6/IO+0/C3u7oaZbrHBf
LmZBaDAxzz2xIa8cHrN4+HtNW+UAzbI+1t78mMW0x0/IUH5EcPSwIxx7mkm9smAS
ri4UT2lTW0ZaqWhKgLJSvE2PfTThB428vRVl7aQf5CiHE9Vdi2GQvZa8aXQQSLra
Nimtmw4Qy87ArrWGopnVmonWau4B+SJlNNJITZKwmS9D/Pygc7aQT1wLiDhRHlTX
Sm9AEHTL5ahJnZ1Wl1qZ25vQhhxeGyRXi6aWuJG69EIvzHqErsGn0HRfxmkPz/cL
LiVOL8Fe74PvoHw65aI8PI0XzMeK9j8ImQ282vOgSW5bDzpG+c5ZeCUrUcFdCIpG
iDVNDYn1jFsx/OCSE7/nV1HcJaYgJQ3tVE38eSI+zDd8AynxBfStaNxTI6H+OTU4
H0OzEQrRXBc6UD00Vtrsg+gBosDADdGpLZNF0uR+uqSEzwsuRoS5S2rzm+VOqVff
eay0zvA4LTrokmvlI2rdPzX+ilHtWjbuzqAn0/vF6gK78SrB9Zwwx9Yx+Xt5rYWk
fgc24y/si34UKGrdJ4Zj9q2PbRWOyQ7dxYryN7jerEkAd3+y5vKD72zRV5UU7uep
oxFGn7mxMv1r0VHn9hU/0JEfP33jzpVgM+J/nULxyjkUPKWpQJMXtdCEoWkXO7Tr
Q+i7ZxzxGj/b+HkmYSs7gPv9NImUPi+8ww4IibS9b23PE1I+dAP+S5SgU5IpwCO3
caSb8wqTcmFIQhzxW6bA1RN7q2HEANUHENrFhsUZpySfOh8YRR1bmpNkAoQem+0r
2jEdoxfRIKsZXO9tTtzgcu3YAXx/XSj0ELly6Uxl++yWpf1jYt2eYK+WrSNXaZw8
KDA5Oa9pB3G+Xy8KskuUvx3nMbnAKvF4ZDaDMK+pwPT23S1rLsd9edtO9KEbe9+3
ETlWmN6pJvSm9yACLta8B5HU8VBXv8OE4vU1fSCXjFH0k6QAdJt6m1kvpRgd6K38
E+JOcSrXlHbaQCJIkIe4mu64jryedN8k7uW3+SDke1v2+hkyDpWsEf89QYewhq00
H19fg5dEaFeTnYxzciINbyg+aVFPWG5rVCe+7STqyNy05P3K1RAYxFdWWrKy3L3l
fNqKQhrO4a54PU8iNFjMupi9aLVL64452HNKEPCz+xo9i3wpQBhwTmNVdk22hkFJ
X/HBEC3nH2ht7uyKQRleh5tXlNVomtpRgZU/LX6FwAXha6JuLV+mzu0t0pz5hMTc
2SARnHhA3Eg5rXqkZ3jQbs2mgg/LmjNbrONiVQ4NJIahF7PAc3HzBpyNkPbE7BR+
tkCMltskYOynQVQA/TMsnKH4DQEe5Xkb8+P6CXLFcBsfbHLB0v01nwv7YFaF33Qj
gR6TUE9W5cnMNxh+50UNiWlZnaC4AbOSDLoQuYT4CKfR8f9D0Oelz90W76cR6rvD
qp0zNGUXQ5CAtj//MhTBd2ayPlLYVCpV7O27LF73/oA5mgMmKnDiFpHtBvJSCoJ8
pKimCrn+VjrBFWSJB4WRB0MjjErfQSrqAryRvXzK5wh1Y7NEhrULI4Ka28PJhZsH
XRL0XFgHxO78ZVmWPo3rBGTU2FpuLPL37BoPeO0YuFNGNXEbWtTpTsV8hzAMHWUl
Fyi2O6ZFy1cmzkqSXRtmT7pW4EKa0T2u9/J0FqahZ8EcKrNGVfzkzBWocYwdaMiY
p41TWNS6fBWUbNaeZrmpfLWFFv7C0R4P3s0sQLkiPqRv8wJsTZksmaJnteL5SSSF
8uVwGicNSYfYg0FIiWx9+mbdeumseQecPV+Mg8ohmkpqGzoJOzvFZBDlOdmDsYz9
wnXrwDDhYhsnRH6hrbqyXr0Rckg+xrKEUHax+byrUcygc4VkN8fHYejDLvKi15ZN
FAAp4JGzFNM3ZiuG9RxEQ1Nmw5FDuicxmO3z8AW4BVvizCsjAnKMW5CPdT969408
xCRliuI6gxsjCkFgudCNDJDq3mLeqEWAV39iQ48HuoKrRnHc4B0tU7fEiJzIrWMw
JkP0Al1x+iqsF6AaKRcS8KTt3uJr939u65BO1/UeJexh4vuoobB5B/SXf1dgc3CC
ukjjIC1WWQdUVgmkzjHsU9Y7KYV6hju25nKE9vKhEGwUiZeRYepzrRbHl3qj+Ov/
YX4WiLTW7zEzMSd9JE/RCY0lOI4NvS5/YhupesA2basGCpR58WuTF9zcdtTqEVNn
Lvbp3BackpDNBbUg0V2qBqE3fvWT4CcwSOFrCM+jA+jpDnRLSTNO90NcI9HKG12v
2ob+PZEJNU26RuCuIwi27duYfvGY2Zl+1t6laBcZbC70r7hrG8jJgquo9rTYCRMp
ySVb6cMSJwwGrB/I1XAqe1gpALL5OTAvCgTL8iRqRt0SItBN9g4mFU1rEK05zU9N
UXvDNT3XJerz7Q8dIx0e2OwVeyypXTY5YecSlzE+ygZCpyGug5nmYJG5u8p5J7rt
Ep8MRNYl17omAgYo6eUS0ontbymTcsOtzeC0m8j2jqIg0PiQjXBQ5y/jbTxTDCTp
eOLaS/3nhsbXkyG533RzUrAsUyFIfv8xLPrhFMQQgQ/1smuEDzdqKKub+3M03pQ0
y2GVS7RBOH5Xu4E2r3BsoueNVQlfFxkB4nDJ5aW4Lqz8AmcxEsZbb3R3uKnhjxsa
p5MsF7VZtjLoTzRX/VKZGVng4NJuXXeaio2R3TXpJcMeoXzZVuAYmSR5eII/QLH/
XzStzgRT+gyWWiPTozoc8yd39cN2ZJKgI6xDb0KbPkicsTmTI83e/X4LWq4OgncR
7t45JpUrgYP4b8wy8JFZRl0BBKE6HIJHzhL6cd3e8zm7PNGtiQeLugj6GwtBUk9C
5faQ/+AYH/vg/ugV1iy8WImCarizCUX8IQy/irFJ4Dq5jx1aJheXcgj6hmpr52uc
IJkP6gX2F0FxAMe8GasryPDZ7Gn469yKhWyDsHpTKvkT1s1aI96XcHwg0tak1evL
ntA3fGacoaQwPAQnzJDDqkxvfK8egQynItz4teFhdjx2qSsIsxu000ZE4I3ssr6F
Je/vz+mBnad/uvsQJxiEQKL6VSQCJxWcqRNVQBr5CqK7p6zOa1ilabhLgsQjLWiy
mI+YUsEisftxLycKifFJ1r1aZ987wFP1eTlhqwn2eDWcyDAn7mPGjirrhds8MZe6
AMMe6a43TyMG/1D61wiEu/W0hdJaV4x4ZxVznthC6I5xS4qgviVphxBekQlLSoTw
8/8QKy1EuQxEGUI7Txm7eHy4cjYBPLaqpYicy5m5uFBSOvDRLcwU/VhskqeKDJ63
xkWWw+vvWPzECfge+xTuIu4y+jiD97RXr2jZWCBTDPwals5luWvYpqYqKur9CQdT
9Cd6zx4lU6kY3g1j5k7GzTuCyyddZIK8x6RePK/ilOj6rpyg5y5N4wH3iHXi8Uqa
4hhwUVMtYBKzcg3eQ0jg2fLzYHu9C0bvcGWCqVahkgtlkP+D7fQ/4Ee7yK2aQwqX
jfDDhkLp9I8bV9UlKZiVdOXn0utUoDBHkh5N+OlVXaK9mkjyGfDQjVUdNiYdCFCy
db5z1x5lWfHRkT5iH84NQm2Jgh4GjhRZ/0C/J6e+ZPFX/o40fNwnjDw+vK3bgqaq
rv+4mZN4ltX2qe1sxkUOhDfd9/hKZcHPfcEQCDYFIM5rjMHt62SCqD9nOs04J5YY
CFDzB9kYZFPu40HFHho8cFYEmM7IJh98ACC0+ZkU1wLdpmH5VFcWPEGXP8UL0DMX
PGaQnPaRsgGlSSP9vXpfy1rqMW50yUpgZRO23MlO21Ud1NwwPO6szgU8wIriOOOr
yv7lftwD2GO2UecD1R4KOi8lUoJKIR/8T1fHHfyXy9bbeOQy09g/bj4UMHUceaP1
avp8ms+HbXvUEvt1ZvsGuj42JMT++icT9U3U3e3n7/Jwc9I7/nJ3bp9gu/CKhIlC
4ciSF0tckjl7qzg0HCP5XsFvpJzlowxA3IF4aArOdUPN2I3fUaXztbN/9UnPsRMT
XtmhS0TYSEoPfgFHiiD6CaHtnff/JKsZtwiTB1htZ8j4+76AmSD4AmhCa0tt4NIp
WdapEQ/srd5JXX+hl+J/888nftRvq4XG+Wse+wmGhTD1nEhlCildTOY9LqdzBt32
2FGG9sIc8hPW448pHG66g6HFiS6ivMFtCjC/hQXucgys7nH0p+XgyVGxfNZKia3V
k7V0Z9Bg+pmDMFwbzpyC5QpG13G6PNqBfFqsrUf3wuYLyhpgaIvPfkHKCJPHxxT5
pDvI+z0Mkz029QTp6CObxfCJXXl4Kb3/KIkkG7hVsBbusFyk1A2+zUc9764AafhV
q6gQ0YDhptSTt+k9Em6lUJFEU1h0YjZR6EM3Kx1L2SMakkalIK/FKkn8d4V/AH/U
Nl4yN4AIs0CISj2cTIGMN+JASMAPgjOrNAwvrtKEJijTEF8T1mwKasM9SAWD4xmN
65C3YIie7kKJvWfy2TZAB7UoCPIQ0DglBP7qSh8zpdvVXNGTIL4zigkpGqbvjQxr
sHldE6aSZf1bB6o5Sgf5jPoltRapgKfNvz+SKwY/gfWJGUzO/jdehDnCIFCdEoib
TGlCrR5z748D8kS+31gsDZKMB6bekF4sxJtPChcGb1yzKnza/6VM7pU35B3Dyk9z
uRse7x0sO0nyvJhlYa/kmI6H6iQTJWRb0Y6l6GkeMkkKn24xi2fcXlWVCFeU3CqH
V+9GvLex5fvXIKD8O2aOl2+pOa512ibiAKYtRQ6dumIRwzBmds2aDIdM4RJ2Stf+
nU75aEJiUbZmVr4ISnBg6jzOHA28tsNlZDad/ftUBPbBOovmiP5ZmVFiV4CmZEyX
gvXD/grySKYlaHnVv63znq0rZKeU4WwjWWWcmX/Y8MnFIjxk194KKZjE1rfrzTpF
cvN6eqj6ogzFc+MLPGb0oGlktbJPgZdU5yhILk5lAz89TVRtLvz1vu5UIf9eWfa+
WYc2CzJUVQ/Zk+JXsaxfbjmuOyugF1NQ0Y20ZlE14HTJFEnjcNMGOJZsLS8Pl16S
n0k+3c3ZiNcay+kgPH+CjPfPExaIqzgtW2yBbdVjci7y901lTqFAxhLCIez8Q7W5
nWyUldLgQ75/uFu2wFwhHxAw5FrRH0EcrQqaSNUkHzX6taadtewxcbMx9YUV6++w
VWUqiRvNBHrfEi1iD/jyage6xo/h7sG4LyEtIbuj2Px1/VmT+JkCUDwxLqyh56u3
xIm3ZvW38rr20lYa4THJ1R/ngXIlffOdSuWenEzkJPDxae4/vHLcdpuzDxHpVKKl
tt04Yxy8kf1M3foNyMT4As46OoRj0pB7A+OuW+0p9i05J2L+VH0+ZgkNDvsaZ1ew
WgFSzZQwC/jVzKPP+FsGC3TRPti1PTBHIPgbgQfFFkzc8VOijBETgJdV+SsO6+nS
DttvZ72K0BSkZYrjPGVx2nh3rAzIAzW+YEaCHifoeNoGq4VynDmf3Xkmc1pSGUny
PCw4lfuzSPQbcwK3CIOjtoE0uGWG/mfMLAnvKrH/DjWABm2fyiq9iYILxSYnq8zF
w15yD3WRCYJzs46lhBHAOyZIaywtG3EsoTbQkFhj5E3vqFoA7R649CncJI5DvEE9
/3EpzdetR0YV+iKnBHBXWnqiMJjQlZQcf9BG2u7yk6Bg9pNLnnMLYab/6817qlSp
37fQFu7zAUWoxKPZiIyowR1dXz05bieWn2xijAE+p0NtApNzj5g+nuN3XOSu4Bui
W77XSpat/Ht3gPd0RUr4lnEwtt9tmiQF3TWPTkTXAnNeQrHGjITBrLQBZ7wayfFc
Kfg5L7R4vikN0mmh+m+U8+Nnw1bh1G7zgaW1xzUyfqCv4v0EBAJEMrRNS+wbw6+Z
CjHGT+cWek1GcpojksHfJ6hjvjCYiPKjuPnIseaZNjsffS33oEZvjlTeIkOBM/Mg
+RlFoVK7FL7oSnqu9vmr49LDC+0Q/zEk3BVDL+bpVgzIcjF6WMFgklF8YizWweSi
9B9Zq4L7gFExSVyzeeE0UNKFl2J0aEUncQGp8wInjQeNsrF3LriCDe8dm67GeGmH
t+1/kxQl3L01AlTKadgefuT8ZHLjg7Zi6zBlE+h6eWtCmTp1ejfvwD5FjPcwTOu+
Pxx1RN3UosJ1ewfHiYIeNQ593JMPtwcaz97UekiaLrqAoYjHiKJDDx49eGj2znZT
fffL+FSLap3icsaXMkxLto+ln6fJ+SIXFCfSUYV49BTecyoiBZxZQ266wQZBHK2H
lLqvk7duqCcRiVN5GAhwWP+2xve7BfMwThR+mKs+6AVAJ7YDXlY5dMh/AdN4rzYz
TrndXzCP6t2DCy967uKEH2x0xIjCYIcV1YRw6eGML/i3D3BEAXSB2fg6YfXzWS66
KMAxpHBuNRVdmz3HPSgPb6eOgW6PNPWg02nPiCXAx+dpwb4GJrFCm5kHAnoWTVkR
qpYj90Z+KONDhcR9VubNjdak3sr91WnaOPs/06IA8aKQQtvaxbHl1iI6PG2fuMZK
wHuOB1m071XSiKn227V0Tly2MvRSlD/gkKV+AHr9GiKCFYbRIrdlCkQxkqRhq1Nc
p8XXoGuaUWT6EbHTTM2A7NjykS0Ov4NuTP0OzSoRb7e1R2BbytbswFYIYd4IDrAd
Jh8XjCTTUycJqhzOUc2GVW5WgXK4FG9giJXm5wE51kGiK4kyS0KNmWsAquBfCeI+
EpofqJzruFBDgAXvv3qj21+WgMt0qdK5Xrb0QQfldIEifZDJq6bZ80ahVSZrAVgS
6KfPxg5IoTbb2fVjk51VaoV2n0eDidHItJgA7Slt8HI6HOEzwPhcuVnmqAmfXgzz
7h6PE1JMsMyXtgC1K5jS/HhI2yd+qNMsFhz2nZz9GX+Dn/3CbUe7Zmlu80EXn9s2
GyypdohWW5oo8VLgeNBw3bs2No3mVJqW1YKF3VlOYD3snZcEhpyc3/ofCip7mhks
YFSlGSUw54eJNkUmG0YR27o1Z85erUh1drnIZXuQRW5XRoF5EVfG+kSHcKmdoM+0
pK5Y39ODYPBcAjwTRPnPzBP+vACZP7ayna9DM06bqpAlJLz2qdLdkqxxaOdJ5ie9
q7By7ZZFOxy9KZ0PuUWvqc8ITqfcnfYLFZnysosxYaSREvzPCoxw7jFzje+b0mUO
E96lwFuKqCiJZT2Rz2Kyrm/X7rrujYHrl/SvTH6sqzpqn0Bv6QEFuT4JHKE4MMoH
1fAoh63I2iPOQo+J1aVJywZbQJZ5jcoPxy9w2/b7H5CSoaP+CsokGNeSWtMkkRxR
qgr6ap24FuOEdlJ7LUuN+zmpMRlaO1FvXa9KPKQdAdIB5KU3cMEPoQiHWaVS/9Ko
QoBdLeHHnfqrQUlVfMCvpB2MNA2nR+1k51OmrKQJrczcm2Jbwbohr0up0DLCHZJd
kw2T4P/U1YMTCjEMC7hx1DcEWOlwWwMzqISb77Gj8tLp4t42fqXm+0Tx6vL/rSZ4
Ra4quks9qxXAkLtu4+uKWx0i3SSklhaGowIhMH48PANXHpi/SDrYhbVJLv4RTpoA
FIke3IyHdf3ncDN+7j2+vc12h1ykBmXcu2chv6CWNWfCTfl5ybgw2S+nWBsSvTOJ
PT361jywVaKhnouXhiv/1wS0PeuHiTjvqVSY/7r0rhfeMOyMgU5rX3CQ8MbrIZJC
DMWVNFQoN1F9ojmJiuMna1J3VPvLunVOtVbHrdYDy6X8a5Ir1QDGlJu/ocz7evLy
hKHhoMoodZrulwdVM+xlQb0tuKJd2t/WKul15vMg7D4n7KizHaWwaKzPQH74ER8S
BZtFCkIq4qat4gxzCI5jeYGdwsW+zahJYnXU9DvDmP6prUg75NMNPK0GYOqQXhSI
VmsWbFymXTLKToHhIGq31vEVAsydnniql8m7B+Sj/gkdH+4pf2lUQvDvGPa0YJav
Shvgu7jS2szKVrqIRDFM0LWqO0BDi0+K1aDoDrltNu6PEiDrAzkmCx998UOCP7km
IPMiIoeLqhA7V+YEtjNykinDKSXsAlhpHXhqOCLt5raijemF9bNsyqzO52janqgm
0AyghKBTckCtWuu6SYn96N45Eu93YGmN8t24Iv/jGdD/JFzD6C6nryWLpfX+orVo
Cj863VjmVU5UisWDdLO09x7avAxKOqWfjfdtYsUGaph9EgrQzVv8my10eZ0ouNdh
vClGUYPeaarB2Wxa5hm6KeJrLJGuWidl+3VSAacf8O4uejeEEbxzR9SGzdQwBIbd
rFXYqiWyK0TINI87sORfFlpDaiQ//jc3w+hpxs+y6dWN2PkDvPfEj5ql+FbUhYuW
OYw0vD8Lja43HLFGut3k+veO8Gjmu8dfxyuY50cE8yQ7ocddDZbfQLCwGdFrXuIb
+tLwGSKy3YVXWjXf5mrS8hsBKi5Ua9Ma1W0vfq7HYdYymvUnWL0QZgUT9W9UW779
faltNoLgy/1cP2sXS1lca5Gn9V3olWiQvIPvOmXgDmaI+yCo7xYq8wDkbJmybm/l
axPjtHbDcRb9xwX3NsJklx7y+BMpPCWFkn+8SDPqbJhQexlsuo8NUm7zisaz8Xsz
X5hairmxYG9px0x9GrKddE1u4EaD9vxLKk9i+t7b0oqBG4j3Uu3VWxjcOVXyqw+A
Smu3onlXCFGNEHg3ex8bK/CKsGkJVCGqDCC4k7Ya+0C82fVkTI9Cm1+22Bd0ILEE
iVL9tZQ7cAVJw4FrVMt62sogeYgE/zqW16bTTFoMxV/jEwGtKawlztxAxD/seGVy
IgupeSKLBZHo1F9kKoM/pztJQsBSbQgPYP5KOHP+LSiB1G0Q0fhglMx8UR3ak2ah
7PoVSN46akwYOJ/xgWqAVhRtXmGs0wcJxNrUhpXPIjbDT3tJbABdUw9Ms13ouep8
mRXA5ypcQE1iGqfR1Y6uE8MG4iUGLtK9VwPw0m+X7RHFB3Li87/J/minjLJXP/mr
vL+Vkl8Q52SP7nIda2DBZNJOcitcQ1h6IriM8G48QBJEGDeB/e+dYGEV77esf3v4
gfzOpkQ0dBbFzekNgrNXlqpRnOdDcj53uIp0xbdv7/+yOZNH/duuBzfpPvt8aNWz
OdOTFDRKsSz8BOJFgnqXvUsU+dxyqDcSNdumABb+RSqLBvU67oIGy9OYCzvPIxPk
aB/Vg/EYcxH3QgHTL7mB34fTtafCSabdvFqEhM5qNKGl+1NHcPWR/TTPY1+VZPKG
pqZmr/oeYZusLq2b1uesD0mMSicwZHUm6raOXCzLYGUXJ/7WAJPz86VYlzOgvwLO
gvbR3S6TFl+vd6VTzd/QCldwQ4t7KtZ/VJHjWtu2mtNZ+md+7ClklqNexC9cGbKw
hqDiyT0hXWIpLgzyWfZfwZ1mHBeKMtpNJQz7uJEybEhmFkxFsQwFmcmPgc5rMWrb
yfcbQfNNqwRKxmraL3vW2I9srA6T7+68G3fNxLOmd8/+3HaqS3/vZq+qZy889oxk
+beBqQQm7gkKPqbIeDHpOPU9YXqdQ0+td/GQSiJNa9zBYlUxbTKJZLuBmPEjobOe
dpoPBxZ81ieSzaXM5CDxk2NmtcbWmwVrRmQOguCmqjDOhDg1a7q5j5DhVsR7qjlm
Ui5+pDojhSKjN1EFIdkA/SL37KMzhxlmatnGQsB9RoIaF9BVvgdYGic7ssU3mZbK
Yn3ZuBvRtLAfurJao6043SyhthAL+MxjsAfwbc5oESBWOz/3JjOekYtC828HzqCJ
ZI1amK4ZPok6PRrZwmNZH3R2OKZ8UuB6xomMXBd6fD5UqLnGu5Hnds/th3daasUm
b1b2QirrkkvD0obq0LwzIsUX0PzuODt+H9eto0KLbvkc3fmMcgRYgFBycqf+XFrt
i7jNtuu/Ctf+nmjLW11I5hA78VfJPuE1i863OdLLm35UyE0qEQqetygNQH1vx/fy
MrKJprRT6TsCFJSRWBGH5DljIaFUEEXNTQNLO+HEyAi3XPGYBBJ+g01NZn/dc5gk
fzhrJ/++xHNs/J+Bqj3w9abqvZZGo6DHApWfc+hN9/kFM/3M1VHQKArOd+V0gn9Y
bVr6BnvZ9mDCmQH5MWeIW9u4dse+t5449TmAaL2fLONtroQ59XhA53SDpR6zSzyN
M704VVtJRYkE61vSmNxkmVWpbGxWWFAZQksruH7LnDTaoUGKEVeKvk6ATbnsq9fe
56wWcxNuystR1aRHNQR8QQpVIq+6emf+quKN53iHpXlLjwhbRMOciywmNug6DLVL
CISfCxA/WYA+pr3RWypmaxwMFNzImYYyB/VQ8kWGhQ8YYm3kK9vRSj4Ce5Y9rzUp
FEsIJrnMfZW0co5qB5LmQbjlia23u73wKGxPM/FsNDmWDhPIUfJvF8AsJJ3QVvPT
J3MBs+Vr1tVLjUDn9Y/U9KF90iAzQ3YUYpqGsbzjmS5PowlcKZMQO8NxeZFbz0Iw
cGzInAVxKvMc30DeoXQCNyP2Yt+9FN0gosBlqKZb7YtEKCK54JP6J4Bcz8fPLHIp
bpA4T5oCB21zMHeBgq3i0ynZoEksE3Gv82WiU4BIb4QKHudqu2eIDh7k5oxJiPFa
m6jurbpT4MwkIaf4bvJO9eb9eTVfSnxESCLibc8gbIkZcUNkQfW1JUp0PPaWO2qj
H5S3S0sYOBCGOXG5tyCmaZ/JRijkBauhD60IJVmtX6MQsxW4IzMqrzvLFucxZ/+f
kLaLSU9TGvgCkPQcRyAunCkPx1/caWv6xCPA2IH5H795BUec4neGelkgF46WCDuM
pDQe3Nok2F/GoOefu6lyuyRjiE+4Raqt5DDocyqJ0vWsDO0+NFeL5SsgugI/Mwmj
6/nGeBPQrSiSVFvZmQ66C4aCTNbT/sc3uox9w8zM6Zfcg6XNuktSYyGmtCXSF8vN
/PrfOsE1e2jE+24Fal/hic8L3N2AdfR9fyjYf8Gx1RutSdIg9b0wwX0OMYiUjNAa
n3jJVKIGvG3DlhTTAYqz78PsPXE1q4Ehj058uKaFeSmdjlJikO5PyVoBmjosU2Td
5VOlunmFchTQ24/6jfymy6+ZOQk7wnUOGnlDSNKgZjfY51Usk2u8N7vQ8P0gms4v
gWjJ157jAZX+i3hDV3o7PHmQvNZkyypuM+Wy3laImYJ3HLUqyI0E0Qvoqv60YtqT
xN67ll2GMMFuLxVu8izQkH3QMO116PplBRAbIrRIvV0PwmSvpu2v323/AQWgslaw
wOnVNPPjX7iNQhdnW0uuT0R4GRiDZGkYTExOastixojHEYwWanX9N6t7SZUYpJvR
Xy4LIIMBYkJ0o6qijV8/+5d2Y/K6J8KdWMQfNpGUhOG78bsVuZ6y2MRd/RuiNAYI
v1ufp328Mr84XNIDps/p2TzzpPPGND4AKHj6mq2LnHQWBbjEFJ5fxY7ycMHjRW+q
eiJd32g+Zq+nuhipv5Xpad+MIetPQJqEubPpaDUiq3HJU6R6W3tnIRdsHa4VDgCg
+hDojahMY8doAnZ9e9ZLeB5YtqkgRagIN69KD/NkEnTAnaFkzmjvyjfxV563SPCy
d/CxB666XNc/G7p0s82rusvcXI8DyGZat8YhwYLZkHj/GntR2ZuP3yj2Nlh+wvpi
haIR+Ppl6s06RqZndIqRUnxb49SN3tfr3TvIduDlHyijY09VE0oUJ1Em05fvlPVE
MlEPXubdNoPRORWGGE4pnAWLPWlPbw2LdrGLR72vjbkpAFtwlBdb040TUuR2egKy
NslZJ29/QBweIawHx4w/gyt7CNpfa+sSkVb6reSvQTU+if0iJckHUuZgA14MGYhf
nN0AQt4R32iJM/90TQB+Q2D4SxTAdlqWvYJ1aQ/n030N8xiw6nukfWgpaCCqpNjD
Vn9PM0Rq3Q3I1CIpR60BzbSsM6Wtn8ajoQRVLXA2dY8DolV6ToR9rHOwExYwA04u
K4mJlVJUfkg7MJNJKaf8a+FWn7eJdJ1vfmQVo8TBj0HVRwFkHZFMkoEjZHhkPm+3
zPS7eSWFQYIjbSSHtR6H9J7Ll4g9X9A4jJuiSxZT128ZjzZe4kKvSkl2yZqK+9Ga
wVoDJN51Tq9/spD38BdxbAH/TDWiCgkGoV/qqsTnOAuMC+QR3F20SOuSutiG9jkI
sYsd5qGERkbEUJRW93lKYEkruHfNWM730OtqytIz97TEPg3oLv1S1IEwLLG4QmPF
mW0octO8WEH8s3fh59kFvq1TGVebpopBU5yQpT/x0N8pXMpHc1c3lvFY/aXsAkzb
44tPYiCVKhQsskHpb22Mi18K1O+cMrESqlwq1pDOqoeOVlD4fmXSsTcXRfvCrOep
fje1tqTvRr8NKJYBtf63ZJNxX/bdgv+be8qU7hMeWsHPXgynwtC3k3DQlXol8Zgs
+yQrwPtDQdlgLe8NbU9LkuS+CMM2HLIcPIL6s0grweBtKvG/0bLrN7HzWjLHlB3e
xPDbEn4ol2V5+yymKe0UKW+p6lPBPjylrpQ0iaum0th4FwlJQv0+WlQ9hRx+NVxx
29J0Blanhb2tKSrPJFt3m9L4fRozaXQor9e+HaqY6rYEUWnwnNn53P4WEzULuM7R
tqNfk+WkBzvZjdckpy+UymUkYsvOmdLcy4exu1ePJi67K/qfEpx3lsYMkJOo7eU2
MtsR98lQekHzbxAInNcSInsLFWgmn5Utdzi1iMiSKXtO4/386Bjutg9A1eFLlxXm
ArydrE0+6R3blTRs+mcJ2UEl1cjA9VF+w9enpEPN1X0gkr5K0x1sTRfPcNZ3Jnyk
aeAPyoYGaJZXvmwFM7k1trjME2l4W90/hH1sB5Byb8pFSaqos3G7qe/a9DpUJ2YG
ceD7njoEmmxF5mTC8EhSDdUwMcs7OBTTn5i1qzPU7n+n9Hh1hE7vxA+VZ5HMzz6v
CG4JhjgK0Jk6fQhtTxjzFtteweDc6v1vJJXflANddgutx21toWI7jE4a88Zgn9ET
N37cvRQ+CWYVOrE5qrpUTU4g5nHoGbfTBWlIku/XarspNb+sgkV61jrvTYaIxoIs
ZOEx3FbFlrUYJhfS9cMenZfMSATRoRnibYWTOIkaz6wlxKKURVtC+fm92o4BIwvD
FMqXs8ZfRbBvP6+AuAjvd/4SCNsK5mYpZWQzY8E7zcpp8KxjHyCwvawvCiLeHCVq
hp6PtfQH9OA8t8huATnEiamWr1/P5ybQt4g/QxR724XneTyOmqayvB8V9N0ARq+I
Y06QJyDKgl0rZI0FEuR0pxfW8yXlw2QgdCo0OBzVKL9+ra7exWlWc5C0546QSJUu
ZF5j5tvue12E72LSlJwxgbvt91iVSCh8LoCOO+Wu20Zobl8hOopjhDsnlVPGQXL4
ekWt2cqqPtl440FiDimPEYKlb9sXNYV41c0jOt2Z6T+d4CvVV39GR7nL9LSVQreu
WCj17FOR2FV7Jl/DAnkkHC5zRl0mTpysfKFTswwOx3eUSZB/oFOTXVDWiaicwRBi
PTPKfdDPfyJnjbz6vU27hjVGTje+1bs1pjZtz7R49LQ71ufUGPT3322uMaI4PT0c
t+/OUymWK7308l2apOZNLWkgvUVjRSlJpl9rNUafCXsIQnMu3lMdhIb6vOjo4IRO
6pJ5uKjh/CFpGX6Z7CM0yjLLCeIGuYl8+pMMLDvkng7xWAHxACi13Xz+VjODLIU9
50lKoFoBbqTQl7RBe+3e7NKnzeMMtxRaujNTNDWnSftUk9Ns76K09AJS7MxgfJXO
0PxLCcbqG6onaPb2uatA5F87yQYFVtoy9ciD57r+iFn5gOOyBPXrttIUPQXtcBvQ
BsqVhrP5gOx727qmif+xjPxu25C5SD1odZNlu0Tg0oKkNrI9wyijBqzuNPlsSg5M
toUS1QJiI0IlipqdPVsn2ISguhr48lbmNtkaq+WoM3uOTKelGugYHNQGZe40WqDg
bVEIaXfJl2vHo5QuuhbG33MsAC1l1ifDqmPwf7J0yoxtceeUSlHfl98cX5y6nI8h
Dzi22mcIB3DPcG+OOlbn7lbHG74oabtsdAJg2zQBbnquYusp7KEEpzoUcY/Nej4n
gqDZzjMYL8CnZmL7itTH5+H/7O2Dc1x0+uDKRgD8jYJpe2x9IHd5/pcc53IbOLxE
2QAdnCI3vYHMAm9YYQabF6gdY95x3MXyfHbzHuKJjZnqP8PB0bAQBY4rM00+i+T6
9iA1RgtR7kyVroZwQ9OYtTgjmuWYZijlv5+JJ+WwTZpIR7DCUOCuiQ515bVcaGKD
pVkWMn93zA0dCFmy5bnvmTje1oyGebqmL69O5vW9TlDGq1EopLqpuR7RV3FUX21s
GX6tA+4Qqky0F4So8o0TnJu9AWoXGduOGEyfa1Gg2fArZSvJ/ynZR2jd2EctzNIO
AOfmuKg4H/BCMeAD+sNLgfZzXiLPnJw9eHix9nx+6ikeE8BSc554VFym17keABI1
VuDQ5423mOfg4kpo5MtJ6qaSJIZCZsg1QoHjGcAfS2J3O0fLg/lqYYzuXYadAhUC
pnyTsQCisTrGo2T86lwRIXrebmhW1cCZYlQrc/lgqkiOpwrtXlj5Ljff8buTY2vH
EKyBmR7eX/v9c5QfcXcJvS695KZJ00HAcd+oRfYDZHNGRRITbbjzAofqGHHTCeAC
LKBY3gAWz8hETbkwg/zxpIvIqjfEhmZePToLYKJmce/wDGwJa1h+VOFlAV1g/ba2
B5Isr7QGx6xqV8SkVNhyFur1QSwZwV3NHjV4AbTmMWpNzIVSl25oCSHdg3Cqi4hH
YlBPc79+iwCzcQDyaNv/umAGmH5cVf1eUTivC5RxQtoX3bs1w4NnoxBoBW9Hc3AC
PvnqXzC1cUYk46D0nW8d0uKnCEEuL31FWOGhsPb7EFWaBQK94jGYj8iZpgEzRkBb
X7AGdPi23r8HPxNMJpst0dzu/Acw0xU7+nIKKxCgiUc3GWR71aybONMwyl1pUfyy
opIc+ephPSc+/6botEAhxOtbWf47ZmvciaQntD8xs+GZmChRYp6AbK28xtMF3/iw
o5k3A2Vu3IeaDJierzwmHmipA1H3tiCO2M0xMK9VX87+LU+ClxOL4rAUvQoqQLSs
9EIWi9aEIt6c8w4oAleTqcJNW+l5IqZXIbDBit78P9euwZLumSnOXffQk5ES3eKA
svS7GfKmcuVVeg8PQ72JaJv/pjLm/Pbl/wak22FxNbqeUaBhBa0O1obZX/UPdEyb
rEodyjRjojDx0McScXbnTPwmI5Rnba6iE7M0kyFPZMTjPk1bpj8L4gEbq04VS4Le
Z/n6w3V7dMPIRWuCQGFR2iq6qEIvoEQAJjQLiq2f90fEOcXS3lhLRMfuZm36dTsz
s0gb/vjlCB1un0J3GboDw8Zm1XV0qXBlxhv9l1p7jPauwRt8dtfajQl+bwA9rQdK
UYqCi+HKbkDUUmOZO3BI691SPzaTKAomDvHaLa7b7ClYNECPrvBaJTatZcjXpKqj
MpdnhWg/6DsbV1RcdlFPFrim7HOSDEyzyr8+FWNq1ORhX6LhEhzkoYeFCP/8Cfxn
8mTsi2BNX/n10pA2lxp66JO/WdWD5XPF3xGWfeQ/mSGH1xXPMSh8CKdLaqIInUoL
MZaZJEYVAIj2AYCvpOMu4FwhVC9srOy77ApHqrXKJOBXnA9D+iV8lz8MYGPr/zCL
A5d2H50Asw+tp6+OzGY0AhIaVN6ZbFdmYJlE3Y6mXbv5hZlfXH0uB0+w0Wbrr9pS
ltN7/dssVz+ATkKf6AdYFod0xs6T6laW3khL2ku42cZBrH9I8trIfkbn33pcG/fW
/yHMC2SjK82HM7UFyGdLi7xpHc1eBMZiFiIziuMADessgGYm5BphH0muzXC/WGeH
07JSyRQXXUxIRO39orF6/EQumbG40u+i2WmKNcJqXeidlcYybO+iaONeZyHg3fc/
TcDbjcEnHVTJ2x5k0JrXXq2Cyuwy9XcVpiSF79/B9l4BzbprdMZPmuj8dz+vZ1BV
smGxrS/hY5BNd2pwKLGzFOhj/6fhW60RhuHh1nzziaWoLYBS8+KI6n5sMS4JwQHm
Bv82TlNoHZtfINisLo/aU18nCBqCoysaj97FLcf29YCw9hq/w3gVtH+p7swMvYrj
yqi/vc4IWNqia9K/kpzf0AdfLW+7nIZ6ggswjE3iIGO3kaaYr2JJNjhMKZLYkXNV
KqLv1hnu0Dw5tPGHLFpsUws9ijlSHhMTXQYncOLUkdYfNGN5zL3QGgUZ021ux6F6
96DyGYxIerA2p2tAMTAoG+tS0vc01D/dIo/Omgc3aPOxq/HQezqAHJiEmSbT4XAQ
onux6YBtQZcjN5nSlGC+sJ+81j2bMAdcOyowahFhbSon+S8YWYNg0ZQC+4KCKkrt
z6qDEzI9tjP52BX7UFhj3v8/P+KzcFjezDlokESHWYe4oNLPvVy96VfJmS0l1fZb
X7a70NZF1/vkbvrbVkFGJIj0321VeeMEZ6rFW2bA4kC45RfodH6c1Hoi/RpJP28L
BiBXN656JLwtGuSizU1UsxMP6LDocne4gUC+24VwN3OmE6DPG3ApQxTN6IunBZsP
5CijxfjtaX2XgRRTAIqXhxle+TdUvPHQuMsNkVKpVzJEe105MEzNwOYQR5AWJRnF
ON5TKzeMpgRlsCROkrKM1gtJ8HL846i68uDYSHHmburGy9FTYxxmaKMihztN2xLv
WIyMP2l3xbUJaw5bRQEGM5XHWovz79HUAxbxVu7DMLv4Yxcu+cNldmRl8Z8k9soG
hwKp/VUiOCEXdFpixIA7H8Njnbz8WwR338oLe/Um3xP0OVq/oa+9UPP1i+nKT913
Ix66V2Q9gU/SkVrBeOjZcvAYbeeyFqZnasd4FT0y02FN2DNoGU+raZn+sE3pAZpz
BVmrQXBkYLmcMiihkTMRERYDhq0yMpTjiu+3bEBZNqrCQKz3OFYwglPBvc5xr2Do
nsZ6MVkicwbLSvopur03BXMRNDEL0tbpOh4WbPOnMGALVc81YADVGu3l/JaqqovE
aim9lxmjUf7IGBguIiY/o8U6qUH+uYvFeiwdv4eH3f0YiMpWeGs68A1Ax01BQg28
Xr+dFn7/4o9NkmwIRDKxOL4/FKul2R4K3snBv4PMPTQt6IYzUUxHHsIiUEg7QIJO
PyNjUBe1/h/y1xHfwpfWMwOhQ2NUljuuv9mXCJXIStlMFJFXpL3Wo/L+ERywalom
aLFXgCU5T+ZWN6LUsfjxjrPM8FwCNEr+xijVyyAyHoMJumLnbuGJykoiLzcBVFRn
W3tnXeRjooPgLTRsu1SbDb9ow2Mr6I7OZfVlILHoz5Vw53UNdj52tSQ3ASjLbOm3
ydld/3Y5Y0LYIvjc5y/utu6iro/3z2X+4tvvMXc8o4Lpv77wpn5v2z7AQrIXPtzg
C7sygsKk2xdeIARS6W67xNyJ5UZ/T5WZWH+ydnFAVeSmUuw+oDQamt3MyZtm8JxE
uEZsZryuSY1X9Yd042rcePzonmc+r4WozldF6zMrOGj2ECQMFAJrtzFdiIwWHFXU
QYnd+tBb1QuKCFvCZb+lrwNS48D5t6XcVUvrKCoVxXtEZgKUKRptJ9LZEFkKkD2c
aiUX5juu4GGk9xKfbJU+8kLlcnayRM1mrfs2nXDTa2HIrvmn0nqOiDcJmSIIMreu
qN269nTbc8wulnIAP7mpQuwzgvJPF+kQj7FIF+xuSkfZyFsaGnMZW5S56TINChes
9lt2/3UTecK9o9NVq/qUe25piW2JunLHRiyYNxD9EDfxYcAg22nO53Ul+ONA+yBs
JLcJTSLDGo3WsrdNOBKoE4C7ely5jRRdl8+TYdb/WVAL4c/0LDXBMFjr8JcHr3U6
yAi9X1AfngDbipDo5IM6PS5k+BOHdEX93SXoxxKcn99X3nLikW2V804HtoI94Txv
KNbpRd8f7d40lIWIDHaUhANrZUg6Al3WHLeDQ/OyAXEenJ5t7FWsqNmvjtLLOZD/
U23FVKSqpEV0XGJySmbO48ehaOALyJnXKWxGdLYWyz9SUSMXRxyLdORj5yg134XM
lzYchAUiHOZe3rb7tfbuTCwyvS7u+EQ7rh0Rlhiju0GmvoVhdbH500qLWCGF8M3/
YQhbB067jFO+zpQu8l2ABOVmz2JVybfJvPwhMaEqptuY+QsO7ckWtTyPZL1B89aW
rPcIfoLJTbXDZVUu0d4OdTZnbKbxsQMIM4gMizV0Qz7lG3N0SKE9I+lqthoyMxQl
TOhNlUqJNviaynao1+H7a6IWQJ0ueCYpmY9s3CCnU5jxMurtrH9MGMWooGomo0pc
l0iik5X42M5Gc/0RbKRTJMTmUPKmxAZKLD5W7+jFuIoo4TGrC4WCw2iYaixCWhs/
EJ+4HWl0HCtTh6PSdwbvyyEzQc5zvOmo1Ec9o6SrYBCUCqW3HIWu8qCJq1FuTpXz
fhzdobYjZyThEUS/uq3KO63lX9pkAUnxwjIOYEYXbyzr+L695qoa6am+5XvxFhAJ
0324aYiFwlk/rMi5F5gEkz3fmTXKsh7I9gKmH3mMqYJu58G6h3XVGaTCWQoZ8q9n
bofKUT39yGY9wzDDjibmlojE3ul4jOwzLA/6/JmWW2iNr908EWr1cHNWRaseiUps
/Pzkm8QkFLuWaE7hAAG9sjgLQrj/jXMLKdc6QFWqxwXXORsoteDPsZ/azPo/oalj
I86qWeTOBdmh3P6TbXosg/aVCwprSmfHu3g9eAKC6Z0P3NYqzIlvhDkw7RqF9dZi
wmybuotB1+xH3ClkTwgIGnQYVf4Xxk6mFCWjDV+nACNaSBIPYz7E/ACVaOmul1H8
LNo/hAFqQKob+2AhAOp9NTX0krahzojocLq1P/BnwCFVOBSz0jpgLZgnWLIoEeBA
bjIBdIGm5vbpHL4bzM3jXFUhGsHlZfOIoZUctwwIzgAycOQsHd2yvv6gX/fwasqY
Tg+zfl70SIrw7vN2BfO+M2QazgEOCgVbRGXGZtM0ilpWLoDnOhxMgyRWRx8r9wK/
eYDek6J9k4H8kNDSXuO47TmtgI0CBqXZC+nxbvypq/PGAotuY74dbzLxFj8R2aEy
Z2c9JNr+gKxqWTm/DUVbHNclbZnfidvh/dzp5waA2H1ADjPHpAjppyYJ0RUsNsdF
oQ+W9YsIkmwBiV74DVctS1rOIzdjnV9H6HS6mIfssDmVndKp6ABX5VL0ktJ6d+a/
Nhr/08cLS0nN8/3SwJ7u2LufqXlaEg25iGHsBnvucNxCu6aQPU13I9Z9MKDV1nOn
WOEPGBjD3Vsf+eWwluWpRR8AXBuPiXZRA0qbRtbRWZViODgIViFC671MIImSVUax
sh18kI1O/fponcRxDG8ES0GxLA0b4XvhCpTiji949JwxP/oZsaAQitSgSCXMqUQQ
TuxmvchEFoF+SSZy5zODdzDA+QUkghGLFbsWXpPA2EvPFpvJ13jNXYyl9IgR60F+
jDiY8l8Icm/AGhUFR47dNrhw9EI7rivEBgbkoz90MvwJc450ykacswvnYTS3tFw5
/3S5bhCALJWUwMhlFijGE3Su6kT4bpPpKilXekV90DvXerCDBkNQNk/esRiHpVB0
29+1Biuo8X8xCy6PYPCvMriBvsgwvfTpXkvuYgGZZnnRDsgXleXzk66rdR3beptg
W7yCshWirpEAi6Mxir36FvCrsVWK0g8T9ClHMdBHmRepET8KvQaWbAfPSIyTcoSi
xCG59xc9H5rFLY0Bahi5kD9TPjEmaEwAfQBGkNIzfXrv9W9iI8UF7HZCbpmJxYrE
kLX2l7lSm7EwEVOybWBXcHMOLG4DX0Yyz8caxZBhwUqqabEEqTRbO4pzQ29lwIZB
pr5g+GGTcZTdnLzhJ5lRnD18wTmX+Cyb4AX4Y8jFScNJBiKXsLe/tyLlhIldtGgC
FWqZFduXc04aU4lb9NC2w5XRUoBlWJw0cH/736ICJhvlty9V//YTY8KAedPAdvsR
nYZ04KvTzJfJb2h6KZjLOPEdTKScW34gr4YU84fr1G7sqqR1C2adzs8adiYgK84L
vZ9LQANSmNMp6WPqFSP6ZplE9zv7e9S+cAIl3zGvfEO8P/LF6J+zGD+MknGql4je
84lypSc1oxqwpweZUQ9/Op2KihNbkW7+YhUPqAlLFybicxR4TeVc4xsUjxx4FFq2
7mMEuIYWesyAsuhwFwzczDXVFxD4igN7fvNtxljBn8EoEeeWvRLnPIJaEJin8Ylr
scnwM9C3i+yduX4C5PXdBAqK4dyZ3X0SrgrOeDhe2rkUEYE3y+jDKz83EFi4DPKo
Qql4DSJRv9xskv+A01rMyC/kh2zwDTd6wYcjEZxVmh5f1skQZXZiac3dbCYdEwin
BUI4DSE2fxdfkUbhUD+zK3mcrp8Co0K9U3TOa5mX+opoEkxc80N4qM+VD1EryAhQ
oaho5QfOt0VDqEnIFUxcjJIBEgXcG0mR+ZM+dX1IXGQCkckZAxPRyIVqYm16XNNo
mcMdW0VXpqfYn3njoLOAtoeTmH5i5OWvAHQm3AHo54rhD1MekG9+431VlZfjWjCF
GhTutrxN01libl+gMGmuHwbo/e0dFpKgHfSOiqLwixkQGPoTmuhG6zwlLVbQW449
G4UcfOwDhqe2XL3EAUHxUH08Qr5UKOAAO3kJSLMG+n/2nb9j2F5eXVnn5xupZKFh
lF/JoDaeAOd1rk2aniRwbMjX6U25/msccZx3KTmVRfiwGp5z8KVcjGuwiQ2+gQx9
xCHnOUofhnOTXH9d8Uj0w3mxY6MAKmLJJjodIgC2Wbz0+mNvaUWjPBBEQWqrV4J1
NuEY3OxLgnQzmVdUo+6XS3rVcwQGDIqQGui6WGhnglHLxz56WRfRLXCULFP9OH7q
aL9Nv7Z0px8srGUg2TggihdRQ+43Rha9vTZsU8RO4jiOCnwenHYLwj//MPL0u0Ss
8ih6BRpOKhXQsMKc/tqylaRC4UJLuidA8Sr8tUvIigSusKLJgXjBT3ryrQ4/Yo5i
g/cQX9sFEUSX5mtfCIu9bpsLDzH0mun06BSJ2Wulq0snUbk5zLe/YhPR6+o0gmEc
SqyaDo0SDyCfBN36gi3OBJy7fTxVJ8m9KJTDF/7t0lcECPFt8YnN79GowjpLoaDC
M2jaHdjKW3zkicgds3X/LDsFNpVlJWamQCocVfq7Xoe7oy92HN27pxK4PQGP28es
XAelDsTdV5oxs52Z2DkVSDUCeBkrPcgBeKysMqw2VKg0fNlK4kD8zP1drW59Dewu
jOWo1zAcb/cgsks5kSl1zSc//5eS5Uxa7OatGB4dF2bwysPeyIpoV9lQFfxsp6+h
++WbGx8PHpwwQSEpeLMwYDF0wiy3twlV09mR020bnmddu4E11D0frfnlg+DjYYoc
R1bFkgqJuzGcn4gEqJDlenvWVqzng8fHIJAx+aJ5AOcumghjxVARMDCrUamZN3CE
9aKT/pGjJMt/VF1HnL3aZWNaTUWf3fJAol4HnpXueovGRYHitzTClthYSX6fpm51
Lfuu6goOvjybS38FJpqQ2Lbn/6VJNpU78riKEyYnGG0JyaOVpani2r+nI4/EWaZG
CQPbRg6O79n+gX+QA48uGj6HmPO12+fiLPeNKvMxibr8TuR5pvrrAebmyvYV37H+
M9pV1FZU+3vj1VF6/BaMgGAG+VrpT3NWwpa8W+8aajnHJaj1PCFT+UNujOUsivTk
mosSqnL/3WXF5vS0fLG5YIJQ6OyyD/DY/Vvw72cvWbWwmzi5JheCi23D5a71PR3o
+z4lVZsC63mOdxgYKs0WTCTqNhkrVfcY9JC+Y6bNLojjlwQNLiYCgal21o+DqXgH
sA3A+BIWdL3GurQXiDTHC1j3pR4VUKlrXkCzHLvFb0dyrMFZsy7ouRrCZGyaF5YE
EW8xe0jLUodUjIS0qEXOYVQ3lWfsnfD1icXE3Lb/AqJ9NkzlhRXzHsX9u1FySG+u
Az51g4wrzvuS8f4N4ThNBpyzMUxNJCPfrpjGcfotYhhpgnt3eDLao0XV7wZLGGij
k6x9vzmsoPqVZ9uFIp0qwL4UzCn9merJGS3ia8IqS9B+eY+jkpXBHGOHkWTXrc4p
ME3zOqm1s9SY6V1FHq6B8hbmlfcN8WZfabap04G3PRNHdCm21/rwTOIRHtfxiNoU
PARTCj4Oj8RSzIjQ5Dl1GIM9pPGL0V9bmGpyFt9WgCNWn4nlH4u+UyiDqv5K1Gna
9UaY4KIjsvj93exuK5sz7qB8M8iDxA63DvoNijZN0ohAYgQgwyo3AVID1/xBwQdx
u2vj1JumPV28n4wreBdBvwhItA0rlO8+gACRWcaEp5TeVJTetIG33kaC/cbBz9st
EobxVb3DWtGC6ES9EEFgvovbZG0m3WG22Co3JoWuptYAyTCtku0EWqpB4PeVh68U
KKUdUMq/KxzDlCnvzF8hc4er/jkz1shwVat3SqeV+s5veTVU1te+LSVJD2FYz+EQ
DrWhqyllCm4bKa62JDkCfxDUt/scN0w+7S0vTSWF1f7ocNlqNmFBhaSg6g17J5jY
SjMcAfX12blGCKrnQTaEPV1GJNfpzBAhZdNeCPvgnlbbpmN0tgXFNE6o/HALVTR5
UJrpztPlAukEkhdxpKAC3uwZ4Flj4RdY41lV2n8EFLpb4KHO4kUYLzhwI/4H/cPw
FahFodJ8cNnsaN53A/Lu1JSubCk2Qv6+zqmvC/8cukEeswBPmEanVm1y9DhAhv3H
b4JbJSMN5lnWAneFh3rVE9djnPWltHHWQZEaqwa7kqr1ZJ8oG8X0oiirx0K14To4
6SI839lOGTUbNWT8NB7OhdH8tfAAPvR/K7N2U6cJrCqjbdBsWCLwMURLBxr08Cgv
fYmB2TcDaomsJp0OBTxDJyaw8takOboFLQSb6qET7UclmiJh2As4sbCdoawOqoH/
0g4BdcH5y37dhdHS2hEN1i8nHe6spMqK5Evn9jZPNx0s+iycbk+zXEVb5VgIiGRu
ls+QpEC282DYs3DlLmOvSiLlsFU1VGIu2On2FOphfkh5gI8fqEUA95KwvDpW5j2o
B7pzY+w8qoEgdePqVsnDsbpzZnb2AGyl12RPFOVXwe4rlQ+VU7/kHPeb/dxkb5n1
Gq5J8xY3554tMfr3119Or85Jq7WYab3IMwH61vIKL1PHe4tiUSZiN5ImeHuM5eHf
daldDr8f56Z49owBZ4c19kIiyTHtTAkDZa6cBT0f8kvSiaEK9Qes2Qmqq1P8z88b
/Wxl6qE9BY8H0a1IdYYo5jvMEWisaHopFIC2OMWFbaeknVkHvdMPWNW4I19lYHeM
QR1YmIoMMI8EqS7GTr47yD8ihPflX6+QdGr6Q88mbjLehD4Pe9oz+BY7uV0bmuWI
RWvKVU+tMtxQwuS2UV2r/9Tczrx0XxAfcy5d1kgDkuy7CE6P0JQYaAzhNkVrwC//
m1cufvFFs5u6si2bkqdFbEgdmeQCKgNCrFrgXgnx/DNzdhbRe1h5MfuEZtqkk+Mz
PzQv56qFj3iAlW1DUDSpwwUzzvD/xW2nG8CQhW3645z+ot5q8w0janvh4icLZa2u
2j9GLCwfwBWRgdnGGChNcghpYsgzepvkFjD9gKe68GoPSBtJ6qMzW/e9FJEdy6u9
LdjTVMFMFimmQoAmRCEax5fVque0aS7wznEYif2zVoAAHPAb5YkyL7e6BqJiBxYq
2rXgFKsLdZz/LShJgYbtohMlpLA2jBolxRpERTmo7JGPkaNoQqbrwM0l47QCPn5L
cBc7h2NioltNNWqVI0f8Jcx6FVIrDIVL14O2vCICfv5T8EEetb2GFlEex30vdU74
SO6CPwL4ALMpaNpdhR0GHLfr60M0L+llK3brt+9+76hM0TY1XxRfVTyi7pCVvxLR
emaYDZKlHq3gCTvWW1/qYwSiuez5QYTWvxN0EqDQpdGFwKI+q5o7iKfSKUof2oNa
3X7Z9pI9E3/S6IxjqWCpMaBz449FlRF7V95sPfU7mq3ea+Oe2y3CJNNtAY8cjQeO
Tx74NL3JWgBhpKp4YBsuYdYwA5LgTBX+0inmKIUjKnh4i64w/Pl2hfey/DF4UgHX
hm3ysCNnqTeQQMhPYv0hCxNGaTwJFZ7VAF64nWLA1kPhzlB/kdxyutocG1MOgGk/
V6ka6mfRDyhuRFosBBUmB6ET70XCSur2EcrMSlzybjkdat8+KhyX8x4DaqvEa/lN
YcX0R4SKHBoL5rrDTML8pBC5rwMbR9KbXq2Kqn6OLGley29BBLsV21mDnbQZYT7x
4piZXEquj2/EJqGwqh1xE/l/nwqJWaghxXPgdSFjJYqViMKcQd5rNeT41eJGnu5T
K9d02M9Ef6u9jTGvFAv6T7UYl4KCSpfc8dvAhgH/S9dn8Wp4MBO9HxjVIhO1UhEO
2YX1Cj+XQUQFasfew1ImxGTKiJI8gDKBvVD/90jQG763pNY+OJwGN4GN7fzA2Ge5
7VXuVwdzd9HYRS36osUXKEA4YtMIh2a9w0ne06bTZWxTbo5tLUbIvxIwUURYBF6u
kTUv5ecVU9APZ2t76YvkDSUjbtQ43oJYjPw69xyb9amYDAXvQthnl1kcq3weR8IQ
IgFFg36jWi/Zu5vIUGsiXxLRKwGOYhhXQAvXpIMBCtUvcn5HI6cVSgiJFmcQsQIh
01fvd/KuiEiuzyuuHMcinWmmZKZRzuWQg/S+2VFWVRbuMgnfWHp8es1mis7XqdF8
hecb+AfCWD21f8dZQTFmjo0n19R65vtqLzQJQwz+aeX8In2iWZww99piLu3JnT9q
i/bCNYSo+e/n/AQjb8TJmb1303YeBpCKjF31CkaPhjNs8Ne8HEoYddENZ4zlH1qv
L/G49S+6orfUk+/6qcGqe8SWtR6So79yMsG7sI+L0KcojdCR93wqLiFQwki5krGX
MCCW2LlEse9/CAXArHGf7BksXhZElrLysLv9PzFSRiiGZTVoxFAskI4/RNCWkagS
gMEyTz3HyQjT26UcS/80IRuE72wt1iW1FxOzRZajRMYdzNZOFajKebsv1FVhSRZ6
uK56vrY+1HjXMzxU3QExaV5Z/mDmKH/whuKRiqa121pCrRxZaWx7xt4HC6E+nRKB
JjOcaQY5Bg7shAVOQlMhx4HvW2beXlJLOVwBiPyjb7SsXsx05p0kIqV+jFRdaSUj
hjUN6MEhPMVy4+UXL44pk1Kmh/e61ISQfYE8se3rd1sLEbI9zYxR+YFhxn90estT
T3wiih9NAAxP3yKJQAT/bapb/azUFh54/VNpMdoSikW227Om6zJcRwFU/SSTXy9o
9DkPYSvREZFLwzGs++wDtWHrsH9pB/kDrucICTE33GjfX5aqZNxsec1n0FQsiOdi
PEHOzKAUAMBr8ts7S1lDYasLSmDQl2Isikf/4oY37qO7A3IsUrL7uLzXTkbu88np
XdWYwhnJQ1tP5dOF5BCnUdv4ssr4hYe4QC4VPQw5zeHegvir/rJ3qwyaA/m/zPn1
CI4BsmokGuxa1RLRgj4sTRQqw24ltKDHoopTSBG8MFZbcvhxLusgFAp9XUaAypPR
vWjsGfXtzQW+aNIeUHPuDHCY8wVdxktvlw9OIxPswlpUOktXJkpUlpyUXg/kK0xr
DxWHEApGFJ0MdVM96SxDaLrt7CkiEXM8IguegH2Ig42R6tMe3CO8okl3eEGqbXNS
i+lyFUalLTkGWaVdtashQiXXqMlpn8NBMZ5yBKKOKD6p45WE7wbnW06L4P5MOPVI
K8D8Cv4hQ/rvtAG0q2+UfiJcKTe+6RudpmI4vQe+KjMjvK0SAhxYH24IeCxDMzzU
q+L5lTTSrn5KjiUg5kDng4k0l/kH3Y+3mq03U5XLHj9yjIwZRqYxF8ggTsOOHp6B
7FGsUKZRp7Dv+TsSD1ItD6YuvNDZA5fXWQIPeVJC1xAIe3XHtq8aTTchRslRp2hh
fljB/u9XR0liZrU1DV+eir4VNNdyGbkcEIuZ1kUcsWd/LAOJPVcZL/xoUmTIJi+L
ykkOHKBRtM7SE3wmKRF/mW9KHx8ezufENIzw9m6k6KXjGQwBj95ZuepXuzWVTxBO
l2pnIYE81j5NWMZmx4lArxzJC22y7yXRyR9gDRtoYQ0fKx73Tw9xCk7/yCqSsnfT
wIYXWks1Z23z2oX2q9jvpVw8Xcpb5MJVTNb5+5VP2GZUo1LAjIXeokRLdgM7pWaj
XF/75payrnlXsvbde3+i7OnKF2bmfo1S2sz9wbF0PNy4gbpAHcMd3VL72tUXxVz4
uzpUpsVn/jJQDKkFJz9PX02G0tLoh4HqJNvK/GbH6fn+JMKjwO5e3/FhV6eE3FIW
6o5BHBwPSD2gnhiMoVUCFKdXCNeey1FW7FREHzNF0ANCpr/tXYpHZD0ovbMy0mjM
gLsIEF0zaAOI/Qxfeq9hftuXJ4b8e8qRc1LaVOUJUOSpCLqOviyoX+F4SeNHuIAu
nOaflHBbp7yg3RMb4UVRUW0cTms1W7HGKQZRvV8mfPkg1OOFRb5kumXM6NOwUNp6
GcKnJiXW0XHuP0w5zB0iGycmRKDdlCdkG2Jf5A209Zrat6hiN7OH49yvdu0g4/Fw
BM0hpnR7EDXqpt6kqyksw4/bPclNm55yysuLpueK1AvnOd/401nOxVVc3onwZ8UX
RAKW62p6F+IZ8l5dZ+sCdc7KoccID7DdM6zU6OdtGLFY+WqS5NyNywA5D3Tb/+Uj
Op5baD5ViJj5fA4p3iLQfshrWL4NJjQ+3vRSNqNeoMS3/9wYeY/NjdhkDX6uIDjp
nakeiLDcyKjoMGzxUitkYIBacYBz8BGGPjIXh3HsEH49Q5fEwdLWLDsmxM0KZppY
QbGlITCHvBQKiJmFPnjiGhVGA/R2YdHhLs5EBgMqOU58R7cNZ02IR1lwp/D4InhV
m4qyc/hYPmonqynq7K/3Vb5TRtE0GWnIZMfK942MDc0EzaxLk4Xj2UkbFIxVtzEs
9c3dXR2DEk1cEWuuOGwE8qqlA6pYgQP5Nu6E+88siIpaZ7IoP3an1Hf8AUkk+Pgz
WktubQxig6HlZYwrTBC2/4ePNjjBL4V173txYsoCI34+y3hPqd/c/nM8B0mAaYi1
tfTR+hXmazBL0+3xuIRtOBSUfPmV0hCB1CewEwXXDDTW2wgGNrQHL4eicIkI76IK
kBr2sq6xwRV68IQFL8s0XH+DfC1mDUXmfwtV0MNmkqZo2Pd+/QvnMfEiBJsIS+bC
BSErgFLSgzQVTy7G2BfOqKMc2FzNsOGnK2FCci9w211a+P5Q+dQWrZz6wPVSWsmm
JxX3Zcz7n8ybEdq0D/eFKf8RCSj+usrPm0UJvYvKgj7vnx2vKzyV2lcyyFMMwYfh
XzbgW+Wr+Sgwokl/6rUvaVm8vOlQTuyJMsyEMYb+q3DlcejPSdfptWRgb/eQ2hxd
2f3xwQSaraEmv1MLHjtDPZLzWVAIDtoDtYd5K/iY8bS02TCVqfwFjl6z9lJVVToe
xK9BtUI2GSRY+8j8lk7mg9N3VBcS+XkHxUtGE6f3a2wubsrsaXQqtwgGYl87kFKq
/60Oz8kUOtzF1Jc6dkLpi4Ij75SX91mngt8OnfkVoW988Cwsz/mgyMkA/CsApYJa
TvRqKep50u54oqFAlA8fafWpQUht9kMdKQRJPaKmwMu6z1J5cqLzMpkO8LQmYxmJ
/8LYUBCBv9iTK89bBCo8Ori/M0AyEFxQnjj2Tuhq4kgNC0xt7dwiBD5uuu3TjFmK
0k48IH512G/GFDykEoI9N6pmRPQVl2XwZ2P/s8m2XStPl16WZResq6Y1Cv10ZC0Y
ijyUxc6EVnAsttvYlIhInlJgao7Wa2vHj2uCaH7beLmKXHAbZmCj+d9VdG12Uf6y
AXcagHizN4nuNMBnDiemvpi7nlDmpayYziRox5w0MX1E3jY6bfidRO9PcAlQp05q
lwFsNn1ifKt0rV7f+O84TUmxH6/lFwpex0d8ddnyIyPZcFSoe5wbtrxYtjW4qpdd
iXDNPvAcOoGnaOq3ngVnEXqbYIWqyRCRsypwaBnkFdSB+Ujz647u3oWzK4aPQ2lK
cTzKOBbqE4eleFxf/4HCV5v6fX8KIPHmh04eQe0VC6aR6k7gfeJ+nnPBsEeL0mYZ
mg+OBnzBZNEB+gf0j6xsb4D2aM0ba3ZVxsllgYzEnqT71m/puBehyrLycZ7TJ/cd
PZtTYaQTKLK2ME/4Cn7A5gmd3r+FZZchb6NOw3gZcnski6OWvQOa43n7fownk8rk
5jldHnibrfglNjwDku3uB205mOKPL8JNvoJxzgf30OgfurVXbjtzRW0ZK3MP2jVt
5mmaTM/emZAA6NwMZzM5H1NCWmgFlNSi6+E6Yg0A9gpu4MB7U1s4r/H/l8WtSZs+
Sv0jRtdlot8a1+VMJmvI7EL5j1TF96SEa9DJuSm+wsqCECF1TH44iXnWwC1NAUmz
M9jrGOOkRGGE6BXezqsZ31MzbxcP2Zqd/GogFEeS9d28wDmDTUVSMpCFLFFqqBjG
qSFvTwGKp0Z3B5JEaBSf6TQunqkoAsUNuNu5RibdGE6F3AbCSOMsxulSa1+y0y7d
b3Kc4JA4G4mWa6y1THlZdbsx12H2DxcYZOnuMAZw42gA5eHU8kQgQRlZfWofQu13
metVHWOZsSp/HLR+VJzxJ2VppzxAAN5cYFIx3OJzHKxn9tcAdasC0tMBL7pmAAFR
4L9ywaCD5V4qKaHMc3zKgDsAXfluMQo15OwhpY4sPHKJecL6R1GFzHVHD2cQSOiO
VbJVmYGatGMBeOZa3vOkuZGVe17ctlbeEPymQ7DeKjDLDb08twagrCXChJLDP53U
ctSBpAE8u3zTf6pz5yy7PDXDaszwAW9wkU1GoZrWHVnytXeyeoxoajhA7SP1HkmQ
CdUh+9eGAK5eue5HxvAsQKRZT6o/DsiTKNS/dTkxMRkuEsFFyHXDf7bbj9kNgIZJ
nbIgZQ61bR3CwmhFk+YJ7SiCv6NAOLST/C6vQpBcVYbclaj8D7v4YR/jJFiZcfDa
1BP+YxLKOrxA+Ue5yh24Xb8u1Qsk6u6Mby6TNBb92QYV11PA5o5p+zZ99/ErueYP
UdgK+lRhldHWhPARYOWkaq7tGC/s/jZgIbbB46GwmxuwC+IELLLsgnJ7FKCeGSq/
8F5lvX3YJ1a0T04EoqmWO4kIcibuV9YbIScjJRMjYFSqMTV3+BmKaS+JMBM1s50E
K/oM+CwjG7t8xpzEQi5Zxq5EyU9ZrYPRy8efToTwJgXEr1CQi2av9+8/VOYPc7Pf
/7B5XcwJ9N2RKTnYCW+Uk8OfOZsUSYK0qG0cFXSX3uDgIOIGp3JHrPCrrahQkD+s
0Qx16sh83FfXZMD+eq3MZ1px1Pj0wCxwSMmlv/Ey82bpZLfasfsjcDvF/4GRZjLD
IzFp8An7/TQ9ZCpbkzzQzG6eQ/i28w4keOQVuhlEGhRfXCB/AZAFEDYXqbZqscv+
VXQnX0PAVlWR72vmox9IhviDnbv1q7h4n9dhbrQEVdafisHnUb7P77KyaOecxp9x
xFv4Dp9Ob7remTk76pMd65huj+SzOS1wP8r8BdUVyh6Sq2vwDGpZz70hPRF7qmnp
ui6haMLgvzPIlphbfK03+ADmsx9ppGFIDzgpN1/TWOc29dQGpZSmleOaBA7MCG0f
2JAuPlQg5EeLhbxBxgE9ZV7xX20QEB6MC7V235Gvqn9jzToniqxtBPJCofeMiSnt
rWjIuX0F9jRrvR0kEvqNpwE9KsiZhVAPyA6yUZ7VCkS/Q8a2YurqBTzeJWX5Coj5
gm8hJHHss9KJDIXwkTCrWYsUStwV8z+dYg1js6yIpcLA5s24KnV4HQPBgwp3bXI8
MDPTsOcx5S9wr0iEZ9BvhygyePaDLxX+bx4ONsLTFpgSfKOQP0P+xxjiIxgW1bvG
Ai91lEZVg2D4QUHDY16+LffDsv3kJhHt7dNy+q40DBx0rxhrxfT5pBYwldNijL5m
5Pp+fsY4z/T26mvGgNWQu97aXNx4P6dV/+/WsO3FnLE8rMXNkVowD2asUfX16nbW
2Zi0AIx/dQ/4vM7Ya3flCZeDiUY759YvMpOF2BqRsVYxJRVZ79ZjaqFeqCL6ijCa
njjwlPKCTray8wVHtF+d9/O92gg2nmFrewCVDDk2rXqCAjDD8Btn4RT2RDdUDL2V
M+4kDIM5uTCdLUwqICaqw2/0+hQFVpve4PL9gLn5BhCxhf+fwDcfsZhWQ1Yx0fO+
RGMObzu+dQMpiKEZOPFF3lD0FLBObTeyvWjIiGR5My5QSlZbMUgCMRgprKC1PypY
QxuEtKvWgMBH+0+lS+XTVc0TNHwvDLuHe1HaAgTQyFgtsFHTHhIMkkeZXrWkvytA
dbv1Jdd5/zJ9nLLwJWNT9R7Mu2DL7IS/+LHzoIcY7BuaQctP0tNxMXzS6yNyc2XK
pQp3zKmRh2o5cpG+2RDo2jULem84HikCfo0qSBSQw6onF8YT5RIOuA/p5n+to6s9
DfvaxqC5rG57/vMw36QFc5RJzRC8L/7qPaPRk07mvsRvh2Dkx8sNkEARwjULOBKm
avZPbHW6U7TP5TkFsm+lrN8kLCn07ub4GvRBwrcnWg1vhhfapBuaW5jr0ty8F4jN
g/myuC+h9opuV8xKR3Y5aYXDgLym/l3xxPavPPIM1trepx6aaY6hrgMj9SmmpFoK
oo3SvycuvAFeg0ZkbvfrlucNlXIgYBbosznCeUGFeODvG1c7ggFp7TxlAIyEVax3
CuLuTBlYcNoiQHRScG9daYxz/Rj3bn6WnPZNF2TpAVatvJUNSG5Zlsp/XPhFUASo
GNjxl08KbiCeJNKPYxxCIaEyi6HnRxk/D1EN4tIzAhX6APe7l3cDg4rC8uWggFfB
mhiNpJ5vC1WpV9cDMDFIKlh4+DQSH71CC4K49pqKEBllqVvWT+DMYa47tVnVIuzV
pJxFuRequgbafzv6IwW02kE4xSdcx0AztImPRlb+vbz53SxQZp8PCRT/b2kJfOlb
Yjpr3csLUvXYf8Q4KZ1IOIujg1/zhZc2PoCnJZzQWh1dfvyV2CgSdA8beVepV5R+
0Q7fCqwaJW/R/fvWm/QFcpiP3CnUUJcRhlm9Aklt7qWTSH+LIef86/j8XIZL9nak
pUXSFsIZxXE3eSH4vLQQkgaRu9Ha+S9qB/h9ew1J2LVdD0o0OGy2n6pJ25o/Zuc/
14dzlkcQMRPcuXOelY2Rj59XTzszs0SQ5sE6p6dDGCT7Ag5pb0cVBpaXpc6Nnu1g
q7XF2acGHyNDmtisagD1NQPK5Z0xktgvSAHThVATphXCGN/kSm3+maYL1kO8bpt+
brARMHUj/BGcsoyinD4ahloDO5owAkpFDuRCbA3X4ppJKj8hmcWS5yclVqbPG3aG
7JWJ6nO38V2CvomXAXa/AS3DCWhepvsAWJKYhJCYOOatDH/SxXRLXxB1pXBtSWW6
8Et0YAyp98HD/qBuM+Iz5rGLQl/ENKrMXs9MIpvM2RiwtbCgYQiUHpu5MrtmYPdu
Yd65yVnCUKxWciIQ/sn8F3jGQqMhuVhm98TNmRBBZMCDdJCWh1xZeoXTFQYze4Q6
vdCebEgbgiew+EHtkIAGx53FldSn4KysqxVt7Kx1CsP7jRlxAUNy+BOZoYuapzVz
Qp8h9FMktDkn7+1ef2jOd2LbD/JjcxBGlIx4NrbqJaZ/zq4EYcyjgcyE6NlCXMoK
X1IU1RUDUR2YbZcw3yIpLITdeL4LnR1b+69qqbxWOrwb2FgNfTUISCYU0MW/2dAe
c8PP+6M3Kw8EbgiuzdEySok/f8ghSU4f5e5NlmLDJUonQMIBoCdVe1jKE7t8H1cZ
39MUBJaQ4iIDfX0kznZ8juLNxQd4Y40j5S58GJiDU8JS80H1TZj0NBMmVous5aWB
Jvvnj4cyt6jV217gO8IznsJ9V8IFY5ZmLVTfsmdxj2gKZlGTX/O6KD1s28VJrwbD
dvh+xXhWm70jQZFn6wxwblKilmWC74xu60cU1hr8FtEVX1m/WAJujY6Y5MnFkYaf
LZa2DfE8KWakgT8hkv/AtYLR0zfWcreRAQLa4ztEVZpB8tSWhFqoTTEz3xAACveI
QMMGN8gJRae4R1M6NJJRlDY7Z3t0Mx2qM5vEr5i2wOYsR/MKNI4uH63OhB3i1+j5
4fysbVNAv62cpH8rD649Ft1W41IV0GfffNRGEZep8OpITE7AVdmJH8IL/2tgUmCF
eRCYgeNB1e2aU2a0KbGFlXE6v/VIpUiWvJ6GLUPD33O933y8cvNBo6CpX1ZMquDm
7DSYvXGjPAQVeuq/PVtKw+w1BcQX30fYsgi/6PfpCO9dCau8TdHrwdOhXBfqS1/2
1zODh1XzKLtrJx/buWwRzjF9TMJaVIX1/4h0cYjPCJWVR7HGQ971soDugl3+PD7S
QzbzPQwzTgFfNOFebE4+8s/6GNwWJCN5gpf1pWoCwQdb8x3za/qJbVHHSbCpLaj+
mVOxv8KcVuvr3yuFz346MK3DeUEmn1wMw4W9hSKtkyQFlt93O8EZ0ArZmB+RD/zq
/FyAFkv7/iMEaTeDmWYKymo/gg2yTdGYS1DbyvrAAzO9Ox8LV0sYwZYDVlW2HWcU
YbZ5oVW1UwXZ9wShZV5WtvED7YmwM9pM3Bb0WMCKrp7+HT4lSL4kxWHFT/faQxCS
iDCKrZmFD4isCCOHM9gSg7+esNlZc+VFd1UZpo+ogu3y9Qx5St3bU7JoTZQ4bA+O
9l6XFMNUefM6O9GcTLZkG/HjS1CceM7qgl945aakdMYWpedOfP+g7KeGbwxGgo0k
3L/XbY5U+5j6gH8Vt/YBOSD1qIRPfku/+JxFFd9N5bghuRxYXpJ+s6gzIkO0Qy/T
KqG0fsMLR4fI4oh0w/56QP7PYzWm32kdNQ3B1m1hiuBNhecfDCzQGxmfk+Yccs/v
/ArrEDu6x1JVuVJ8uncm2unr5EHYXfp0r0bVbpnj/M6NQKCBNaFxSg6x6NbUCKYY
P/wSpkGQJVmn2m0MSwc/1OerH5dgyuQXvYvSCSXHpnXOA5xyr6ZhAcrWrE3k+iiY
M+QtHjAqo8koEijQ3iatjXZKq9K6Xw27w0B+lMRbiHesuqLXp6XmEKnPQIrE4f5+
Hb1h/+KmS8/dNS+Djr0Plb79ZzwJsUs7g7TRnXo4OI4JmX8Tff3jATyjO9zWyUSs
s9XwTq+LKT87p02hnPenxumhOAN/tItJr/wtBWScYlHYBTjuYpVWTsinQKwkOE+j
V9cUG4q6Jsdv7L5aiNb65bQlsClw7YszXrG4mdwo8w482GK0ttzwjXDvDuSlg/Ya
qib7Ap2gtfPORCoQeDXYRRxScdYPjkEDPPTXZ/nDGrQcgCWbfpZmdd4ix/c/YEjx
nnt84laFZ0LY/97sgdcTo5akWpW813T5eIxcLIBBUggLrZIrEJ5efKtyJ6NH9sur
RLCuIIZzsvf7YrutbBH3KAPhLUo3EO4mUOU3RnWfexRuRpix9jfNnUG/J4J7l0Cd
d8E96S1OwQYkakWCzom2WeCobBEyMkWeY1mBH4S/dGgO0Mcsn+ADzcue9ywusw+c
tC2/jyMmsyb6cSdMDHGCa31E5a9jYgA+Jzn2wseqoImyTGH1hS3px1hIelridnUG
iu1t3nL+8jAXihge6fRU7FwHkK1JeesGopGha5NgnPLGLSMoeNjD6p3PiPUB+lCC
ih+KVyLDwdRvajmnDN2nc7Ef8LMMrk52g696pdCFIUXCg5vNXy96B2pm7sVpT9YH
MgMwgyXaPryLRdscrksvXwRPJ9ltkxEdf//GUwAVO2QfyNL2zh/09PgjfX5AEoQR
oRnY25l2xY41JJoRcysfrIavrqggr4JHNRctWUkp25NbVQ15aeXn0bomwG+AF8S9
5tgNoP60azzneueRs9LwBC6tBqhiMASRVUl8bM20DnS2xY3zbsqMRDov3EMwsmVz
nMcaymEc2+U13qJvWADg93u0A7z/UxIOeGKa3Q07kqH01L5azCLnWwhzJfJZ4c1V
1HwWFDIQvCUXEwbrjMu5GPoXWNnUX0Rn2Geinn0XnGhVRr2kk8ap/BUv636cs/QM
eLAoKk51ZFiEEdcu+NEKIxXdfVXCm3XctWz5GS2H6yR3OQQ+1nZTfjdHCjvxNU1C
oFN92SOpR2//Pa1UqmHHX4lL27ZMfD15wixLD2XpaqH4vhzRiqR8fj5fVLvrUidX
8bAEC8eIodOH/fpiXONal8I9zbQuTSnEYRUnWbEm5pSe8z8CTTxHv2MC+7YF07Ly
042g7q12zfUjLLTxVG5NZQ4PFmaM8err8IWgV+LO0+EbE4AvX4K8UUs/ckA4CZbq
+JwgEqbhKgFVtwHyLgYc+ep3o7MTqUEZyh5OfwfdfLAHPWJnryrmt9IOVpFPUuBk
5yJsTfJy9iwmtyEAfTYteL4r0UMpin5qm6FXtSYWH/DOztPRIwmyJxpKjwOaLNPm
r/zvGL6PbJ0CU+wr4wVY3O2M8m9jNiEgJTErj2cGk1Of+jHAtj4ozfifqZ6YzJyL
FkDVDleVl1tDd/VEn+5fVFqrf42PypHdMg9n2B9i7jQdHZRgm7bFe1BRmocYzcTZ
Gb4q3ux79j1cIqYyRSq0kswnUI2AnDhqxrI59ggvjaEkZ9sP+9yHpzrSEuU7t67z
xo/48dVJPLQp5Czdj3JpZ2n8lTn0K8p+Wm4XeFOGwnie0e9D316QBjJhqVrTLmDu
5DtsziRqUxfbeu2th3q05XGiqsHuxODfdKDqgnxCyGDKinkBLH2VSidpNFHY0O2w
Zyig66/ZuEuXw8rEV6gXVM6AugZXqOwdy20wBGZve/awoPJE/g6ZLSJ3IWTF3cRE
fv0DJgMcBgi0z+aZoTcU58kbfdF9ftwCXS85ONEifrYwdpqcdKrV5xXkXBTKaabG
tO6A82zJAR6mK9WRZK7GWy/eKTeruGR5aXw+wZhBta3kNJcw41rOk0kgZEJEZV/h
soe6DBNwNl8n/aRkZICaYEX59lV+Pdu3gQg2cNTAq1CkDUZJdm4UgcH/VfuIFQIQ
ue0LPB9NOvWx29fJ2kmD/+4BftY2d+OE022aHhnqmwuqX9e0grsG5XcgbYBAvNsw
STR+//01mk46GkzV3Jnvlp8ktNkcq+4+JbeGoa7401XbKiBMzKIJZxik0ZzrEg52
UUFJQC7GIt4OKOVz7xRQ9DAjR1Mf+ab1yMAy25QM+ieTALm38af/u8PKA1Kcwjf9
WRXeMOHoD+2yWNZJYK3Jm3N0ZRthbjK65JYTeVbRpojYL/eHHXGfSo3HDHKTURw6
+l5Ijh+y69BGb7vHdMAHZs8DT9DRPNV08jfX3wqdJEpR2jck+I576akqtXrHvpQi
6s1ad1A5BASX474t5TB058iUC2EBctnRU+mMLieDHqH8XMHPx961+CcVk0UkNnEE
VFQokndbwIcQrYyR06tA8Di6iEtAeGH3bGaIDM9hNqLVUke3AadV3RyRkfVrEd8c
f9bYwc/9Si68Dy8sj8LUGKRViveWfIV8AunOpxDYqY4JXP0euv+JtZIVxydasZ/V
y3JUNlhwaNavtO6bH4Z4K6Sfml6mTLGdvsdy9ifWaMhMw/pfFKG+sRpS/K9ilBy7
lwR6egFrbeVrWFgGYwMC3bNqnU2oJMkuBaXhZxqdPtUfqk0g+CQYbaXsulNRw8n2
IcxDf2OdXV6eXtT6GKHPzVguDxbDGF5WGpzza/01inx6yOQ1Ve0dzyjN0QRf+I/p
lBckgoPja4j0Jy9inRZ6Twso5wppF81uUd1vNMngMIiqPT63J5HO6TyDspEbSwTk
rBpdvVJ6rikGNXOaFkfWY8d2JCVgqJPiHOmb7lgEfRF+czgImYl7wVzVKPOpacyo
YbzfDEy88d+1hN/PpQZQ4uvGvSAu/+SdXei4gypHAaRVpWXUeiLJDI8DbSJD0BlT
m4UZyfkiK+jIzO0jd1L/LaA1C4dWpCtGYMuIazriPaZTUZbCbE7zIWFfQy2rMtKF
4zZJeDTOAfufeyCU3VBr6cTvsJrlqPeK6jZA+EheEFsFj642C7LKryWdtMM5T+a+
May2KWfa4pTCwSfb96iLpQxiobDrvR05qgHwp6Pas9XGBfu0NuF+nLknAbOV33AI
tdcVYv6NMOmIPp4G1O/2sSE3kJQpWyYhwym2pje+HDzUh+yQSA/9PXk/ARDFvl+7
+hiyuP36Jj9KM1eIJip18ZCQXktsPdTqkjal9pm+ag8Rq3TOhM828XHjSpDl683A
pqr8I8z6D0JEqDip1bz0Wm8DMduZXIGT/Fki1w+WWwHOEwGdFox/56SkdclXfqEF
rAtmQWYgq50NpDquXu17pEIdas/Qr+8jGEMFMuxlJSpLbbfXJODsdMJstu08A5oZ
7kaf8gdhYWRo8VaVD0N6mTwMsqO5Nf5/Hig5H/PaQpzBDeBtw4p/Z9+Zf00TO/AH
kJdc+XSLsJWtWkk6+gShOZSiQ82nH5gT8r9GPhP5IoOhwKztn08AIMA8nIuQ+QyS
06DWQVwc7t03R3Wb6qyAeHKw77pt96GrWiEG5VTKTplv0jNqh+xDwhXGTNoHjdTW
T2lTb1wMEuUR0CeP1YBbWKxAvH/fL40t4XYMdlS0jj+apiWFpf1AXpWpZhoq2Fzn
rG7wNiNJZbccSxFGnqwEkEsVWLUymCocrzkgnhLmgVFA8aqma+6N6geuve6ZQZHi
yjq/T2tkZy9VHsxenblNito/nivnYOdN8ddKUUYdpHmK6N9D0g24n3jln9Nsqu7H
Puw592mBIYcsXNLOCzdGlIfhLtc9X0qn2jac2bnpAqKeLP163lunW7VwmxZgCMjj
lGjssLyUgSsRar+Rh4SrDtee/FgZ8DdqT7iqhO4BpcfEujQ4IWIMAKnKoywuvpPM
ofKpyNnY6Oj0I1JGqvWgHXDFV4EVZoTGQKjA9TyawcOAZWHRscAc/g/it26UKkye
mRhbQ2XbLIS4Yq0HZl5bSwJ0Uy5c3mWD4wAH6Gxm7TlJpa/VbbvHI8AiD8Osb54f
/3DM2UV+bt0XLMUOLl+rkQS6e8PICrrqYQCjng3l0vSgpruQaHyN2714ft+AwuXN
vPE7SPQ98sEplUNWgp8of4hM4vEdt7Nl3Jo9etjwc1tZihBM2PQ/nR+cCx//ISR4
/nVl2XrbQmsIVzsnz0HpMdKS26agFDM/Xd7qjrryEnzC7hCK4opFR0/2Jb5/8evi
K9y/seoxzTdKbaT+EQPcgtdNyshC/+2Xu9C+dhFUe7trUXImli0CAr5c8qzmVY+O
+l81crH0pgXqq81V29kuqqnvmzk6dD4hGRUEtYYyOdvRI11T7Br/nzqLUg0nlWIy
uNO7Z9N/vxrBIzlIWux8VdvqUvK8jY89WM5BpSjqKl76ixlru2pneclUF1OtoUS/
uYY4QqGMVx1Uu8BYDi7znTSXbJ3HR/BRw7XWpQPwjD3MlJ4jTHSs7+f/nHtzt/gU
XhJJTRtmN4kdN6ePVhZq5C/dAgy2glrC8MOTVIX4s1xy+VdJAb8qt2xsVmosyQcT
gqIXnSYCPFaCixVD9wdKvyDOM7AsDkKo5xjtU2lPE4/VCtbG1skP+bUIng9M4fa5
DhMgn/4zL/NNXJMtj39b2ATB33lz578EFNbMYCwukZvtBv8KVlu879Wu1YTTrsTc
a3JvXhmufqRkjvGeHZWMJwUn/t1e1Q7LWpvfC3qfAiirY9taEwBproYCNxEq6AXm
Vfabf2aNAMqMDnBUdF4LBxtqXasITFYu93QMYJ4lRj9BTAUzGXBSDTDjMlfZ19Uc
sZNjwU10Oe5oTMad7bTErOXsa7w4bktLJRyqxTZpvyOcrxXdHP+y0pfalwDzNX9j
8+BrskonHCdPlWSqL11vjTBlnWeYXx4NixOzIn5toVs89TLHcmH1gq2CxL28vcyK
uQeRwoulzp0r6RN77a+5NQPJ9PbCjNKcFJzNQ5qi/r+kEX/mRkmi0a6ctRqY0b97
Hgw1JFvUowkxiNzbxd0W1RBaRztuniVtfWByxaK0gZXIBQvvYBUj91owVqdWB+8i
unJQOCqYUrH3zahhnU46HCqcH9+vZLMHjvZx+8rGPpg9VV28yO0e7SdhTZQ6fItj
NqgIYb0wYXKS34TBm1YbdexuF16m0UOmAxbP7DwOg4Sw82ySU8q5zZkNOovzDEbS
DNYwIRRZWFaKXw9O3GlCHgNMKGLiSzRrO/CESd+V1WFXmTHe89uXCL9TqUjW9oPB
sKwxIHrnXde5NLMXTkwbRjiAtxtlCz2MWK1tVL3ezLzPXNwNFRH53Na1bn7jJUtY
+HBoW3O/108iCBjKpBA/XZF+O1fgjaAD7vl7YZcz2F+xrJ+exsA0ILCstJhzbBaA
ZKyuwJTEMnyXIf2YlKi2Hou9WoYk8qRA7LTmvOUrI7oYfCB7YzHJHMr+oaiMDfz/
JxTnrSzHEt5N3L8kBnRoq8Pa3E+fGTFDA21pe1Ua/IL/v/Ub2x/zHEJsz7LoBD5Y
Uf14YQB4MUNP9SViDGYQs9qbFHK3hR5N0fvWdXemUjsPl86UFPvp/MFbUlW1dPKM
VQGZpDcOG780bdhKF0RLL7pku3lPH1zEuUjF5QoqwEuLiRCLiVlVdUwyY4tCRYCK
5+By1QFDk1rgd17dt3IEhk7SSM3Gs34f/iSazTqGGISZncENUEh+IH40N9AeqC6Y
M95I71zbDdt6VEol4KhyMMKhcQY07+kc28nWZt5o0afuOxJn7NvB4JZWy2hubFAW
rpbEiqyf7nwJbu+fr8GQrLxHB3qWrCxA5iqJZA/NNna5I7Gju1Qy5M+OvSIiAkD3
e+9bCyNCDXw6Q2lM/nzfmLCeJyKQOmcetyRqBgTsDEeNTd/OuvylCIh2noyV4e9b
uv3qx4Eth22UpcTRvWz2kgIfO9a2BEF6PKsd2LDZrvhMqs2hufD1rX2/ZZujZ4FF
IfoGYlZZsljwqBmjN9phVPPD2WZvbsIPLJ1sdv4PsNRAasWht3RNRvJHzz9WqZue
SKZmwjkWkBXmNgsSeHhekXbkw8UtTR5Vh9EntVH6IM3EaoFIpEDKTTuER/g4/+aQ
qWMu6wA/7uZdMrgLkAawBEwcKPHdVwSGip/8/gLu8IkjvOMuh5jnM0/K1oftEVPm
4YXAcVfWApWpFt3RbRty8AJEm6QzHKDth7BOA2oJXDCHWtikjH1KbWYXO5GsT9PY
8WbmdEpiZDj8Nb59jrjhkV6bd8p7stjVA84dnX1BfU9SA0qQoQV8ihVM0Wzm+twF
aLuQ4T2OhOBE/rN5y/eAnls09pWGW52HYTYjVEgzvSKWF5MsV1DknIw+Yygu2o7e
pPekAVG9p3k6CyF5qUNxAxGlm5mhnd+sXmEAxXZ+JPDWlZuuhMTsYvbHpf0GYM0/
IOx8ZNyy0P0ERfsNwckCpZakVOjqkkj/y5N/HjD992bN4YoguFUX1vN8EjcGBQTt
FVoz75+kIUMSk8oGzl9DODU53dvOezE50/OLMukQJ70m13qlTzTchVCydM4d4aon
+HtgjAnRUtpsmILA4wbo3+NTwDXNdnOi7LzJJqK23JlUzU2NYVUXCgFMhT1vxD3O
00kw12ZRMWz9x96OV9KZePXSoBVDikzlLslWK0i3tx8haEqM9scht+sge1PbIsvH
ka/cvCHofW+NOuJ6glPfZa8IMDpt3vceA/6ZSrz8VY4f8B9pKP1y/bXAcwD4w5zs
A/2+CknS+5R3JMej+AA6CToq/xF63oxAImD1xBLgXAJ2CypiFVbdcDLBnixHeI6v
S1WXSqtGwKym+9WhRZE/KmRpPzg64/Hfg00byh05xJqVqkSIV7qPuejttbTe7MRG
nWOxE1x8y5zeo9ldjRTcOSEroHbGekLQ/LjM9flX+ocwGO4zN4dNskWjyICkwQ6g
TteYARuhCW0DgfY4EZ3rNB+MO3WVQTz2s2xRYdtrh7PoOorj1D4c39PzGaZeTo0r
gPJjYVVcwL22kkujpsHTcPiZMlwIHdN4Sk6KrOpGDB3nWPkYvP1zYdpTAzLu70z/
DOh4vW9MaqzIRMsLSOTGlR7+8gyDkarSzVHiaIaT2HcHuxgEIxGt5ATeDtJWNNZu
gpicU6eOsvxepzKgZNrkMshak7D3M1znJe77X3RvEVNUDyER67b+r8vJEqlINUZA
8h1rQzcKScbushlLOwM8MudeFDWk29j8AhFBx/EvG4XN2ifSKa25nRaecPWCrSDj
2eR89XaEiOPqRo31p475xn7gxn7nBpWkmBK5SVzzp2b/ceq6/8nEda+2tjA0KAFt
59mwJwtk4UuoOjyRvtXyvSxgtzGKsLYK51NSTB35Vm8AD4cCRELOXRoXPCuyTM7u
CjBpc23hUZb0IYI3OoooJucjkE0cvcBaIOTBC01kcUngRhzRCxRkk6QufMoli4NM
myCRO/Sfrwbfg5rNZ4qDJG58cD2wAmavDw7dCwKirMjpXjictzb+sajI3Bd4PK+F
GgUW0KzVdPcM4GDHck5ChJK9VNIr3yU0H3uXVjdhGrgiuV9xS6r7FhPB0KOHk1fJ
zhGitBlQKavUzPDT0juScBpyYOMDaNtZkb9vyATZPKqnsVxc+jMTkZCRTyGkjOsu
7G2+kbjRVh2CKN85XucS/NSON5n/5g8zirUEQnhnOeJ1HcH/yxiNZIWTkAZyBrSg
rx/Kljq5Wf3luoPDxAsjOgkbiT2TqYeyu3JkUuvSYNKuQwtJc2vXyR4XBiKDpQc3
j87uxomE+9GAtYMcD1Of5PAKa+uVJd/dOMKbaeA6bgRg+v3DOUykUTCNDgyjZYAw
274E8Q3h+AupfGxXW5PRqAi+7dnJdRK59oiajWSFldKYSU2AwYmV6JFM1vCq+QXR
pTmEQ0GDIoerOZMxIXja4A3QaQit7Qy2CvcFP5cECWpsotj4vUTufjnx8MTwgXSb
imsF6c6lGm0uAPW1abxJFB7ozt4nxrkDYcS2GT0kScZBZbeZWUgwDMzYgYajLQh8
1j6lF3Sp70fHIt+r7AWOTfHF/ul6fjLAgutxVM9Gj390t/2UxLEdckyHVL2HFYrx
lhh4Ca2iomEgyZBuN4B423ndImkTfqCLc1Md1/k/IWXYW3iYcIc/zok6EJre5Ivw
qecqSVcMFdvcDeIn0Dhc0ztG0Xo1UMi7y8K7VlXGA0dGgrkh1oUwPbEZQE19Qve+
8RdkiIBbfUwVeqttcEwR86/lDEyXc1yZ6fKOM1s+lmLp7C8SZtYUlmhYUT9Rjwwd
w3eiwPpzHwZrz3klDcu46R7zfUrFe/5f+yzDIBUzVgzVBgwPzwk1xsoQEqlxbDjK
h6Q/OgE4lPk3aVXYf0K8u3wqTmhuMxi9wlDi9wToatdS0PtlDOUoPmDgnzusT3k3
Q+hJO5UcsMFbUDmLLbrKIamizg+3mSoJOcLhFq63liliDBigsgtvcpy/yWiko9Av
fTsyESq3yQKoe6o8hIIGXMWifTe3APmqj5ubPFbAeeb+OfhPid3N3WIDd99EbZ3I
ghO0Rv00f823+fqpGxCcXI0sdCLsr/bMTtH3vCNTyUiomIkLEtOwsETqijPtZSa3
HbPT9CuPstSkVOwfONWx3e0HDQHSdVPajz7jnQYgjCIxivU58MLsrWY0+HfWgX9i
X359TKMxQfSxlJTCfz/tu+Of1p0G4fnGGqCyxeHfAfELtp2nJ9ad2V1o7Y8X9o4C
gXomtyLMJ3s9MV73GTCcSl64KfGfb4baxI43gRXyr/U7aHGeWWr8kFmD4ohnXOoN
7PTPFXaDMfRVp/jS+pYun5ehBE7SAbgVxybVvLFNv1ZORn8E9MWhFT8xDGUeq9Qu
KBjKgLrRvk31dYNSuIQMksZ9lceGQasnIRxCIOW2ZbcJkFR/J04No8t9WHN0zWRv
WghQ8gd+M08Epr1jZ38fT06GTI5URiw1Smhqs7jXTE5xhhP/r1sk3N//olQBHPjX
0OlneFZCxMMC4oXzsSWiS2dr0Cn9pHcGU8ty1r2DWbo0+wKBa+HLl6DNO6ivdKJC
81AVizaSnjVIlaNWcJcnGbcAqvAD0JdQURPBTwL3eO0pZoN0sDA9dY/ysAkI4A21
4BkkTdHm5dgAABZ36Qsk89oTlgqBn7/0TjLQiBTS40Xl+YuxQ9rO4qVy+iWAKbsb
vilbYHFr+daqJ81Rv+3JXIEByB3th96fRTGqM4Q6Onv2tZqk3vnuZsoezdqnTnvr
DqAyYlQBymxQWCacZ44idZaXRPcA0D67lCElpIeV6WD9dCzon7KvxTChSKZaEOIK
66G8pLqnO5soY2KzdHSCZEr7xvidaetWnAd+zGmqj5qcwQSV8L2QSBEZfhYo79WC
St7pttGTsg0TZE8i5volr1fEJzHv0isvjeNtd+Ca0dYUJBzMffmXKbwxlEwimGCf
KtlOwOHxe1D5nu6VD3Qu/sTIttbNtYNjo8E+r2labxKKqvH8UVpTPJUVSzRyT1lt
lhSecPmwvG6Rv3/1+HcznFTq9iWb/EjveC0Lvf/iWZ2+4NqeLfOGefJTIslzTb2h
rwOoxmZ1pVYMLNjYK8OygSQ9VAXOGvcZ1e464z30t3KQgt6f+/Hx7EIcZndbONf8
li8+i8iokK+imZrKl4tuwWgQ65WmUhWBtjOLSs1DRSaKGeWZgDk+WNkV2+3SJHfW
CCD7peXMDgOSvaISCKkaFW835GMsg3GgmhlkFcMdvQQnDeniSLNeR71slt/NZBU5
Dj9BrsMynavUuxfAbZ6C9nI5JvmtkJ5uug79SBHqEJZ4y7Dmjz9uFVjroig0bEiY
rvLl557SCvcPmi/ulvEFcdsIcGwrxfQFaAon4JHuzsaX5kE7W/T6E2POnr8Ys/fz
PKwd1q+QFKhMA1Pt30yAkOgt6GkAJ8U5Xyk+f3qdGGDf97A6gDEaDfYyMhNr/Z3+
5h60/OnUD57oFcgnkA+dgTitb8Ug61wgyvhVvM0vxgMoz0t16wBhd1cSvbGnDm/a
NYYVg3bBtuhTBv/oUI4KpwQC5k5JURrufPWLym7l+zIr43WOxLuJoE+06oay5RvU
EyXykM3Rakr0+cT0HLEWn6nNxaugfbgGhel5BO+B86q14dX58d4Z4b+HTdwA65lT
dwA0mCL+Q4queTQP0LzL7M8IAj2PgxoNyk/UZ7nkBhYCAzhrKy+bYibDNHlQ5Pk2
FZtB4CpHlNmGCIHMENhi7hkBhCjJGfdX8hmknn1CdplzxD2mbLKuygO1DepExi9O
OyKmEpZ3c3oaTbDREQsKCYmyvYZNFsXv9Wgrxlox3StHmCCyfSA4uIrbpzGtMS6O
O/5gwcnbdy1lPuAXvcAj9kRO01kbO5TnG9SlT1UMP2+DfSPDRPsE/jHrx1VKbXzT
EKoBtet4EeIlYT+Sy2EHtH4Z1c9VxL2U6AMsS86qmDLz3qO1LmaYNZT/obAjeArD
7ItbPTBe3AnpMVDpPB0bmNQ6r+HFZWBG+pjzJk1Qf3iXcl8S5LLXt0lnD9qCHbGi
NyG1yxHUJ7l5SfB8Iu2lHeFGwYbmjBjxPwMfFrXFFmN/tNJMPRCK8kHuWqQcJfYy
LzMtau51CVc3yeyUUAp/zvQH+ix7QpA1mQGp4m0pQSuazZGzbBU03qtDDnsEo8a4
cvHswCWYNCOESA1bRnZ4RudcYh34a9fbFis8hRXFp4GSPXLpv9/o0Vns/KN1tOHh
nAh9kyet578XhfbWkd4hauEW6jsM+5/7KvX65MfSUxHyGSkAljKw7S7BAa1zxq1e
fthQ+HyHvTU4x02bpW7WkT6gdXHRBIIls9acf5yA2id99Ex8FdIn5vhfQ1pE2nba
qdiNUUhYR8tDsZwbwgbDtCeXfjcfGapzs+4FgsmKUYyjPxwLn/m9wivZxBSVkHpn
eWVVeaAA6sL88y+MGPeGwX+Slqnm0Js/vpZtDpjDNtNiMUZTL9pWO+0hoXtjt24K
lcWCqk4bwfh9c/FvvFWNL6ya57t4PXLvxiv/L1NL274CKAEo+loN8Gok25je6OQW
hsT7PDrt3gGEFGT1avDpj6RDAhut3hZozbsAMmxv3CaRqIpnAxjogNuRHSujL0IV
juVXnpHnhaPvNbi+8sZmxUQDbNtEvdV0Dtbd1p6lLBW5LAWgePgEuP2zupYXcOsX
RCuZnZKWEn1VHvWxNvoPI8829W27OoH1uJtqRvzsRrnDZJroK/BYEIzhMmrlYMjU
HBXzc0zRXyvcifNKsBoed4+io/0CUtcsSjx2hyxwxRsnNwBlTceUMP3ypXRQsWqX
V5AdPpgCjQUCAESpx2jIzh9/pQn78VAuu2tBccnshJuviWnmGjI1rNMBYNxHnM4B
DQe28fw4r4E9PEZUp9144DxISzqLIgFkDW6dAO4UPKguyyD4SlDxsafgdXpKdTPX
evxv6WrVODPpF+4i6ACOg3BFhMxWbawE0hDa5tob2pzMyWsvr1NaX5lvb1K0jnMQ
Cyhip4Vhlfy3HJ0aOo2qVUd88os2Lmf5WPTKmOBOmRy6YrT4CmZ8vd8jSUImT1sD
eQBv2VAVmTHMDqhqYqqaGHJsvvWlp3BGr82SljnI23dsDcg8r6sGsyeQTy1V3YGw
/W5JAIUq1+9Sd6xIMDr10XlumW6eWRr5nByQ6vv5TPxw2F84ZkkO7LGMptdwVzdi
bfnG0yasD/1wSp/fKPItuqkIG+twh9AzMPmi8cS1MPzdDevkUKSnZtWXak9eLUSg
jj1VTAE1Irp1GjPitfhOrAWJWv5902XjNv9CejEDIsVwJKEmov1InYQ9PzH+a4FS
3Xkf8hmvOm3IbskPDbgzZtme4+XcjjNgCj6fNrlkBzymgm09hjjmA3eWcqzyloJX
mmnsdCDYCkxr8C4N5jOJ/Du6V+E6dOTTgp5NloGW/yPAHgnHQnlqCY7HQ6OPviF0
WbIOf+v+qM5O2xWWyx+x0vGKyG0kbIcZZs0Yt5OROBJsTThSqZA12s6zlQazSH4x
5u7a5tSVXsraltD3J/DEGLEqSvqfzWVFEERyYSnXl+Fzzo6hxy69FyszbyuIqjhr
ZEhtXELxq/KpxuQ1QtDLjks2CNDIQ9bo9OVJj+lRJ+/CjlYQcxdcgGP3LQ3jyOZ4
vKN/OQiU0+2WHPYN3IVyKEAXq32rfcAF1spvVa2Awj7SlTyqZcSX1xvWXQ9XYcXD
cuNt7n1Ey5dArsW0CSvnL0iREcYQxva7DSev0XJc+SpAPNrNUcaLapTyxABQMj3r
MmZSRG+ulUerHm+0T9Ah4N4Y+hBg8k7SO/K/YD1ysNGWU3w629FhlI7u0DcJ7+fK
ZzAfJQ9k2kISPkIo7NkfYz0rlaZ9ZAeDQRCM7jugMxJclN9G99c6spizAQZe7KR4
cAecIbSwI/wI0pA0bgMOsfuopJoafI2Ziutaf83Lu7S8lAfCI3EkoA3xCU8kPxBy
3i/z7a0licsAg8FeXjtJ0qlt/ffc6LZD55w5Ys+nEx53OIp2HQGOa9BW2uy+41r4
MKlx57yWRB3cXOjO7apd6TvEwJeuTBvwguG5mEvXOJmvMfUKWjrlRQHPUhe07XHu
nTKcpWdx7gr/vBo4NgrbPXmrF4A6ss+3FD6kUFIHrzqsJAVLDiJhwdR7KPhyVlSh
DmcSRBhgG+6DU5roM1bZspd6BOjdARXZIMwf1rv6nM+KHvt0rQ2KtvV7b3YwWjZy
s8FdUDTJF9B+RluYalrtn7AAqyogSKT89ZHgZ5ERtrcsRS4lCqvesg6UkB+jZNHJ
QoOvxwOJSTfi/dZ+8rpIShdnPGbcVwzztTLmZArc4jdSuRasiV3x0/AqysgnQhVt
TgAGr/W6R87MzNE9V4UlGHL1J+7N19ifZl0UuIoRsCuN+smgfsauJsynhHLs0XvG
kIedPAOBjkSqHRiZyLruINuRnyRQAfy9aeOA9ptS9DTxD1AI+quFd0Z3LhHiFBdX
Ptuml+/QSFVQ8jxrPV8rUKer+xWOj+fLrmTx5bNc3r60hv9QZOSx7ZDa19YJ/hsA
WY+W+lHirKqxCs90jhibWr64PYWeR9qEQBvmk5IoqBNluc3m0VoAWIqgy259QdWj
g3e1+T624pQuCs/I9aSiCSHgeq3mmMw/3OHL51PRH29Ia3BqKHIWrs2svwVrDiJl
B8TRkGKVsUK3Od+5wgyxctrvfF6+Ba72OnnLcupMKUETq5rYzx+IG3zEwfa0Xcoc
/xwbJjtbBh4DGLYXRJ2fLVNyKar377OWQ/MRum2AJm82yrPzr1tVkzzL3R4g5skQ
8LOv3z1upvdWy8yLhjiA5cPOr9oL2Goof6ZunBH8mpF3FRZUIqsMt9y+gJJ6hK2M
mKY0z8xTSst2ZLQGVQre9UdF0yeBRnRbmrrzt9dgtSozM5XEn/tsKU2V8JyZxeYj
i7Ebiwj/kMoM9nz1bz3OUuJ/Ddj0L1jXRz0Az7d1hCg5M8x9PxLPk75axORtnlhY
L7c+emmuZsL2gSoif4PQIoiyRvlsUuuxJ86nGb5c0rwHN3XhodI7H9QZkHX9CrlA
p7+CiDDjFUEgVz1kCZqdYCS2F16jJi+7/Ox+SpRRCtU4RL0g7O8JuH80ni3NhzKA
0ogp0i4ZPz9QmEphZBgqcnfbCptFZM+s9tDKnCJuOj2lZ2lt5i7qa5riQY/Z2Jwr
2R8KtLIWldI+ntKqWRN21Q3QdcGFhDvmFYXEvmbM6R/lphrULl1Xee7EiOajcbGM
ERurAE+Ez/22olNy65lVs5oI0499Cc7uXi+rN2SQwcb2xnTy7vOamTQIVL78ptTI
4ExzaW7y8Y+WjQ7+vdICcSv2ytzjCFCxgxotx8EssWD41b4+QV/E14Fw6TD7Ds4W
n5D/DIg8M5lPZjl60xFSQS4Rkf0GNcH7JvGV5BH0iNe2N0FjzdItjz6LUMyCisdH
G6UJ8QsPg5AqTkZMEy4R54WURUhn/BXb/sq2javYxVlFzK2063n741+OElc+YTiH
lNUx3VLDWVjhnahiILeiZgJfk3kOtfQ/crfmN5R0yEOkxasv5eXll6d2SiyNxxdI
Q1FTuSyGPQjT2hVlQotdSGQzv1/535+kCsC5z9yEFPubZVFeCPh1I8HkvrW52kOw
a0GXkvQBxAkje8EEf4JKPhA1Msmyn6i0UX8ru7/2qTBbA5mUcL2/9URp+DH4bt/Y
th0cY3+PD5riSl62A60DhL2QUyO/No7bJIDwgBcPfjkD5IaLaTcSsW2IoGQXyZ5j
RRfSBkirCMzGXobRMPoYCdXNeIn7o3a2c2aDuIWzx/q/3hPxv63z66YRFtqE7FKM
yOcoN//Fn2duR0LgXKcz/YplpHqIm1FWFB12TxMWTr18mNwqilbJbSCyiiyLJJ9I
YynPTVi1i9ERhnhGDDjbnA21iDZ5xTQnsFOyXzX7KX6QYlpDrcG+nPH6gm+SCwej
8+LIilNgRgm/uHiRyQxldaquK9mClp55eN62q1DKNbrNP19f9zYcMqIJYdibSG7N
U3ptylxmNsqnBUk8eTFOTJUxaL1sHobRK5Hqrk5t/0MSbvEMMaBRt45MHTGa/DaK
636HlvHv4glHhN1VDl1Cbm9U0aWEP3cvFQ8rniA4F7pVVHrxdyvLyCFClNScVYRC
zQbADS5G4m6yxyaDX0pr2DqcbGTbfVby0dJw475PGxJc4npqJMusOxpw4L1VxSSq
vpEAzi9Ll16LdkktoJZHL3seRtXt+5c7QfIBCkrJQpYTlJJgVtOMifUSdHfa3MQ5
ukwhjGDELz6pJi58KDlFTK/MPhb6p2xGNvSRSO6e/VgpTVnHsnIpcxrbfZamjYsV
uH/EZ2nuxkxz7EWcbXMzpp7IwrkVoZA/LpT0KiqnMa7jsIxqhfUB4dmZZ8hYn/d+
znaosfdFr4+FbAAmHgfSw1QPUz8rY4se5ki2YkkRWqiCYgnVE9JRZovdh+dWQfQ2
ZfPkTGqxowdCu+wa9bS0ad2Jeu20C6Oy+Dm8fnMeE9vMFZeqtqs9xQYLAvTIWKr8
tsqDksYBrAck9ff21V5wUHtqQQDntiHPfkmFJOc2DzHmmpti87U4+I8stNG/V8NJ
IpQXbkGYxRnDDOPFW2JX/r6a9JJyBOUUZmvYI3jaEw0mrerWETcxn8X79hdX404m
qxyN0qbmeLx41k6/ttffhl7Xq6v0d8eCQGd+bETqBOW2YbmvHus5R9fxQsdvizb/
18XeV3+6mhXlUNLEhqysrZAWDGTVJnXVIg741EsIoS5iErCDtL127t9nPE/YBqSS
gBrCkSTJriCUuLih68zS5Ie4LgcVS8wrQuUQGOXwpdJcBIUY8tcReMx5SxFnp2WX
JNfnyp/ntta6iuYNIRKEWJYvnIyoclDR2HTEZSl8/yAs6rjr5pR8sKEvhRpwabXV
txKB1f6E3x+17MbCED+o8Enr1WPXEtP3tM6kA4LLiJVVWJUhFXeiYidplV6p2Y+y
bRkAt7Vgcs2EXA6YUT+JK/TkGRh5lQX7elLEi2iza+CBafyxeBGJ30G3pYNf0Pu4
Mlp8guk86TAkQjlRCeUd0k4incc5MsX/DzqCM0wUftmz1VtAxMCqLEtegmG/q8Yl
Ar6egreWhaeTXNy+8ZXPpAm8HunQkqVS8TifP7RJk0qkSs53xL4eo5ggICcFdW1x
2QnUORhxfnUu+Ax33E80ibM6GQS1aopsf0OAO+ucx18mBNTI8x+DWIvE9I1g3IJ/
UzoDC2EFHIpqA5Ncl1xEvJwxs910+k/bAJDuYQfHwSoPCTuhmBX92saOZymgheUn
4QenZmZLtHecczoL3PUlpKDPLdLHW6kZJZwy7XZVSbGrAB2u8YlFqlNFtDn1Z2cR
TC2KdO0SFXkCY2RFLh+6kVJr//62v8l6+jF88wOoWTK+455I+t/5z0A05OOI0qOi
dBjLpHEBOxRn55GRAanTLd2q0WNlokEMQ9327bdNfWtX57j+UxavwFmn0Lfj8TLX
XJ9+zRJp2q9KTav9pF/PE68uGwCckrByHGMATo6hLlOxcxqy5UAOijfw4eihq0r8
iBUC1z2W2DaGMCup4g45zE6uIj9e5L1XPYD+kP37lORxiNeogdfZeaCYl6LHOtBH
uusjoRZfzw1iXM3MgOZvxDeUp8srIsQ+H/7iDlQ9irdyIeO6IEXNet2ZmJimpF7O
C0OG9dVCd0ScO4Cn9B0MiWpVBSPHrHxIwGomE7K2L9SuQ5R+g61mMomqcfww6Dd8
kaJxJFXcNg8RB6X8omdcWXuwFk+ruqKEskcLhvk7AXozUrD7bd7Y907o4sF2IK4l
LfKvVUuYkh2wEyEw41O6loG+aXUqkwkitnu+BZxQnDpvvOcWAkzy2SccCEtG9KIo
AwRLLMmdL4R97TiVI+0+IA6//dU7zJfk7u0ErgFX4kAB3L9ZnQUkDZoTmiRDm8uu
o0rS3dgoXKnNutUB2xNOjWXlWNQ/LDcgEjsSz6+hB6bTZKnxJbWzddj4qvHYzoS6
Gpix+me7b81nXJKIuA5JPJWxQF1OWrc5kfTfrkwDuhLhBHsSv9aIDCWYr8xFBb/0
Qce9qKPwpIeTHSyz/OzfvjfTA575XKS5gKVA+YBW/ebF/6hbtIq90QbFz8zlT83H
x4HM0hZoip/1FiGUe0wGNRmhkwdTxlOKvH+pFPEY+Wy91UZVOiQ1ieEvXQ/MLRMu
B5V+le9HOj5OKyybrN/mF0ao0yXsMbcZnblArKOinSHrIFq8BL7sW1LJhAdTiSpo
O7sddPmMjnTiO425JVjc0M5qCWiPKCl247T8NQSdy6TY3t8l7yAshnBOlu/xcu+r
F7dQ1nLxnxUBXcwzXz2LmtoZmpLFD8wC3h6ToOgCPFhWOAnm16Y23AD//x88XRgH
sFEbwZMgsjPPt3eDaXk2afNbk8XkfRRZ30CGEhVuk4mnJn65nzsMSBpTASI1wvrk
FV4whTsJXZiVqMII7Gh4dNgLkheEH5jPh9aRGfKqbT1Euvr5TajnJpkZ1lEkvk1K
O5AdFtUYRIoKlHi9DPNPzYfoW+C8mMFEe53JLmHxtQAi9Ei6yYOgJngbvYpjU/6S
Mung00Na1U8w8+u9rhepBEgt8g3w7ru/YULcMmhzaU+488vDY1F6XU0Y093+OtEx
FXiKejQ3Br4Ld+M/he8xry92Kjnx7KZ0IhBNbJygAEHJsST99ZuBxA9o0BNLv3sB
NP4HeCUdLcaFYZTFg3zfNgezmEGaTBT7jH6zlminXCOE76ZxkXfuJFTQVf9QOyit
Wg3bleo6+3boAJebe9Y8dOWyKgK1rO3HHxhf+e5qeG8Auhwy4xChMcrQbgac6LLx
v/f8Dy8ORgkR5YNkLQL4THM+6oerh4/7aVV70QBz4oN3ZZSGsnejIhysWdiyLR52
4k662IvE02y6eQ4USf5FPvWJoChXoGuur/A3u6K8gQX3Jvo65zAKT2NkNMSJaKil
ixt9P6gA1jWYG+A04SGbMxrtE3vvSPU39kI1rfSgL3L2DUyRmEaMKsw1cmOHbkd0
wIjJoXEVycJpl/Mlyr1gpF2pi+wS/X1yFbpk2pTUl/IRU6pNVDV5EIF6pvfWipj1
LwOJBzSlY7D9e55UmZZ3P2WyFneUDcXGWWJulzl28A06fTMTuz7EqtSXSccghpGI
EUHqhYqnxLQ9/r0TS/ZFq5wfmWkBiu8ygJwPg6Y3xtWxgkBYhdeU4OPaxGdKKNdg
qO3ppjeeb5AqZKpmNtPyJp/idblTnYcU0XAy7A34ARK2OxbK1nHFvnesWoOMhNqG
dVl/6IgsLtWKx7nqDSSwwKm6huG+1s92nhtkMpH9ZrnkDZdqkO4Ok7MU0/Lvnukt
ZsFUc6BJkK8oE/fvtd8wQwb12DQWBZO+PV+pH0NGmQq/yZkAXIukYZNDwy38xKiO
27PBrQFrFMDpfddVx5hVHgrCav5n0n3CtOQf7RLOdWj1maxsHj6of8CFUTGd3Bzp
O4MtWUYYcSYXOrrunlCEEhoAjkMRTd2sOPltzOoN/D+ijIVbDfbHtCN3hyAqVBQI
z//YpGMJc9swWFV4OHiYIbzONwHxvJvrmgPlfX3dGDxyWeEfqJ6h92GA6CkyejUt
3co6LOrrVbMXyJQx9FqfgaeG4ILVXTq3xabVI0J8YIkjlhkupp+Ku6DyKbRkFZk3
bXDL6Lp9jl/HB/fPG79DMGwaZr8LLWRXq7U9f4UuSdwHCKmAbqgHiiDxOgZVfHdE
HLXcjZ8u9Uhroq6QLqwqlKsMUGjQlrk8Ohw/sg0jv+cR3Oymngt6J+xIM+fbS6Pa
66DXhZWHxHx/qUIlW5Qcdyrbr4rxDLLb5arH/g5X67DCBYeW8MHQzMSNmR/se2mh
zhD0G413QQNOPWHjS3Yf2myAIjDMQFEbUeFg08DGGYTeDSgep9yWg+MiCjYVdC5l
9M7JdvF8jE0sNt7/pGXxdSyQNLbwLgsj2G0Kp5eTtBA9INiMye5VzreeShLBIwq7
LgI3zg1Vc1yw60IGjZZ3/6olograxHoymdTXBDY+MuaNnBlwVu4WmoLCA7VkQnn9
J4OGHdaZN09izLrpF0vFjaDNVBpgbxQwbOYelCK9XizcFuqAQUbm/JQlbudscgNG
nulV4WLqSsgcKhEBIZUbppPFc/xrxfT3WUqjpNsJSphZgEPzZpJwKZy9Cj5BeNM6
ZsrlA8bhRfPoR763s3F6u/W6I/KvSdZF7GjWRVPjVx8odPKmUrGxGI48mfmQBeb9
CJOCDNLDxKqqm+fi+DHtfjFwCxGKVthkAItRZENu44Mo2mUOI1Zljrsn9ZZtouKr
SS4udiEl2qJ27SCCNUe/C0xu1b22aecugYPUfxKiT+4Z5sl7rtRHpAWDNOSNhdx1
30/NBxjQLg4iMH3ORBhxKcFQbAVEGqqI5/liIeJV/jLNw2QcA2bMqFjpzTRKHbTf
nPx9DDHD2Zf9uM3UovW/IRc4jydcS72Y0NE485KeACnCsTch86qHHz6STkNU7KJN
V9i3QSHPbnbJ/fFVrAWprdAbq7YPtW6Jui7fCHdsxNWK6V+W5XvknKKl1LRlwclw
DBQolOcWp6Wu11Yg8rb95mKl3mGAOEE+4St0fJETKNeYDh6wzVFHtGj3Zi138VJu
YHK6+gsteNGGxJi9yi0EPMPBwK2MD+b1xRe4UAeX3AQrQhKg2edTh+tq0RTiLOSw
AOr1Xn+poxNZiV5o8jEC84p6OcmrXohOpf5vaXOfMjDMcaqz5a0p8tBq7tTPBtpk
pHaK7mSTnKHZt+hZ4pqiec0D8cYIF4U5fyxzLhmofV7LXwr2RNbRA8a1DWP6Nel9
yarIbUvxuz7+30hNOvsGuUbdnPj2bL1QIq/brtM7kNEAft2SJnu94hg/cF7FH2nv
TmQZJil+1uXembrPWmoGRfmXHGXGF4FPgQFzaDtWg5VBaPzlGHbCbWDjX1K50x35
dEbMatl9P9u6m2lc9YdZsJxRDKYoIAYrZACdtruuitRWk7pj1CMONfF2rFo3yBmc
vTJ2ng3c8kPSpgMmC3wm3ctY1X7WMTrbY2Ps9KjtCKARtONGRghMsOeTCcnx8Gi1
otSkfoDV/lSjenCx0QlfFg7y/evn4O7Xc4cZ1f54IMoMdKOazOVxGXdHOn4zFrZv
P+zU/P79h3GKLJDWZhU84w/teOfRfkGDOsXk3B/LJzj+BbjSt/fUaT1TE0GhUs9r
o0nEdc0bwtIp72u0v1Z5UYK8+Us+c/mQsy0yoGAOsQK06xi7iZNf2EtezpPc9+Wb
bDXwWCND246LgqzOV8G/0OyAhPvf4slra192C1UwAkiztgXWgQQYgl67GsjRd0SL
fOUt4xDPfrXgrVUCl7IgKH1cY3Mt3hHabDkZwvSojqMKCLdYZTbkMJRKZqAtRIt2
mUucIyFW2sOjerCuHCoMdAnpj1B8YowwnAUGc2xl3Qy+HgTG57G/Q5TV4rVk9QHi
kcuvV9JW5EKc9ZkhpKi+WNBxfaChazv/ydUJI1YHAWsJXqsgx7P8tYADuohJLgJn
K+LcGH5RONG0VxvxNUMTTFI8oOVyUHWxAGje/TBSJLboCO0WwewI7k0RDloT/0wE
Qsj47uGz5Qwp/WAM1VewBKf3AkeY3HJvB7HfrL/F37giFigmUMHsFDrDD1tgCrIB
2Jk9ESYJ8544XTDAMXzMNAoZ+IvRZB2/8+C/4/ATlXjxstv60N2cGSZSXfNAqDfO
g4EVSNxVa5RXhuyvJY+b9ZUjvntfatdzCmQhkQoGAtZPiB4ZH39csvfNdrLSA511
c/de4I4K7JS6EcGh3Trq7IJFE57HmFuXt9VmhMSryxtB4UstZ+u3zZThQj8endxc
9iX5PFmumkXkfoouA/nB9Zgqd6CIC5yjU3cQvFPFJRqJGS9hkcbHKTVK6ggqnABu
JWlYRJCnBrR3pmAOD2B6W2nCq6s4RIspPx2L/iBPcRAl4MPkhL9zbxC+78I5iH5e
XJNjz3EGGE9srnt6j8XX70YAtOEvv/3gGvvKnt65lBKCd+4LI3AjdTqz8AHtX0wz
MYcV7wcPKeMZ9lcDSiGa67dF7cxZW4JrkHi2gP4M2Tsnvq6PjP9xZi4484TyM7EN
12tx4V6mrDlOCFHnp51ONW+kijEt2v2QR3UDf0ta3M5ZniOUZGHx9IzXyWpWbA7k
LaFPKcmvV/RcK/5nAYRJXOPVPfvhWxiMprSlj/AXCHF2ZBjj3qGfCWx4WDZURl7s
lruygo8fsGOV4PG0Z6MMYOXNTzRhmUr/40Loh5VTMC9nrhc/I8JLZNpgX2DgJA/1
S8855Toasovj4SuOsMjvOUg4jNaITudhf8lEv4QkolyduRQtdg5PJyzPjd4zNIP9
t8jX7cVRdJ6g5wPyg1Ia8p0nEgSfME/FsIPXD2UXEpSQhI45LGhPf4SwFYSg0h1z
S2S9dA7xb/kOYtUMdmfoSWHw3ldXRQ84vvL7wHYGmMMHUjuhgTaM2xgl6d/eZMUJ
lM7PI9lPsDxIQ8JoTA4dporSgcanMIMxyfIXt9xqXpGU4RwmxT8GgEaAQ6CDDeKu
AtyvviVDpdJ36BFlnokFI2o5DBzRpo9qA/IS5ucUHdA6mR84CQMUxMJ0k4m7fCR5
kPotyjvwjWJDV6LAC5gMUkttBx8P34SMgAP/SpPoBo7jVv2RvdHnlCH4A9wwdvzQ
AvEAuTXl/lKt4eAUpzmfHxR4jZirFwuvOkS74oOXugHKcBWXjUl++rjU4gT8Onh2
YYSlXSO8pITl7sAlD/4+xJYAVSGkLU3vuKvV17iP81vagHI/7MVmTICn/qPW4Len
MDxfygTx/JkOC/Fxoky5eoLEODF+8f7KsYizvuXmmm9pW9tD8padtkY/DvRMAR1x
TyyFUMym3zAcXfzjlge30v9tybHJCkAIuVFQp7POx+XVK1i6wTlynoJoeZsuDKLu
OTWMIGA4C+7Jdu36+suMMo8rXXjg3/2xGCSBFPK2F9+ernXI5GbRngLzUsQGLwq9
pQD7NXc8sIdaCBHzMGMqKev0gIeT5yEjkJ7uP9Dw5BXYNI84h0RpUqYVs4KRhzYO
vozQ+GTlBvGx1kuhX0g7T+xZCuNI6eTvHjiDFvKxb7a/gLH2o2fP2RHxUXJD9Z1O
+NLe+S8XkZpjmFYQQ8DDWQHGKCaap1wDg+kqOfUEaf9SO/wUBTUZi+peccU7NcVs
7MkhCWKZwerFu0pPgaTy1rbyw7h8R6Ls9RvtWRbw3GeX0bJX4Z8oFAmERQPipBbb
LI/FLGK9/AUvKze3JcpTHMULBxqRiTxxLnstn9I41t36Uo+dlhXGZu810SnHgU4F
fh2ENGX7lpBNstsaE/UOIP9pZC3TvM2OI1OqcrPiNhjIvvmucp+WGApn+spdQva7
n8Ilj2VZdVAyJiLEbPXuiJ/PGre8yTPymBxsyI50m70n3ie1XS+mRD50klh0mu0F
/IE+42/zuxdCsD9MPwHpP22Ni8KsH8ZZhDt7HSRIMGqLgqLxrbGTfD+Wjyne+aiD
NIniMWIEJBxo8tPLb83ly8BLqu3zYKDmct0SUAGcvGDPH7IS2sWbKgjWQmj+bgHY
I52R1tXmIhW+KsJ+X4Xnh1kyuVhEqtZ92SUA1dwD+cHrR56twCwB0PMnbgntmBL0
rn5rVJrNh1KVeE7sDh5RanjqV1xAC+gS5+PZTfxdeglf/A9NvUplgiZeuWMRFJBr
gbnw1aRRsa2OWTWG3ZaPm+bgMs9QWArwEU48TLTiBH5yYzHJrs5WzxTwR6EQnlQI
lYdFwdS5M0nqbIn8TIVkY5/GxM7lPriu8vxgmeJ3CS7RBCXtBFOkBpLx6h0Lb7lh
5XwGR6sR84mgUvsph05xS6/vdbJFSupGwvmlNiIVBjCltmJUNKbFXYRlwTckxe34
jUH0ThhgZc2LrRKzvtAYcswY5bgnmwjwM6IF4FRwbITqLSIpvb0lOhkDWhsOhti+
qcj18hq9kfzDxnLINtA6BbI15h61YPR7hMx97TNwr1ljF30VLHrEswkMKt6YqX9v
43jJ+R8cRPmucz7Afhn054jn2JtiJ3oSh472EVpa8ML11mg1AKUTfEfWQPy1x2Ba
R3t1MNckI5KgjsEOa12uLl0YRR/cqzScj4LWyB5unr02mnU8SzjAe2etwXbCmzxW
L0Y/ioeh7I+0YAA1pdlapHIa+VQsSg3yhp5OtumefHT6wy0PuE9cQlIqvxtollUG
wmRpv2zDKXnsdUfG53NgBab0IRUv6kdgjesUmAaxKW6gIElB3MfKa7bCD+MsL593
mzL2DSE7/UH/egFD0cx13SiUJjgtGkgUWf+snLNt8nRsHvPKoh6M5I4IxCz6B2wJ
/i56tgUD9BNf0SQ2WWL8L0vE2H62MjCt3KvhYeQz7xIoQpze1YNFOA5egSHsxqgL
J4C8znN2IQnk8c5GmtUy8i2+4IvRTvxVPAPKl7w5Q8svxJ7ZXIUYM/67/KJmctJH
PF9o1pX9PzJXAtQb1a26NPpnjjkVwvc/jrz/6PRmiyU/jwCYVMKAqDpvGhtFE30q
/waYYXk9zwrGrCGwXQEdZTrBPL5Ibtkbbflz6iZ+hA/w34bmzENI8sTHmhj/QjfA
7n4fcOJqXKnG5WJPGvQW7dGcLIgyiy6w4W5jAZrTD6sMvZxhSN26MeabPh9Wwo6u
cltmMRZ/Uvp46yYjwV3pBWAS6zGCKqZiGCIaN5LLIczffJSZe7WRkmIL6fOlxUNk
8iLkEO5tobafNHn1v5nexOR+RCq62eBo4y31d0FHT8KCBedoWC+lTZew4C5+LCEE
MThIJCmozRKQj4ylIFwJht9kbOlPkQZrFCpU1MpTHFbqxdg8zueig+P6FyF2Liyr
EeH5Sdf+ceuw420BA3RGU2Yns2srYKZ3fXL2MB1bMYlyEcJBgi4M3ewUZX++kqLa
f2Mh5U+RsKjLiteIWu7LrHGGWDY0KDd7HytxRV2vDGZQhVrfjjkNSE9kTOnidker
lJUMBs6bcA7Jika7AMbGtaJD8tHOpTqe1Du0yLBp8/qpxu6POdUayYl3HVUd6/Jq
3ClFBEKJzKk2NeKecdu7T9eK8VuXZRkBilLGTTgcyUez0qE7IVWNanv0fEan1wiL
oXvP6+QsNyUswnrXGoSTSBQ+Pp3DfTZBBReIhYW7urj+fr4cyz+pSHiQsERVj2pO
S2gb27Z5hyR4yNC2uQhV98rI80ql+trkwQrK6Ew25IUJYWB59JgL/xaqR4VA/elr
tdZVS/GN8pgbTARjvoeCACJLUgm07jDjLhT/6i4JRlcazjE+fFXgCpJz7GBLALpC
jZ7JYUMxkO3SOGoRDLCnSf2IqsC/DVKAUZhlNIAl+E+lcrxSwsNAJ1ghCE52cTap
TcsRfBxdeMBFQndRd0Mgz6VKkCNzJvnytg6hB74UYd4v6mMDpQMJ7+PYz6FkHW5F
m0T1ILnyGz2E2rvHrnPEVV8PMrq9tej1eKV8VFMoO8DVbLwZPd2jGo5kt2oDztTo
zrbbDzeM9KOy/kfR2Nba94yGOwS+nVzgKLkb7EQchvvyso2xDpXA22/XSy77YpKL
DHpLUVYJ8zgiskhby4A1AlUbN2M439FRuvRuflNBQ+14V53pvDeAPuTNzAshxWjT
AOSxquFTPyjOrXzd8b13TcD4dA1czRkrqmBEt/cQAgZKlmuZnJkSuCV/amI7cqAt
MkCAh+nxZ7gHLNvFFvtRi7rxMyExXVGFH/tvDf6oRJch6rk2LRW24zFo2+3Mec2d
7OuLxtW+KdqsQ2WnU1wSF3OcwOfiKTUn31I3tsKQG4bdekaesXyOW80r6IYiKj1Q
eI/16UEsolCnDlFmQDl5mbgE9ZLYgzRcNTJw7jCJvJdTEArislk1sOna7GtnjaK/
kx75uNegPznygIfjstVBNy20JM+NMqY84f0arma5fZdpdxAfnh9xjb0Z8uUDawhH
10fic70shdet/FmkNiKmpJT0vu+gXEYkrC0Jtg5E3we81N19TWvwTgaqXa+nuTQc
czJpyUkndOlnphkTtQNk1RlS4YJb+6wxnTTTb9F0443jewz924pfFlQokUvHKghV
7CMxElCYf0zrOkvWLx8smT1jzUDzaRb3pPFcDkOcGF7Uvky14hnh7kJ3xKe02F0p
KHjmR9/JMS8fSi9PkCxEIydfMSqKgdSjnZZ/hplYwt6aRgKnRhm9zRC4HKEnaq+4
maAzLcaK91CjQF+NIkjEb70W9vdLzRgVn0jstkO5I31n7TmWc8xw4TvRaG6cX3Ll
gwvO+fDAH6Ti1aBy1Lc7fvg4Rp4s/W2aTHtuLdv3zA4b1R4+MKuE2YkdwQgTotcx
dBnbXECHYde2g8AnPrZ7PjW+q7JmCi5eWgMw/pXBdkRVw5y1KX/M7obc50ln6IyC
2gI150//YSlkHbZb3izy2YjZWAxEQe+SUDug278xcJdrGi+4sM6fUnU2xN/k+Kll
03Gs88aMgA4xvXI2ODhCR8+jZD5xckfGnqByAFMGdpXTk/b87GkDYOyDG+UQqYH4
yn/kuHIgj9HNS2doX22ff5iEykdmE57JVq/ZaGrX7rjcPEqZPHiriao4kgkw+Hkx
x1dF59yA7+4TseQr9Ja67yyNCTST+1Ak6lWv2icEM92tX9TXJ8EqODJYEUtiBwQB
Rv33iRXW6rV6qakeY7ChIoJfUixiotnGUOI2AjOBP226PFDQQfW7AuONoXAervIe
hHFIeIhVxtyYfK+YUrwdi0B0ycJZEzaSluSjeaCadydGHF58Awr79VWlI8T+63VU
egC2tNFZTHyBG2zSZCCkAnP/fXTCxhVbwqJvh/VFpbSAxqzu+pxUtHdoW9vSOmjC
C+c4YB9Qf1L2dz9Ab3Zil/1fvmLlpkTTyITL5F6DGrZyKP6/NuCaTsHqtzo6bvIN
DUiDDVQPP/EORtHRnvCBWhYhzSnKAhzzetEYC80rqu0e1hhVQcGgTCjkKNoYJ7h+
lZO8NRoTX42Txl7QK+/GWgqiUkywYU/wuF4/4ywOKe/WwZ/2FznoPZv6pJzISUWs
yLdMknfhewNRvPrC9jD362oTB2cHM9oBrQvjvsgeqE3kqTTs4UG3vOmKYxmyDdFX
Jhduv4dN77xCerEhEV56x8TfVNe0Jf6nc44ekadQgv/Kl8/rvmxfQLN7S54i40xJ
NlQcV+vRszAPXlKeMd9vOjsaWwjMhtVhh2TI1Frdz4hOCdMWCSvtdzTYA/U1iWUP
JFu7HcGyxHL1GrLLxBuHR4IUaDNw0qLnUmnmutOqy/UTv0GKDdDqtlhBmnjOfb+D
A1L5NWeysm0tsOjbAompr4yCYcxFnv8ym2aRCwt9ocCA9U9xQB6Lv2SCW2LOMZhM
dSQcoNgeOixfjfnWfZpXuIHLHhhcTvxCVImiTWsGpPhh6rJcdQX2+pg2KTtzDW0C
Dyn/+D9p57ZxwG5kpaumzIf9Efi34FfZnVBYwSqzwXBfO+9POXWyF8ER6LhlrQJQ
ZrMwEzoN2e8G4iKzCgRjBpda+o+Ke3EY54P/VaJezhYWsNERsTYzFw03ZYPs2O/4
nKxVdvxKH9BwALoPWHCYY627wLeCifaDD2yOmoDlANhDEMtp3AJ4r81mkyLeezyt
xjWEtuqeyAnCp0zCti7EkZr7t6a8oxd06Vj736bp00i9OqGN+gNnYSBZoJmkeFmz
IMvV40F8h6ssctJp2VQwvd/Gv06pdYflBAGBKR0QCthdmrS/WMXWStSQ3lILb0/m
cQU+sAtZd2+7ZTprFl/nNEriH3NTjBTa2a4nF1jEQQKdHV2GCaDsv0EtICGSf05F
e3/946gm0u0nFfli2wPWMnPQyVPe3W3TVYNqa/TBQCvy1W/n8j4LVX9/HRSOey0J
G/WvmCVPtz/tOsa//P9P6O66aQfdVQrgRA0vDuIbW04cn30Pn8ry0xci9fa7LuWe
2R7yglUbdN+C+J2/0pTfubjfXA0HyVD0f7G03EzRyYZhN1+K9CLBcdQmOXnOXMbY
jOBdh8efTMOytBeBkDPhxvzkbbVxrzr9G4vdkXuxsApCUQlzhgnkzEyosUuZ7RwD
XqV5pr0aOwzsH3YWg5LzoVnZVCnxKlKPuY0eB/eE34G/pXOtoZYBK8l/UchOEgae
uUsg122xMoc+xuqQRiMpIImN96rbZZttPn1hxTVepnJH/xJTOA4uvth5e/eaUZs3
O/lIogeLF7fXqRT9TtTEGTuZTz5Efuie+Ip9TyN9bBtqopUif13WAd9CTOeqtty7
Z2Ywy0AiqhYiyGMn0XVE16hQX9jY+XAvgYIR59qkZy4/w+x/TqPr2cm/uDs0pxZ7
cIWEjdeQH8BvNTdClfH7JsAHeDWY+BnQwLfufUmMfbKfu1RLFhDpYbbhzYnOkIyZ
99+AAAoYpuNyuD+YxhGr/18fykVkIRBvrMrn4jvYzQNaVIYmqWaaKTU0w6ALuMer
HSRAOXsHicbMa/biVhQCcWOiTdRXRRyvOqJR2e79sA0h3o+f1NPLMmV90IDI8f4O
Qo3RwOdfZdudrjhX6XZ9WKMqPCQUdailZuJrHTUJo0N7diyZDlR3QJXXT55zohL7
qqOgDAQdLaaomMw6w8ss48z7K3r0waREu0C3sLhm3G93l+260AaLubs+shr4YdQt
bQbWr9ltl322bjL2JTyw5TXi/0XsidKyrVhx1/y/Uey7V308TT5GrGNvMZKLQe1b
4pscpYV9LJVNIHfayIkR07A4o6P17DQmkW24GRcRZImxWhfTyFDFa8xlCUxevqqy
IeXUH0VpUeKN5MTuZFztp0jm8x9HZo//OCd0LH//monNlK58aU4N/b2f58b6Zjmi
Si2BG3WaB32VErLIEwwKIH8Gi390JKzpjnghdjunM6C6Tto6g/iBLAZjece21fiv
y9sbBLRSeUDYN61ICPb4QmfF/gP3pDUHp+B7GMYodTZP6nDfRVpO20kpfo/1Ftko
33hPTvamaYbaYVBz8dVq2OtVmsa4rnYvM4SHk4TX64an6qafhIJw8TIrf4mrQwnd
HO9RYGh/95ysUaCkyuHJxiYcWMVXn19vxcCWzKlGYeS+bGXvF8NZymcl7PAB+E7H
nYf8yXW4H/D9MpCgIqvLbD+67oHx7O4ZQastiHiXt7CJXn8yiN8J9xayp7NK22Bt
bsVaM3ROpR1gvzvAzi31H4kEb5k3+vhK3YCnJFrh7Ci7XThCPQdQMYw1hG3RrG4t
uf+1qVnFyJuE3Qeh0wDmxQp1hMwFmLqCmL8MLSAdjRofc9jIPtiaDkvL44+3n70A
BD1zmyPuFxARI8g4TB1miNklIOXyCLDuLfGM442kfCJnhiVUc9SoZJSE8sLL8DNV
WCblh2CioMM7C0T52XLWacDuUBZqD9cwjCQe6sqL3LOWyRb2pLAxy/AqqFH6yeKW
WlqzMUrqNBUNu2vb55tFv7Qn9x801Dt7L+liBk9VjzpvdPm9UmFNOe2niLbJ9glf
OqpbzErwsqRq8DPfucUeBbIO8Q8Bp3bGwqn7qdGH9be7xQDU6cp8lZmoR7Npm8aL
RHxEQ9QsYp+ygtUplE2QHeMq1ZqBsPWFHnTUHWGzSCAylt6hVgQa9VoV7Kpqmjyg
dTwZTj7uq0idazCeJQxwlzIdpAr8+VFYRQlLrWrfoWODpLvj/Y2tqws9H+5/wWOk
L7S/ktP5Exm1oeq3qqadrqco2D87tZa8Ms2i0gTCPsg4IILXIlH040uksKbRfMfz
ALjz5c6f0r2CSa0u7YJg5qy7STSGdjM3Kgz/8P71EOhsIFSn6Dd6K8BsDSYSL3ig
+ngptUCG+F1QvfCeGtm9K8cMZCucmm8wGafHgT35g/Rln9KiEeyo2bbBTwMLYKKs
iYbmfW0thHeNDUyOlt8/DcTHkkm32Hvvi5GyAjpcRynWuzulAVxZ6CDg9y/80jrj
Yog5Gpz6fsy6xQWMm2MP6eMchxrxzGKvfyuNOaYzJZUKzPQdwpHehiJo0zDbMOBV
g8zET97tp2wcgeN49ZWWagTev8iCdGzfy358NvnglHjOS9O+5BFruvNVVZwYAlbX
J40UBhY3DVEdMmF6/cygY2aq5U8ZcKlpYCOuz6+xHCwJ9hQxoa6oZ8VaZHKTGljU
suxh0nLrip5r1g5LFFuHJAtOWjKRXzfSvBGWOEAU0g5Cgh9aEA1OfHUevKqzuca0
eRrD7xhpbPG/VGmLhc44oKqwpVrkUkeWmF6MuwGd1vxQHv9zBQtQWnpOYlzNMLWD
KLL9IWFQeJRUCsUqwqLkbU0h5KYUdH/Fza2PGVvcYkYCifMSXFldfPmm/brB+yRc
oDKQWro95mzb+2oXIB3CYgDT4RfIWRfdbWEpIgFboRtqckoQ+CogvCRHzSKZvpq0
Dw9ouU4AJDpFUWczVnHzJiLNgehXG9Ni0phSzTSdqsQa/T7wGHBvbdrbOUbB8ReV
Vp6VT6F1J6sbZACkPzqOObrZ5TTbSJfHuIdubG/UDQfTTNWEILCitrY3IzkcvQ5X
ztbNrFKk0IAxRhSfkxOOnMNRi+yuFX15j6NIlim8yfpJcTBlXVfeL4XwT8dBkdNj
oUOGmbaEBDmgfpTT1myKxjMaE+9kIAP/4s4LUUsurEeVLiTSZQUrTAhhqb6uE04a
LnpQD/QC4/HwzU525vklk9EVCT2GqjGYKzanW1q8rkyNyW6uFTRwrySLEY6J/pKt
G/92DXmxzdzfHKt8isdqVhR/tFbRhxJcBLsfNi7M0DY0ZTgiWKJc1VH/tktN2BDO
Mm+BM7B2PusTUXdLmOHHAKiXC0eY3aTGLm48aaPFCmiWizarwKLl1Asg5kF40VLe
sdfhftcT1pW8oiAY+Um/65pgpxzXzlrNykYofnKdf0DZN7zncUxG04V+78R9tJ9P
99YTt/+vO66iTtvuHgdfr9Y+zxS+M0X1SO3mDTRtjgtPOIqqw+gRmH5rM8o6+kKH
Nti5vBDzA1Ns98/GyievSlAj+u3IB7UWok0K0Qn/XWbwD9eEBOnMiJjZLfBMlmkO
3WOWNTLmv2iD2XWQM9NpiFed6ZArVTqxLCD9qrkV7o+KgKrRhfJHVCH1mP1gaVuX
jjmlmuGP8OrHV9SI0CqKD9OL25sZoMTQeRs2l63FbHQXUjJ+9ayKO0NB5/tsooEJ
/uzVtPlcSGQDINHICCHEZ81MaiP6AA3J7wSwO095zJGDE15soMh3b9wSN+rRz7D4
oM9zJtci76zrGj6PftIc4e/llqKj8t/lZ+imaHXFWj7ESrbJnvfKEyIIjX2ZliSK
H6h13XJPgYYl/ezHIcnSM4JoSDvnl7YcLgfA/TgvFdfb9Axr199FE8f0CEcBGNoj
afJm9LWQufFAMphHPK3BmWsilbANmTNMENz8LechpVTDEIHtAg17m3O8HbFBi5DG
MDe9MNKPDv2de10Xo+zn7YLcznJwXZx6PuEdxaTEBaGA+6yBvERGzOuWUBJ1mSaQ
voA3YrQ9HoHN7nmG7rESDDCvQZMfZmaUT7Bn4ImxiJmwF7OecASsG0wA0L1fM2CY
JMZd/v5VqDgwTrNinBd79PgHfKiQGs4UdrDsCL5RTRa60yFCXpAtGz3XXUgr8GsQ
l+vcEsh8A/Hvs3kK+mOYzQul2X1TJSQaS1qmpzjYwYxPJyTDTtDmvIlpK7ekBN4J
Y4h3Lp79cMFRL266RGKivo9KEUHBcZCesEqaffoV97FrZCv+7SMXm+1V59+hYp74
XOzn/H1omq/vVNS6sOmqm6F/ngEj93bHKu2PLTa5GjWjGtekGGRqZ7oip5nae5IP
bGea4J5NzaxIJ653WMx83GN1zdMcfOdKa54od3eInSjGRf2JjhOAEEo0hthbHaFf
W61qJq3N4tGIKNvR9P3RJsvnmZgWOFxKa5n53HAhD/CGDbkmTy/4GXixH0fAaDeP
/orysPLVC2snkBUhseZuK0BysVMfiAniNyOAKBe66kS5qqmo7UWMuO0ezEEaE11A
hXvb29l3B50uK6GvpXI2UkRMOfOqykA3mtYtyEckCLtY6eHLTVQ0ouobSkC8/pkl
knXwCs5UJrLDURLszmF/B5rArqJbiOPgIzGGzu3OPTnkctaBC3+c/W/4iwzb9Y1x
jamJmGHVdbMQXjHK6HuDCg7IBY0Y+hbYz2IKkCqF39xea5kOhclDvto0S2ewvoiT
1jiGSzqAnj2ZXqikBO8jj8KCiJTU8EBEzTPy38S9bFxQN+ICkKwZNRFiaXcrfqB5
v1jpz3ZaMKqq6XCHG4yKfQoXTkeztZ42QOK/shpBidPMyEpLfkbgFYXY4ze/Flnj
jMET5I3pkbeu2ytZYNh9avEPSuQ+QTqblvd2eiXLvN2azPYMItEI+rbDgvpMqd6h
7RnUEIswsCQOvl9wqAd+D5XgDv6gDHXP5w+ew4EQ20A46PRXGju4bvaSjFp64b5H
75oB/V6YiAwYx6jJngeebc7y1ezzYVBor1ZSf3kJX1W9pMO2zSA+8BCAtvXHOcsB
+Xnx33QdxJDXxApFSJEnFvLrXHzElZgCpBdCMWrpc0/zDYIiyQaTBCuk9TsljHrY
LDYP3067N7/FBTVM4m2qebUwaFF8aNclB6UG7P2SyAvOmGeu1g37Fe8RB1/wTl4m
3d0s6jkZu+wvMTYy+xfX+gcWI/BcbOOZQyF2nxUPyAL9ZKSN8B0XsshpETDlEXvm
8mTZfbnLBNpBuzr2yDpKRH+hdp44Y1eIV/XAJn93wAJt1VhNM6E8y3JMHpYrIdmd
b9YWkJrvKywa6n+/84Qgxs2L6x0SLotsNzKCGOFwNIod5mSpiNlfsnDvzFgDsI6J
Ef7SkpttRPnPuSZW/YlBgVj6v9s0XFr09eeXia83EoffyG/lx80qD3s8RAlN0M9Q
KaLIh15vAXTRyy2rAs+S4W1c7blfDdinnzhxacsdos3Wcskv8En53Rol1ukkE+J3
1auBiW1q1I+HR+iCwrGPTZfdmHJz5l4Q4Fz4cPIVErRzTedvh8JzlYi/z+YW5Is+
b4QxP5ipea7FTQrSKyHIhcDTGtIaazVG0hEBKjl52EC5Ov4IFwejz+kiABdPjcZb
sHwSYDngBZZL9i2YkFAsHjmRnSmdKE5wkn141Q0vSh8Eqt5Iv0fJj22a07uL43YM
qS6vAJ0EVNeRftt4n+AfocFnhn1ipW2rASqngVIZhe+ffHN3280kKFbkk8wt4YR/
gvG0OOsk9IPBhpea5HUlbaA5GLG1dOLpUAxSHx0oHOMau+jxIzbOsHl8hUZNEkWR
IsGU2HovSAdmGFfVyjWsN9EwpJsJHdcMwEkw5yLaqex566D5OfHV8LYPPk2kTIYG
QwpXaaq7tZkMNBfN3/npdzj9DZeyL4u+F2APhnPWhel0K7L0C2aqr0iiN+ZMcN7W
mgUs9DBi4pmjn/OiZCKP4m/FOonva5o8pfKns+WKvdHfL9h9gubE0z/eMxdF4f2p
k0LlQ89okC2Uirwx3r2p9asyzxLUZGmlI0oyOt0ZH+0VvJyxEvrugM4zd86j1MyP
GR+3QkYpJ+y8H0OXHgCJY1+9z/fnQncdOuxQq2QRW9ShnKkwAuzBdWLGLwpFy0j7
qBCI21omJwPprdFwAWNQlTl2KM+jbi1SUIwVkEYDBEZQDWjuQ7yt/h0fsr+6reZP
E0XfmsO+CQwfjUy+AdDFIyQdzPQPzYbMKy4cqj1/QDIFZdy6XzEIrJKGQxoOKdVe
g6Pddns8pMlsAvKWiLGj3yvGA9LVETgUSVCodrO8dBG8eNNzTLu3syYjdfIBzdui
RvFYUm5FFPEapzknmq1IFymMfNb9MpxnForLNTwbIj8f+NlLBSRtbry6W4QATzjI
Z9uUaxXrlutVwZF8ImPW/7CcH0995J3NhycXg9bDVeKmWEZp2fwOjr35Mztw4bGq
3QNPz1usPSmpgv8cNukmiqdQPEB1ybE8G8u7+aSkbVarc9XRFyEmNLzjKZo1PXOR
BlW3MKkNFJ/SyK2sOjAVDYhKMDAXaHila5JXOrsv3SihwuAkYzAEMySG4qUnkiGh
lFtwnzscj2Zz0aLT72tvWoOIG07YQX9Rqduc0xvmTg3jHR+z/9wXPQIl7i4vAjLl
KdEvZsh38JYe3SHBUTOIJeq9yT1St6XzE6hlXwoaRLwQHM7JPeenQYVcxPruVicc
eBOn4YDdSS+NQyP6XZDk6pw6etOpl0I/Tzv9sxwxnppsygfPhTo7KJLH8yNwykNO
jkbLJnVMwC7IulAWq5F+gR/g9BJNfYKQm9w95EdrS7niLkzr40J9rufT2FdHqdqQ
NcFYl4XxUoBmC2pW7JEgMEF2AHfdzAZF/fsZkAzJ75/pcPfrG2tcuwgddUjo7cTw
rKLPWl5Dd3ZpkjdeFe9v36mFxZYqNiOVh8xkxx3E14gbgLl1EmgSLxBE4W56JdAV
EpeDyZizu9UDsV3+Ix8B5ZaX1/iMAJEEnSIoBIru1sze/yCvd5xwNk8tfhrOrNxl
3ev3pxMBMHljfzSX3UjgnryzjfGbXiQpTMzKUPNvrCvin1FzonIzZau/QYUKzLVo
fFOYJ8xSA6JjhhQKVxMa7tsObvqDg5VyXCorq8aO/DwiaYVzQHoGlQ9jTyhaJgxh
nuTDq4we9o4NGW8GULQwdIDiGFJ5Ki3R6tZrptB1lENm1RWI15jJCYAPJ+qVfS9+
yREaaQKM51+tSm0lqmRUC9uVe14ml+cbHHNLe2ltdihN13NqsLMILwfrICzYIwid
DfDCTHTykZtLZGPaRqewXuZhjNJ3M6RS6UpiFYEp571+Dqhu5g1ZNiDwqG/sQpw7
TlpTRRLATyptkuD0DIuogzTepLw9vRjSb3K7s1GYLmBdfWb06n/0gAoZce/vW5Re
fm6CzSvpGIloPsuNmxWdgR7t9TsDIE7NRW7zn5Mp3gBPGSQuhimjrSlCvmYAOslg
JDoQN2X12ehPMvYm/Qkkg5JKzkuAiWei4fKmoyDO32fuG4N4KpQZIqk8d9OvuLDc
wNZoc8qyy1Kx1OZqm56Ir805SdLwRFKD4cDvNRg6/DEKrIefMT/Ujc2Nncy9CCZ/
LDM1Bj3tTyTGNLLESMPun9uvEiokihbN43J1OsbDyDJ1dG3tyNeqC3qK8rcZUFWp
ZVhwYqdu8rt9e89Ay/f644aNzxOu2mL5SSnHCk/JOOkUXpoOsCbBr6KC2rc4JASJ
0woMP4hyFD0pmKM0qdmWtz4Pj9ehyM4dpUMKdc4Wfv74u/TPRGXlxqtzlPrrXYiu
MszcyscGnv4aKIHXRqmLa0YaPSPvMcW0MWBxyXa86ncf4oqtDJZqujAj/J8TifFE
IgRgXLvurRX1KjnhtBHWkhwzMjF7dVSG9dYhZXP3f9O603xXSrIiyQONFpk+k2Uu
+66drg5o4pqnkEngZmMISu0C6FfTg6EHKBv9QR2l+gFCmsjDgAjXnm4ECh2/JLE0
uzRApELm6ayTvCfAeAaiv+wQFJj/hIKg81zgj5+erTvS93CjTQcFKadBMnD7M+7O
yxtjA+Ode67adAE8JdMDnCjx4Sqbw0P4USHO0sYbtPgZUAsNVvTkusaSE43DZn1R
Aql86+8I52OACfVrxXcWptbXm8KWqkIIwZsElTiHop7pUExuZSbVTGB4mdgiRPPv
h8Zo3i0Ypq615VIKaxF+00mBBNjrpNHp2l17ehbQvCB9kOSZfT6odP+9Mtm/47b2
SdEWeG9mzpo+h6Q7d7D+z64W4JgZ7bTeavIycD12b0mQxfZ4bMDb3NI1Kr2E3vxZ
VAt70MxxCt6agsRJJuPpwE+7FtZGMmZP6hUArdFvSD4a+jkbKKQReRLOSPV/sHAc
VAzPqX+cn6KzlluH3rvE47vXuTUsxKvkM6SpnKJYgReJId7tx+K18z26z5Nacor5
emTJxH1vYtH2H+57z64P5b4WenAiMGDq7mPcclAVk02U3NhyBUQ+w7GfSNnn/KGu
358562DBnTncYwEerOOfX5Af5pJmQ/q7gKYNFrh16O4PDvgSG2I9XS6G9gYp+d72
dxyhFvUw3Yfqh6MgtjqRS4j7W9f/Jxizk3vRVia7glci/GEqrY8qj53jgbNYaFf/
9OF9QGzbiRAbAGPNswSWtbAy7trY++cxjpjAsLU8LtWEEr4D54Ot5uWeVkK54yC2
gAR62Npa+QAy/RUHy8WDl52fyXUKm7t1G9IMc1Il6GtNkOOuq7vlqjxz5ALrik6Q
VnQMEeOItM1Py6L44cbpLq4CLscuQqYfiBvsBq1zkWkm5IJ0zXoxxECS6CYMUEYc
aRUyxXzItnT7We/80RAG14mO55PGQjHVDdF3su7yX+xZQkOJjBas3gOklRO8isZd
+EO2jmYlX0reWW3ynzI1vkbAOct6VbTPtOO2vuQgH6hRRKb/ksZeezli0lhbE38g
bQ+lWDSRmoW0ZSGNzS4Dpe+e7nJh2LjPgt0Bq6+kwCjYzwk9muS/6eMeK7yoKgB1
hR18w2nN4RVHh87XFVm2D3S8cHogw6i1kObSQfaPTWpauajJ24dZ9ZLownTsAimJ
O98Ungm2rbtRs67ru8D33DbXy0ZlzjVLM6+kgyl0GqgpmI+IOPDeRlmHlr4RLLVk
yx8/Dy2qCZe9VUVCe9mBqPbgPx43ynO5JpTw2tKDagxk3RWys5XP7IMiGosDCuU6
RcLLN6rU2cGYzcxoo30qG+IoRh02Bhd658KDSijwFfBwT5cyEbQLtgdBcNree6Ut
7+z7sDw0AW8RliY5XApwJ2s25qQ3Z+cBoTBT6SDUCV8dCykavMtoRt0xDqFPyqkm
4bTMchOSdRm0ItVRsnNMy3DYSFKOxZCdyczq1+P6kKk4Ct/vyZdN1vs0Zz8JHyeM
skLqhmxjHlmdhmAeXGAMsW/1AjNuZzgxxAQoA6JiKSxs2dHAyWIe5Wf6TBhC1T0p
gYge2c4zrxF+dU5TME8HPB3EFCy7oep5B9VR1AC/3+f7yfXKDJPFMzWE7Ap11VDi
isn3EHXjQm1IQtu9fRKyUdZ9byV6Vz4UAFTGjPCuve6nSAH/mYncj89gy80sDrRd
szDcK1a7oWMUk2xROW0+7S9uYGazH0jLpTLN2qR9IkqzeDddj6Y8AU6Mp2P+CAJf
hg668xBVl6u2ojJ1PT60E+gq9ImyCGZH3U0sZOssWoA3/RgWABKEBJIaF5BW1y9y
mVdwL3XQdtAn4WFEbcKciX98yogKr8pTWBn8lSjySDJr/p/EajEhrlvhspF7/6D5
AUSJEpWF4qBFb/26Bz5mTPVLqbPhp58L7ENuzBMqlQiEjIxSI/in/0PbNbvGXVtz
QQtXc5Zr5+HwbgK31BT96s5Ox/oc9cH0gF7mSkUPx6nYA99Z2bKTE4aUL1nFJWqT
5MieIDh4Jdd6QQgP3d6wfBqeY3N8M4TWU6XdvSMslX12MlEX0shnvljgapmTaMKe
DA4cc9PMbjCENL1f2WvkUujgb+GPmtwd02WK0fLx3j6zS3NAxGDFX7cVcLFhs5wE
4myHzXpoH+yZ+XsPec5SiSoCtdBkY0tJA6/o4PoWleFrB80cJv7GVcACTmfBueL7
y/Z3ZpkCBe44H5guKqcdiUTiiy5in0n4ZmjQgS9x62wPGBUOtuj/Rf/IJ0iVitn9
nDKDO8AwNv2e8k4KUB/jSf0P9AEoyIwYGikNmGHJar4ZFWTglYnaxSPJM1ne0aeN
r6XEN0lMJ0jNLkdsn6buHVCeFLov3AGLIQ2wEjtCWJK0ygUYflqQG7ET1OwWr+Ez
g4rH2O+wOL2cjl/LzU1xKjxJ21NIm0w38dv9caJVtoQiXVcrg4JE590EjMxTthnI
eAToH9d+mqdlmJ1zrwjCUVV2wRl1FUEdZ/9mClJeMynfOlRZVV82o8uSU81UZ9i8
hkNywdR/a/a8BVPNZrEYM5ZsibltSudxNZTD9VNabNMbSynIAFtTcqig/EKlUHr+
vFuLgZYxsMX3GT0Dsm7RMIpmOuGcpyHg9meHioel5dRlo2nb21jowaAr3WMgrjk7
4YFOK8tCfMbT5qawBG/WcVfTUs6cBIQt83wWmGsBMTrjYCtwK068oEtMU7e/6sQU
SxMiNb5cX5zEqC1TTY7b/AgQYVQBdJ2uuB9kswpnvQ4TMC2dbJnBs+XDUkAiHyWH
meh27M95Hj3Wo2/AgZPSFgFSST8OboEt5eFGfIuL14iPGoCQ26cpXey7wfo1LVpB
unwpEQtsbgraxIlAn/YWGagyqMQIGMwvlaOv7IafFf6ZvJEXev9CU5d7UzAP+ITw
L7L/vD5+SI5t9zNB+TM7UbwNtJmXzTCuG9JLmuX0ip+rMjTGdfgoQOq1tLv5BBmX
/XBoOs+I/HlwHak709xC2Hs7TeseRaEeZgM8b3+J9oXqMjUMdVE1eM3VzbFvZOnI
HyNUJB3Ug4m8Qo6j8JejT5wU1xLk1x/74olylFyCWnhE7U8lj32kOqENKJQxJkQW
0D1plpZvy7jlp6T8EZWe1FVpg+JO6eXBYeHf4YPZLyoxUymSkofUtJLUi9I+0Hdu
aLk2KDajw3yslx2KEQ0SS1ZIT0tAFIS3jOAIbdtNuB41ieqM2fDqxWiFtBvQwz7/
mb8s1b5lSbJ6ss/4LtM0IQScYcRzKDZFBdzbMjMRWLPAXEOnVUMLDzQaOysocLWQ
u57devZqIjKapRg/OXpwJlBqOoJy1wYbjHcRY2j5+uWRO0rBQ1+tqE3To/GF7iRb
eAA5mQLeNuQSxDEx8to7fvKOv0qQTTA1yfXXR3xlqQ9s+2QpmTsjoda2s0xRI75e
5lNZMmDoQZtgwMPBcfTVW8lVPA1sFrQne4MjzRgRNFev+JfvXsj4jIeTbNxeVZJo
8lNW5nZ7+gArTZN4ma3x48dlJ2NN3L1KoVYIUpb9hNWQfmNUtHoFy2EAdjteZGmR
ls3SfM9OhlgQEKxFxSieQaWE0U38K0mjfdY74CATodY4zr/EUTPub4tbZAGe005x
uia+BrF7AiWVaqDlRV+rZoRmH8j7L5NZGy11X0oEQGi0Xelm9gv3ZIec+K/hdXU+
YnOyMgCZNI5pd1siQsOiMi6KZx2oEWvaVju7gasefl3qZ0bGokW0SBKl+lBnH4qE
KCTDVdGx4011XtdorqN1CEusn5gu5wE7dmVpd0f1f3tlXld9VErO1w8WfIQdmznp
SYmzPHtxr6tawiapNAVoeSYC7FlgEomHqMhHTtw8ymQjRsNtq+QtyDqxau5BquoC
WJrqLQbwNCbRtp9hU7a0wmPa9PnHynB6kE2hvFkBZOu3nmIL2GLPeOBQLmWdlxe6
cENOmSieVsEh7/Uuv1vD1aZj1qh5bulfjy++/e8LdiiWG5UPsXf/sft4KWM6zmos
Nj7s3msG4qrho4a5EgwhqDbELhJe59Y6yJLfrjG8o86SVZiYtFJvnCQVNGqCiovG
0ujlnamOwlo7t4nq0GVDmn5B6dAXbvWAXaIg1HO0viMtDAahlIEnlwOW/+fmgXct
ndhYJknTJaFOtVf2niHYoA1EfQONTYgzwl3l+r5NMkqB9kh3q/9OH8aheA6ZFB48
KsionISdnCFEV23pazoVKWigs54vq/4MpP3lT1SMBcmHRIgtB5yeiMh4LSJs3OZ0
n5eFJ4XqVFZ+F3gUeTVUWdcRiyhX6kjrcmhsx3k0UxexEOBRZSSG5L23Ow5HFLSs
IKHtPcoHLMwFEBgEOlsYYCCQ/5vsGRGxxQr+zv/L3jqxWX+mnyy9wumfW7k84n8R
u8yQpEddKTua+nW3IC/ROMsv7Ki07XAKkfWxr4++ZsuvDu0GaXOj2Bo1IDJGTTDr
lu3EVfcQBbUAPU5zLW+gLVCzWBwiIbVD8d8wwvQIc3yE2CaqM1KTIkuEYKDJvmP1
VC66as+lpoTnLRXDnJ9bphEYXGV74TDBGTglnRIBjxeZqTy7Ppl4ZGjUU3daNjW+
Wk0iZO/XVNXJfVAChbMgUUrHAObArR5n/RrXYQADE6tUP++hiKbrLNGJf7eGPOVs
3xjzs5L7mRuHtVCaMzDqEoQRWIEI4G5Zf8QuJbT9l/6qDWM9S0c5Lza5posS3vpo
aVz67xQni8zV16R6FAYWh+9dnos8aGmQrdrhMewBq9SSSco5hSpwRnxiBOZc9lxK
ct4ECuEsRtIn9g2odzyAISJXudDditefx4zQle4NsJSXGUH7B30k4X/3Zvg9Ftd8
x12pk/08oP5bE86N+kjoZmJjZML1heaLgfbFzBkalXEkdkIrOWY6IP2Xmb5mBaTN
AlpHEn6keK3bEs6TMhEawJzsHkVt1m6Cvo+35xWDAh848/97zVT7VuF0MUQYtgvO
XUr9Qkf6Bsn5DMwFethmLbEgjyXc+IuQ4mpYnZbDG1uERwhx0cd13awcQAMMxW+4
sSrdfeXPd6mq1ugCFR4lbjN6ZSWc0NDSFPfA827MHUm5kdHNvN/Zbi8hObwAdYEA
2y+uwvyvdTh3lubL6sf200tzDwZQNK5WgbbMVBhun7pWxWWIAQxa6lnYV4A33Js+
O83XVeQA3ZpKtGLe5qoya1vciIKzZKddPcfi9A67Xg/0RPfSVW626fvQjs088ZGl
DAa2fgK53Lo4B/T4PZqETSjCpUAQ4EYW4uadqXeKkCgky3ZlgkZbgAOF6ibomO2L
ZP373xLzYS9sw/gSXNDPc1FbZ4pw9ghHOt13KGJKYxevfR52Z1vwRlt1XUSvAR3+
qmwVToL1hB4RAUhRTBMfogYDTAEm28OTJbIgRuUn3kMw0EvR2S8Z/rDK9ABsU+7z
fwHBp6XNTkaHYwcwCbfEoOnHc+8cgzl9UxHQl8MjT3CxsqaFFvBRjW0j0hz+/7r+
EZzrUPMreUokxJkyY48xJjGR8XgjSAVORhxTZmTHyXWhcx0aLY+j95XBn5UM2PsK
/2DoOZ4skrbkGwu4RyO3Wr5wUE1v4GvOdtQ9Z4xfSvMKv/xm+65hJjtax3sRo59H
x092nKG06P5RNLoQ0tQnGxUuWpYCJx8oQk+hGVkXgwSvGD+QWf4LE/uZEakRX30Z
4maROnia2/aCXW39OzrWKEejGAmWXS1BbLbejdnIeSkKg2LC++13F7AnpVTjRjBQ
hX1Xa5qBXQsC6Yv5Rz9FAXxBB1Y1xxfP2UWUou+R6PmcyhznOnQ0bq8XkUg7KXim
VXGlH+uRXA9E2TkUlo/VMpJBBgARbZJkzFHDCf0H7jW4Mqn79rIhDUa/sjxIFHDQ
XyXSLoDWktN7DKiUUPg9s4be9niel+L6yFEOYOCEeH3v1VPls5csXDDHfaXXAUu3
xCSFxaMSnPF0js5566HCOqMnKicGjN/wVHS5ee7+1rbxzsM6eBbQt011Z1nOlPxF
ZY6uxbZQYXFtdx4qxc3HtTyziTJQTN4S5f5AY8vUJr8AjYExasbr6Jaw3Q5IHaTG
lHxxiQJA0k8yjDGp7TV9wCvX3rNwJb5pEAWKlSJ9jnd/F2k82sTr/m+LdrOOkJ5R
WJsMKTDQw5T2BbpgpY7+caXpC4I88ZW/9fMQfoq2pUyv9NP03f1c73/jrevnKF05
IIkfu92zL25C/3nEbuBoR9D5SUNgmrz3BaYOy/xvXSU3KEWp/Jcr2wcoG+OMlG/+
5gSeu1tX1raGQ8KVsPVqyEAuCof5MS4FiLuCL97tneTz0Qf+F4lFqkUOh/vGJgoC
FTNryL3cZjHkwe1fPdPE2lsbFaPA59aA1qod6jQcMk2Wu/TOHcyt6fQw7u9AyF86
s2/6Ub23LT0x2ujeql6UkuhXQEWMB94o3O89lpbJYk3kVai6V0l9uyS7z49lZXV8
rBBbbs8lVNs8lVDdSiALCDQNsFFhfg7ZoMNh1k5wYfOV6t0SEif6OH6iqc7hWvPa
DtN5d8rhWMVMkzXImp5fLZGWUqYIeCS6c0NZ7RdkyD9ULGIB82f+mLVKwOt8QnfT
Law8N9S4laxs8NBUYfT0WB1F4HxuTrRpGZ1VkCDJaj+brxoQ8MwpITe3aA/6Er6B
FtPsLt9SamtjkdadXXtJnUP3M3X6YIP9Pf2roPsJj/SQkZZ9TIlvTu+0AONQaBYd
azK74H+Tbm7vex9RJB/r87ObzKysW/grJmQ1NQ2KLpaG37swIOdfEghkIpPlklwl
FWFrLXgtHHAE25zyhw8vcQNmdYCkwsLHI+o+FBWoORpR95rt2G8Ay2s6YF9PN7kO
mJKDw5yofCWzZXkQjSqYC9sPqZI9+z7iY4uyJUjNV6E2BTjUwfWfu1P9xvVdnJLu
h/4qsdBH0ylbJELvHbedB+v4qnPvDKc4C3IurSHevoSH+RVaMXsGJqYhUvirljav
Nv5RxbXeoMwkCLkAAhCa4DDnQWUK9irSWTNTMkZEkZs5cq7VW+boIDD9JB9oJb3K
eS4XcBQbHu87j5qFaD/ENn1Bhm/xMS9q06ncFRqj8qKCa3H2SgQ0+NBzcfIMliU9
1SkcFqxJsQS7zmu98txbuDYBPk/zeWrLdwwxNtOZNNxA1pZU+rPE5IUBFKQ/4tRb
ib89VvQoUjPhRLSJ0kZkPMiXQNY8LV2P8Y5XdcvxBTXg6orPZytMMGR4ykDLT6PH
tYfHjY2J99hBr72fdP4WOuQU+AN9Gw5aNdkc1nPyu/Fdp1MpQxwW6BOwoDfcIepo
YQrzKjX307l+yeRuHyLgL6uL67zqZqF6pgqBKeqYZHkH0Q7/UIgrzldXolL0O0sc
Tp/mc1x6l474QadJY5bvdA5mMkY8qhrqymvY8oXSpHX6TUOXQrCMzOaIYElekuro
kXfCcNfWRtbGjxzuOHSm1ca9HaTDR0qUw5jgdP7i07ea3yUD8A4iw5QMqST2qJle
0wH8hieDOfyRvcw5LtK9dCIGJGZDwmwhiifK6LF+RqxBDSATz4ppCbuWXNMhKwSh
RKsD7NTi1mFWhNY7XT18kEh1sJDJ3ukBYYRn5KtdF4ej90UqrOjLTsciXnEwhZb9
gFwxGlwern8vxAa8ppN4ZkDN9nbx1Co63FwIn750LtfI4glreitZivt/MXHWf6c/
Na7hfKi/X3cIFYuz5K3PuZ1NufSP4kmmvTNCjzdRJ3kp8VobDH49A4Z4uLH2GB77
bH+iiHXgWCpRETjNLqy40lKItC/iAV8CHZQRaEN3bbAekHcQJMza171lvB+hqrfv
crjD0U/SWZywlbGNR33+HXu06jWkzfpdg+UpViNp7wj08M8Y/ybsSYwDX+s6mS1a
F8+kwVzH/aCTxu2XtFDxsRDTjLiZuNmYYT/Js3oRQ0bysmxcMtnDFK7V+pgiWL0T
qi/e9c+RGJNqGAhvARB0+EtL31tqLAH/uii4woeLSt7CNK03iA6PxKE7xfQG8+TY
ZynUTygOsplD8CHVrSv/FfLXwoKKUAChqEUwkAoF8GLTBXvvcnj4YeFRb1ji1Z5e
3lTjcAIGEy63Xxyt4rHp5A452+BPj0UfeHwSURlwNawdKWm0zyN9H+Xh2HfL9i50
0VqgvUSMB79fvLApiguM7PpMancOcDo3pDYcavTm7CKQrW7AGtEZnmL9x1v5BVc7
pfV2zvC48H9uiickclOTdm/Y1EszVj2Cfyt9YGPZoU3p0MNBOzfoyqV5lwDL5Mrm
xU+xkKu2KBMvOzsRckhixRtVNHB7l/GuR8RQyx5TYVM9Y4Brp0/CSVfQszfZJe5s
OgxRO6QBeLCTQyj1M9bN7XdVZ8YtPYMDZ9vBA0IiCaRafV1sy5N/0fYJ3JY4fOjx
LZGKtvm8Ah/L2+IWt+tzDgRWZCtb9+WG8qGKF1nWiLgL7BzywPoO91HlvsrhIFAc
mtn8+aPOa+JdQFUw7SV2o7TfX7uA6OWRxIl0bdta2Zm6wMddjPylwo7TQL4SRg7s
45/awSd3JEprFf4z4Lv8ZBOhO/xIk8zjyrFYZDZ2ZNcJecK57P/mKkUFwbD/wusw
Crr2uOUnvFYLAkrC9La4Cgs1Je30Y0STTDajHGlmf6e+1BE2tjWs4CKmvF4pgK/m
p1DbsT7qt8Nf50heBwmF2SnlvFDca4VqP7TBoS5i1qDrToxwwxGnumEMjHD80QMD
k9U4LSAJCdfSWJ7o/9j+SvEcCQhVY6tmY9206Gl5JkBK2Ky79BOWakug4hsI7yK/
zb7qwpJjUhBIL8BCj6JCSbzMqSMCWpdzd5nmBgmdxocka4ETZ8kXy0aqRKSNi3/P
q3jo3VvQwz1lYGpkxhZBa2lIpsAHHlzX3sKUuHiAtgfRmW4dSCm1GMIRsaJKyfYJ
Q7PUARiE5C2+vAR5H6xEqOeIpB1rOQi0YFE7DZBikQzoe8JrRve0eM2YGdl0KQHp
QB+WvDhkUayWP1Fz3ZXzqH7kQnWUpWHl/g66rjYJW6CWHSOoz7HySc5HRcldY4Gk
PoDSM1+OThv1ShPvxmKQeQOSzlUrknwNmllZccywzleSpssBrAMvA0LKd/ctAnZv
c3t/geLhJ7qrD2m2XiNnvhu+Un1fTtIXsQOV1dqkunnUxE0McyDmYQNwTV/xfaR3
udR0rY5OHeboQ2AsV4DU8b2ORcsM8xtnDU5RcdIWDa1ho3hDPTsobU2mCVuTafRi
T2h2ge42Llyfr2RQHhTeEWMhw0TkloYRqBqYrGBZyVJ9XXEgcTtzMcU0y5HMafUn
47x0aW/0BHu5COV8VVL8HZJd5QqekdvqrzXeYd8p2jZuOveRURzyr8qNunfJd7aq
q4wtYhjHe0l7lYHx15eiRYW1kKvAwPhpZvB59qwe3rfPasaeo0qZfY4MoIAF49aD
oFWAFWsqrNafZL8jJ+GCeI/53hMyceBl6Uxv2bCwTvQ2NVH5xQ44IyfibB2YLzh8
FXHJSKAHRPgzHTUwy76cJi1oDBLRg4ZdLdrMePj0SXIq2diiDDafxel0q7beavpC
JPrZLE5WnfeBWZhDi/5+rVrxLgfmbK/3aMRl/B9sw7bDwzvIMXaBVeqlxfTcnZLQ
9cZCIhUaaSbASh+dBqbiGHW5OPVZrO816MQi/PGWTCZ3rmWs5NrgJxOCmIEhULhe
0n3WsLvXqG3ajLrKiK13rQwZqFN91UG5coU2dRRBNsgkUul1mS0WBKPsfKda8yrb
OAunI836Agp2RyCZxZfvWUq3kzLasHxo3peckMuQnqr3QMa1eEA0xv+v7hpR3Lcp
sWehH1q72Gt5lQc/pAmpcECNBkUYOPUe8pWW+tN+OHswLu4pg5U7ENBt+CY+pzHl
wW+cG+Lm/aMbpM78pSCfN/2O7ROdLJWHjELjEaVFfRhkB+1t1uQjHyYw1+o2gaq1
UFiUD8ykUnUtjrZnzdKeh2wNoKeU/UobCl+VQbZ31nYNGo9Z5q+3KoBnUfPHXn2n
7h/c8T2ah/Xey8Us6/pyIBDAslj7nFu2RkuHZ0pZQ4d/3h8E0+/0u3udJSOfQpfw
ilanNqrwxxPUvBvDqN16HbdYqPxiOU828PzaFvue3KhrhryHYz67k6xvjO/4flxj
XX/vQ7d9qCiJs3QYt1WEjhyyAb/ZKnllGe7+2QIriQcRMRIbHU0keZIOEXO3LhAz
lDJMhLiVBz65g/j8DTQTdWbeJWeyW24ERefrAseDKtYKA8x7ur0A65peQgIeJvqF
EanmkeK3pJ3xSy8ao56/ygkvP4Mgt06hqI6JWoVLrgc9LIKJ8sLfl7Em0Dighvn1
AanBfKIg2cw0dcw1iS5if+b9CcjNz1s8xY6Din2sjuAmkUETm2mJtznGX4qvzt72
dOvluF+9wFCkoOV6swms+dUfHWA5gVkEoG43RDy1p1CyRFJU/uJy/+ZK2BMjYP5U
MB+4p8B9OmTAK6WiNi6h3jikKGeeoROof4hfKIdbNRf9q7GEAWYZ2OOTsXPYrgmI
A/+chcOy1M/Vjs9lxdraRWXT4jE50aC4KqDrKTXrfy7ufm7lLMKDCsI9CT7sm9GF
hvKDDwrJuA6XMB43chFnPOXc2jswVvS51kVOawPUQEko+qs0SA1esUdRH94epaIF
uRPLaNlQCJANaRs4PmuqmPlhqg4CXl7ULn4yIdkiEkpTtQt0JqRMQeHrsUC4MJvA
V1EZ+awb74yYOf8srGz0i7xit+ia9DxVSXxqhsbN1M9f324X1BHsqi/R20HXMPjI
gouDEK5KCCRHH3M7HfqLyvlwyuc/A+bTlr3jrDwBmC8aKkUKL4fE+U+bh3trtQlz
8zqt5JFjKN1IUYzrHTUS1NZ39SNiTlWvrQrwrIMWDhg2JYEh0tXmLx4/q0tf7ucU
QgBR9kicpr300oAHlT7Q5zICC5P78iC+3Hl7qNy+WPwkuO4ikH1ygMVv9LSjxB0a
qTcNlb6lG8yv/q6SwLEmhIORNSJg+ldyUNBbyjMoQPqlKn8xeXfiePLFVJeegxYc
0NVKnKnP/ix/8j91jBDVnP+yTLWSo3i5F3LsZ80HjSaY8veVaF1tbZ6jTya4lOKQ
a0X6yms5a7HHF5r8nQLiWFtcMroH3NJ1gotIukneEpHBph6hAElRTa7gIDyOxWZ/
Pw1+0FtEvoZSeSQZeBoVmn0Hhzh+38W+NP8dJYi4mtAgXoKAB85o24QWgeBtckAS
3Qgm9jV3i7N04qBv2D/+umScX1Yi4Vn1Roa4+G2nB5wlOSO2ncK1D4prDAyA8dP5
FZpi1duDyn9lwa0f5KV5hHqdwYkKj5elVofN/vuGH5Mk2f2tHw28FiXJ7yVOHKgm
HFZ7QJ8REcQVm8p5G5SyX7y0+8b1JNafsAXH3nq/WyezD9hVMI4Aru7M98AqfrjO
jXPdQfuCXvIINMPdCF7CE7ViXnaFxphluH5Ij7imRSkGFa4oJAJbKr0RRd8Q9qhd
gFSa20LKaqsA41HggER5ExAUFuWleISPNulSEfz2fw8pwihMg9WGMOtfhvnhvyLj
jEclLdVfemeDn9v4tEoI8HsFmhbSH2Jw0v6d+tl1DL8b1opQC5EkhJSRv2cBCpKv
WgoDe2IkhinYpm0vSVK++OT9REHUknaovYKbr7OqDFSHv1jPMpU5T1r9YB6oY3ae
Zf7Mrd4dM8X0aKJHO5pOj2Z9U7ga/qoYc3XkeLasIq6YRnIuhj7DjNr/WXacIJ8/
yhcvNVNHevYOLJL1Bq8oKXBWIX3KH5rjpvEQ4tFFtInix3mVf/HyRVhiji8+5tvt
2orm14Ou6WomXcJX9puARfMSPvTzhSIVWNfDhgwki9EvqI/CrDp8QL+JcjGe109z
IMAp+wa7GbQp3KUymMtUE2h+m1gqzHD4yDUi6S9rBr8MskqP85nnOdpTsumfeoVm
hYbIv8skNQySL1j8g8Uw6HF/foumM/JjXfcQH1bFOOKC+vQnYZszK+BTeunqyTdT
IiZQQoAnAPYV27V7fEQJo+pGQ6liY7PwS1e7Vzb1/fkfGWNdTuH0DfdGoCoDjzpD
gX6G/3JI89RN6U0zcYswleOFgRtqgtDAYvUmCAhGfSO1tSBISRCxz4FmtRLggjB3
rLHGpYoZ7cYD84Rq3MuQSNxoxYcP2H9ekeoouJ/JDxbgLJaOU9+2osjwir3vtxIM
0Y3NbAJ9vFYsHDTHDe27tUH6kWkE9Q2PFjqn7KFL6O3u7Fu1NcD5zggZlByMp7J9
7XODpOSE1D23nO6EH2Y71xRQRy3fc76vU5sn7TIk6Y7w71SZ/o+4AhYcXKZnx7k+
Bzko5eqpJdGZFOREeF0P1CUOLlIFb4E8mMDoyzxyPxQsNJg/qeVsLXWRuUP6TJm4
SYaOvaRosOCbk5v7AQf2aZuz7SB0b0HQrziY3HPXrkZaGtsuyk3/PVbMQY5UOx50
ggvOiQ77c5RcXamvTEojF1gG+6asGsJEGBhTR7W1VmnVfpJRIG4bsMkZqT9MTGbR
ca4thAnOYDP+iCHq4XgZszXbCkeosHYSdP81WmP72hwihsFzvmghbLybV6YsBUoV
/QOGAYGT+vFH9Hvh7Iwbw//mSv4Xr5VicdIkCdzGv1aUUOlzvcOeMHcvUTnm4rtB
NMWZWXqi6ymjWgy554q4ADDHlBBHrbwOxDRSsCEWuMrOfDdjiXZkJGlS6IskQink
RtCptg+zyLO2mwXhKdp/D3UFcTbZ4Ql9OkxAnVxtv+MNgc67Zh3Fkv82sj508Ksv
G58yTMOvPivoArJZKgZ0qmgaPg8rUJf1hbsZuNFjeV5MYdg0/03tc0JDW7CvRIyy
UUR/P7uHLnSPuYAxem5IhuDgGpa4MZogVjdOlwK9L3CXKArelGtUWrzK7Db5U4Mu
zjTesLlpGheexRSDQ6lV+stkK4HQIwmtowfKIIZGhXu3DEsxo5dgsQCGYZQ2RFdI
YVElbz2w1wmJyl4XvI5AHcZlKJRBqtLptzvh9iFPtHH6EERGFoDFx6FR0tEh42xs
AZ7ew09iBOJLYr+y6ulyo/LwBTG35TR75+MOJfk7V5ymWGIqOfOr/EI6a1u7He6v
Il0iNsMCgO0GJ0OnwsFjLVqrtN8BpmDevCt2JUHOhd2zLs2ss9t8JbcN4D/6AZ+N
2woNp1Vr6Qb/PQhS/Gxx9yQj9pxpTopdxgndbpn7zs2RnGVu4FsQ6U/kUfJ3S5nY
cG9re+A1NvHbCGHJjJdjr1vdoJsvNuUJeiwC4Dl+l6StWOR+wDaIr/JaxGF55d4M
+qsGBszKHWml54NjCfMUDPAa1VDmUz0ZSekSHi9XI+lcIgB6f86p3c/qodbg/6ru
mpUbXaHIIi01sHtpRriZobEKqjSL8jnhO3d7rLa0rMYQiQRiEEt+W5FfAp2jyxfQ
aNRDb4A8prpjniYEd1z2QVQWHtPDvXfr0uLBOBUZ6P8R7dplMWLrh8r1b7YXEq8k
5jUrHPQaNquIokFf/TA/1BCvLPj0sVM7dHh8W7y32TWnppHo1ug8K8ephufQXlZ1
/WQql7NW5YCvsbM0T9iWtJcqpdpXTUPCjSSCgdfh5jxErtc5FKWpC/sP6gyl41jT
YPnuHyGIx8YTy3KEyeAfITs27zBwvQhWYIHqqW0059QXUm2UhAabYaICtQwzmCAR
xVzsWpL1gUEMoKhcq+TVgKEHGvwPW4jZOl+XBnkjg+NpYzXmzZ2vLrZq2n2TMXoA
YfFh2zjBnCwi6419T+32AQDPOqcqrMK+EdD7wyU7vh/nkD1Q4PrFmS5wf88APWr5
TgtJ43ccRmhyCG20XVsocmpodjXJi7THII1E1O6YUVwnYA8iFPzwBzfGZaJcIpDi
ULXBRsqFl8xWFZ+p4dtr6Lz0y/84M5QPwh1daYDFz6tk1XGhPOB4FLXxzxnFRPPf
2hNN9p9kcURM91NahN758AwWmO3R4k8Phwgogw2kvSykvrWOWUeTf/L993Ebp7K0
3QDjAdBIUlAJI7GgaPg8MHdYFUkB9FN+8d+l3QoGeaN27ADsinvNbDW5TAN18bLa
g3TcdPxeb3H7EmynFQCzrwzhuWNsA7/9dLeK228ymZDj7zLdNJyTl/dY4wo+7SOo
/4pqmXa4O8OuzvRGhAmxKfWzxEqQnSvqbKpm/yC4zo+rsO/Tk/+Lm6OTAKjbNfqM
xjIboaDLXo5dtwbNIwXOGC7mQAHRGXqfLpcl/q00cEoTx2DL+QH7ybz47BkJ8njn
Y/RBV/aNJk6z6MghDt+BUGUUYUlF9RhyIvfxn1CGVRlyRtSnRbgn/7xgx0eaGBL9
uqUhq+tuCdDrdX0RCOHGHpfrOv+5x3J9/d11oNjBWcK+z1U1/e/p6sstIzeK7Loo
zMuW0U1AkUoD9clzb11tz0gxtTte1x067KYoLMvtfHvPxJ8ji9QD273EA8KUQfM8
tHetXSjhyMMFiJ349dRg45BbXAxp1Vt0cZbJGHGYesacHtk4pq7SeJnJXbh44jqx
7FMf0NXk2sGYjEM39XfI/KkqX3KOzw32NS7EGtNYa89VBLTL16q9xAL6/LW07f6f
LgEx3M5mMWJqiqH14bzHvl4ol8iBWP5kduwSLhCEZgLPBYiXxtwabrl3hxnzmiVq
67RrElqxtVtkXY7qkkCBBoieLHJSIQDAXPjfmWhKmHz6cN/GikKV6pTSvdbf9bXv
dGdfHjit0mPqytxEWmgxU6Dj3kZiGVP2Atlb96up9GTFcu47RKwbFGF3I4s+cPBy
YK64SR1qqX3Lwq/8sMGruITdG9uQRNUASMm4fF/ASa9blAc6ZeudFKoNyRazhrza
6A7U7uWM7iY/bLJBpzxKxBF5EiFhIHLT0SbZzPqvE+XlhLAVBCNy3nKB1QOQ20sW
lpwg3T1KfB+dsZSAWMkCLgERAoRde1hVgRDnWNTiqgFevOl31867MxawhcnCqEkI
ShbjAyfX/tFp5iQIyjFLM9K76Sn37GNKuCU72D8B4gieJZIL73W5ip1HhmCMoTrQ
69/+IpuHbALCQBSGNuJjciVZ50TJdPLTvGk14SxI+iGnfPc4kheQw1TA1SqYxzgx
ZAozvxwWT+j5yuWNb/7ApCxbYFNLj3Hzd328TTUMW/UNapoTymfpHs/KD1YoCGJ+
ITEVLHKYgjG8LCBmGKbnlxSUAzKf8zse6vSZa1K8WZmaY31OmE6Tfs1nxMQBhHon
I29MBmrnf21MygTmrRQ74as/EfB/ApCx/6knDcZcOeyyoRd15N2MDewzwP47lhot
MSHZW3BedtPhNpTHM3LHWGyxbCiLaRbdrQpdXwoDByHSJ4aUUQnGikw9a/Ka9QJh
o+W5HiLcEetj6TrKUh6B38H7wadyEOK+ix+OIFK/2DlDjxKZCqcLYwEsKqFI0HrJ
ohb/42BAETUX5yIZTabf5GQ/yyq/9Hdt1M1hEmQb4PjU02XTi0YW0gWuAvd2VFS9
/OBHWFlJMUlebTaGOvaCJKJ/IieyIMhShY8itQQ07t20e9u2398w+JG78LrjALhl
oPzBmpPR+rXWDqkkD4uWSkuOzVmyNGcEuvlcHE5gmRePQWNfj19bJd+Am7HiOFvC
0P6PDGRklO7OTU0lFTc+O4SL/y7kn7Av0+5o6YKtvXKRksMUyoWc5sn8ml2H6/Lj
QzzmcJ9bMjLhwCNFavsRStm5HoN+d1UxwjR7RTQBQvEwPqo047MGCBFcOIWZr21L
tnNfITKRnftLrp/vAnMyxlJYEUVCnSdW1pZq6EJ/HaPQZPsHi8M7t8GxpYeeWGje
tAezy7phuc5mYOh8riQcMIRQsGaRnPRJQLBI5PBHJghtJKJvH2yUHMI1Kp+V99A8
f8zx7DZR5SkVRDEyyOzPK6tv4cposSGH88zKZoZm+aL9GCojr28MZpY6jCYRPRNB
V4HNnZw5zHtcU0ozt5xRkCdF3I0tDjQoxwz2Gj0z55WDTgizunjGSI2lXVZ3KhRU
dX1sYPcIx9rBG0Oc26q2l+wQuezpjpR6RVnXFKcY9Cx7t7/Ic4wD2Rdhf2EO12jx
HB7AmePk6Jt6n+ybTOqA2ub6BgWPw+5IdBcP6IA6gchUm81IMOZTC09LCv2nXqHE
N3Qpzk6JwbwG7TNuGPs7JhUT+oXES8m+kh2JvUU4BcGwIV8QwCdf/7vDnq1tXvJQ
ORV/cFMspFnXptZChOOgF8Ri6YAqAj+z1vaBBNcJUdTWQDTDKN/oIpVguL7Y3CPP
1aHYRAyqjlKeTHTxG+lj/rCqiDZ2Hrn5gk1FD1wP6NGTffC6FzHUJGr8TsBXqNyp
A1fxGj2yN1QfDFadBXVzXaJ96eo634MtjSzYgvnO0Q9FvtjWg9zDxsExb/+DyQsD
Onnle70nJGqqbcOWEtqwsrcJPDRNpwi0odizQBTJ5/Y2qbBhLYa9RtGNcJ+T2G1K
hFx0jyM1tTTMWDZRD3sApNEJg0w4/HXNteQFiODU2vKwb91bpeeLSjSS4b3kokc+
q8VKAH9TGXVrU1IIjD5wPVBUEW1kKo9vWLcS5W4IMPziasvGmFow6KF5MLya/rz7
Y8C6S+Hky6Ws4aGeQp3EXpaMQcui4Kpm42ecy+K+LYaqsJQ4XDgoC90zOE2p1JjH
9vnrJjRC/73dvuxwmGMVc4xRw6Y3EyZbk0FcWfOcdyh7uUxbR+snMXAWx7k3l1H9
0+KuYEBuGrKRKCGj6+GFzsKMgR1GrZDNu4fhG0zOU7zF1YKMlcE/0HIBhAXX1eSK
7GGxkOdsipMJpQxM1ZaUpO9ScXGTJBHBjQOj76alFpdwB1pXWdgd1z12eL8JcSw3
40p3oNOcHXfqN5zQDWFATEYf3Frp96OearWqb+ckkEkYircJdWwZvE3PEmFlba+U
AQeLIGOS0IICA+F2Mg6iok0mTovEvouxf7dgVcCALLJYrEcLzUh1fu4P6TJQH8eT
KTKIRO/51OCJvks6inXY9JTOfZvNkhXd/ZUVhY7U6O6ETk8cqpNXIVRa0TJP5Z1R
T7hX3bRgCAycl+6et1RQq4NdgKkv9T+qvkJylc1YwzaB4BUwjDgHOc3WOMOqqM6Y
Da8GgyYEDjHnGE1smcSjDgMUQlf8xhWqqBE7N7vdh8fRQd+K5hA61Yh4Vek00Yge
pcdIFxmQkp/oSFB4rGsykfSb/vcBSXdvsHju0iaBlxPy9fupiCubMQy4xiL3YFnP
BRT9hf0UYiCDIqnLLzzfEJih1SxWADobelJiXPt6LDRwg7y8Ey0vTLG1gXK9drkX
kKDvGQCAYJ0zej3DoLq5FHUjX7eCVpJXUBZPVFuj5x1gE8k7wvHiK9RZlB4OO5ok
8rpieUuOm01UHS68I2Me9DwCkVtXAbNWiULTdCpji9A9VtAXT8aMIh1d+VL36b7R
+UZwpm3nuwkIxe334H6XKSyDG3fGbUWdn15qhkmw1GocviK65xC2aFwiaYDlKWJ3
NbsE7e/fYOygMD58aPC/blwW+ZVkBhqiYvCB9Ix0rSpeADwxK1aAqoJ0OnE6LrY8
vYfoTu2IeMEjR0kZb2DETcrDHsOxEs5L3rKLz5a4skkxxwZ6CVVCtGFOPAUaBV9O
g4lppSWBXrSktE+B0oOM2wR4XCmP+9SJaWyxvSHq6yvaTsVCPBTGuv0s7NGGRo9M
E+PYxFP0+wse5VCzrnURwnEriMo65Njx4F9o0SS56JofWWxGk5OYSQTo0fE+w2iX
9f7nEbW0rq1zolDejn/+T7YoRj0vibha/8yvJV9ytYcyzbEwvX/MA9bL3xcYOql/
qlvv/+i52Zcdr5p3g06GTV9Nh/EDFFZaDXbGFPVgZk3xdVFdDJbzagoO1UB6ePMQ
p3Ovg8SxDGQcR4HRQdqDywhAxJ0gUJBPLpXy1bzuKMmLj2a4hxiIlA5WNgF4ksr5
QxM0zGIR2N9aTJrzi5D7YjNNhul4QqwN33Ns1l37rMxBc+9AUdXSfHZBIf71RSxH
lxmHu7VFbX7ztQhFRhkrRAymS0B7nt8i0PB9vdaAu5P7oA3uzn5QK1Fq8MVX5LgE
l3qY1RtWxLLPdAGytK/q7spi3WccKNnWecOzFnk0ewo1gVIBIHFVrGv7iXeH7/YD
f0vCZqXUscXUrn45eddFJGuIKmW8AVeF2NzU6CemSFX9Oxmm9DilDyxh8B+VkK8m
IbV0kKajtGSmHoH1qiEj9IlMqv8+m5YKgC5v3PA5N6lXKLWEA13Gl84yCq/0sVfu
B6GIwXEVzKzxePoYD7JYdujObFQFBo8OQX4Daf4KADtU8/udwW10YYxMTGb2cvop
UQm3edWDZhwIqbgj96kAmFj/WCQrY4Tnfd++mrUk4/NJ8WS3/j7lMGwIQ8FLiSzg
4vKAKly50hbQb3QOo3m72W4PWyuT3fEss+E2zbYCwgTrEPeaTjmsKrrILPD5Iz7B
Lto9BgvLe9TKxfLmF1RJXfQztsFJogFxwDr1L7GsbbCfgFVSAqhKlC9MOJY424uc
eUH7oqACQ48cxb31ugKNKnNLy6iVH15sQK4KywurPIxaoFpI74DgMswUelKoU+2b
7UCAXVOFkqH9nVT6rTwssTbA257WdwZOdS9umPvmqJWH9hXOqMxkz5dXVKvWRJ3s
YazXEAoxvp548bu1h1KPxvO8lxI0vMUccWtkf+wiLZv7b2pPoDki6b04xT71mJub
s38KJ6MezNQ1LvXJJ06BJKCPv+v34o0OPb+MIV5QeCOcpUiVdv+IBdPv3KGB8d6a
L2h3n0X9HRP2lxjvU4YVPQtP5lLrbGdzmKwairqXFQ7/0H9/16d0LADTIq70k8mX
6E8IFcZipe/IVk7tSXlj/oI5eF6OHw1+Ye78SLbV0VjqUj5mwHGoU4SI5rtVc4Zh
EpoqxZgUVRK93DPleH0EVWYvAq3UugjfYH+lu1lCt+1OfHDTh5LxnCSiYsD6Dfem
Za6KdPNZbb7h6sC2B2H/0rwUydeuLDrZNetEz+DLLrE8z4iGSB4uUogW8c80gcXY
KI68ui3iT+sIh8Q/WCiEKE5uciFfXxieQIhPT1ouYuKApru8f2QmjDWbxOFNjFfV
Z0HO++rDqB5mXercMacxziD83mUjjns7NZGh2NmTQ+IehRobAkAOFZtnb4+3zFeJ
Kik3Kq50P/RDlo+4QezKG5fE5d6BE9MwewavkK0GufIIe7+lmEc2qaMykKzkbWM5
SKQONVgD0+VvHKT8/WbhxmGfBqvnP6aVk69Nm+uHEUpZaLPMMTlvmx4eYr2mXlBo
utYtrBxEi2nWugcv3l71MzXqeDEn11hKR80I46QvIBfCXL5QBfJcIDlNSDjbqdLZ
j4KmA1Ij9bxtP5CuoLzmdD7ptjDgG/cocMbsa4irQkgsB9oTvKWr0v5lEfsAWiBt
h2oMQpD5xnsPx41KJmdEHMzNA5O0VImm5rUrb5y3QVv5lRzGsTWoBqFzd/9FpVXR
2owexwVrIXpJhGGhaAhwVVgV8pWBXZpEiulAPdjBftxe2AKqNoaqeTsF/LIikzBv
MtQ2EDSP23McsUDI7jBLJ8dQiX60SpvjRHy3aS2uUEW4OiJMgyo8/K2BYZxlW9C9
uCaeOdV10grNmI0I7gs/TuJ1Uz7mpFCYN648NMjL2yQdyFdySmfp5m4+DH8U8uEC
J3RjDTY1XkY7WLUpqa+uesxzrM/A6rfexjD5G3ampASctRGuTrZ+n9zZV+6M6m1h
FmkkR5pbYBlIfvaugooYkwXaAkw3snoWI1HKKgd94JAAocC6CIqXejsRC/zxDnfO
3dPLmr2UOAjAFLoy+bz8kbur+CxYg++7nOktM6JgQv0QDoeWEBNmU+r6JUHbndA8
PvCiCv1h1Mlm+/ackc2tFeOheiQJPlg3jQrLnI3mu2OtoCBruURBCjbfhlla6J69
eqRE3ULZqKYvooe9RVbMP/zp967xU3wdgiL35Maf66Y9zxqqsFtYNYRtBR/iyKQ+
UjtAba1aPpCfSn1NJB8yeXxvhJp4xY1qgEYOxUUlw7ApkJdzvSEETNBaxL2SzbOf
eN2BqJvAtkVcCbKs955NqnjRACoG+usmSXJuzvmeKiQ9Vl1xhzIxb94qduD9cGeP
6rgHG9NXmRQCaKYyKlT0w3uSPME1Mf2JduqiMiXAUzfqwoqmd/GHnMRUCa93fYiD
m2YYglslpEmHtUEdnIgA92/nn5ssIRVeGh5LKcNdTO0FgcK2aiDYVJQKxQQHpBtN
fqLnymtu/xC+mx6vG7cdrXOP+Um1Y1umqo7TiNCA3QmAsPjpNMhHJ85CG54wO4QK
yfnTsPiRymIPJOWeSioOvdDYL+7/pgDpR2HOG+34pzsH+XQZ4TPraLkb2A9lu/sR
HMDWcqj8HestHemrgvTjJ44FY4+G4+lyIjFbAONBh3NX22t3qq2WM685j0b+SmL2
lBhm2qZN0vl7BszyuB1DQsDUWcFuAaUOQpBZQGHHs4/A8MCyjiY0+p6PUAloMum7
AbugkfQkK/2pN9fqlW2fEkdmiWlmF1yJtIL8YWxF+f0A1lalHZuEudBeFGCMWbvq
XkCZh3rrkwFMcjJ2NhMfy0V+QGzc/bNe7O+rs0c/BCXQZGbYgnbka7HWgGht3ZEp
LAjkC0WNcWq1IJUebQ3eiIE92/rauKA5vRYjhoiTHedxZ0OVkgJIN22tUk+k0Dj2
ZVVYrNmgFk7hn2gglGSBrL3dkLphcLButQc2S4B6/Byww1GeWQkXYrvhcc/gt4A7
SgZyit1KXjsYT2FRi0BbYkEStmEXPggLyYwUXtPameqMGOejkePhv2Rp6lXwPc1O
TD4eZILM5S7BZE/vYbynwf0n0wzo87/hvzzeE1dwLVTCbkrqAnqAclUO59ZO786h
U1go5jb8f+N4f1rBRBvNsUfpUaDvtuQ+0sw2oJ3qa7vjknkrn2ce+pR69Uvi/ybw
Mmg2BF7BzH06orD9kRdGg+SUmJryGezN0yKEKbgCMXPqEz7Df2rmH/f2nF3+bwG8
+MPZetfaZeY8pitV7azcnlVa5Dqs4PH6xrB1b68wlSGwQSsj2+dA2h/WTKNfsVTC
sJd4uy9SDgsyxo579VoTIcwmHaBSgJqmilIuTMboGldylIj7KPayFuJrW0g+DO+i
Qk0dtWvCEf119sfppLHLIDVsk0xLVrE+8jCNaBFG6afYHKstuhV+rYS/hEz1JR+K
jFN9Ava/3tDJ4fiFsklH6gXCEXjeZ2mNmepIG7t7mlr+SfTSyDaWK9VQU/VAVvCH
eE2m//JGKgUKgFP0ncKW5epgJswyF2RUJXajBp4U03W5bkPlp8hk4r4RnP1grVJD
6ZVbumAUiNRW3NHnlb/90AqVI5/L0kRr5oCiDQ8giTuE7uN3KByNRkw6kb8u2LJx
WApybRo783cAHCcbcqjAe4Ou7XT2eqrjCIbYjAkUk9GtID9egF3iWCXJ+ljXs9DS
DYrwhC7jj+IcIfBsMCzbpEWl1mCL05yh36RXoiU2eyq6wPyHVrqZaDU6L7QW8CuU
z2Pq4Ok3s/sXAhke+hciNNYWjA6kHjPqXpaqkGdVNU9p9b3t9qLY5nlqTtpggbf2
VGwB45VJtIx2iiQgT/tvuTbj/dm+7SqAsp52XpjbjR1+nueeW3HEYbeQIGR2fH1u
aPw1OVkBULkpnm2uVWaGiUWe+ykMWUSCwrQI8kG7cg3IUXDRkDM6PKI7iC5e6Lsw
Lcjyf1gYXi6Hv64xl0sW9S5ZTlrKX54nRcwti57ZTs1iELsnA2d48aum6iGZlOH0
VXW3jucqK2c0NWt6/KRBPp/wxPTsz2H997Ajj4WpXCeU6vEzTqHrpHR6Gg7UmbxC
ksYpg2WbiM/yoXr6Bixdgph2KdV6hjSexO0i+e3yvv6kaa7sy3Eift4b7jhTEGgD
SeLJtGEyPUBQAQ02c9Fvi5IVryi9tvx/4+iCf3n5NGATmn27qRD+aIpirraTjYrN
inNFx9bAb8YGxmD+Vh0mJpyPW/HBWmQ6NYEUoCnrykJolHTJ42/xyov54yY5eET4
yPRMICftLy9LPkfvkTRSo1GfmAJCrIvC1Ebx3T7Vh09NCTMoS5DHRyk+a2Omdstl
iD4h3Q2o+fWc6cSe/8jHaC7d/Q2RN7PFcgmG5u0A5UyLKJPFqEUHVBqoNTqlePxz
pHpVYQZHMQW7b8h7/oyxeRaWJKcOiClJ/GaA/3mBX5CSbacT0jvD31tkPkkYiWzd
vw4YnbJ6oP0h2MgTQnxGkbA8wz8ykBXJkYHhoZFcGDw7YXK0oTolZiuEDUFveM6e
f1CJMJf8D00CkIu1wJpbctuMtq/X+jHeUis0xtA5YrmV/cbmwXNtpIDkBXyVyAcQ
ibMpvpdeexflPb5UJO7ipEeYDCsRJpwCwjpUpLFKGPbbamtu6gTKD+r+nXZz42ET
X8P+z9qNgcMiBWxJvGIcTqipr0Ru/tvCCF//JlHz4HUGOWTS+qrQ2oF0RImKG/KY
sWoqKn+UMl7YOT68hiDOxdiQzJ71vxQs9d7mpZomjsCM8RFlb0Wo65vS4cZrld1l
e1S5JVU7hO1DS8HxetSsqZStNKfv05kRb4kIpygm0Uz1itZ2FUTqsflrbVaVpffd
/fR6uoQ3DmCn7HzgXi32gfS3rv6tjwCuP0qiYgWGtMjt1sCmFy6jSoypJU7ygN85
Vyc3POnuEcMloFm56IMdIxr/sY8HbhS2340OVC6F8BqX1pnJwDSYyB2SYlT4b3f2
HwyUcNaS7aN99zKF0hEZnBbfd/9QAfNG/1cqHXEqfO2Q6C0nNofSl9w+t3kabJV3
NSdKlIL3JZmVGQ19V/wYctJsAnKbOk8OqMbiMLUxtmpFQ6msSUny9YlAf8MW3f7u
sRWsXrCOTvcFfjG8o0WTYT0jHmez7JiMmqnfbPzHggASdeenfdb4wh9NdTdrxH/m
AlDj3P+rnyKQftAzar/kIx4Oen+N2LnJRUYydfwXgenIKUvHtovnCovhpt/10u7C
TWjuLUUpR0wtYroyYTRJ3QQGzFG86yJeMUJ+LLlpxMF5vwJStJ7XAoJ/5Y5qYixK
daBSYNsFaAaOrf2nbx8kOap0WICNu1ZulvSC7psHoGsb/WUsbT+X3yYooCbDCxas
o+EinLoxpHf4LGmlA9fzRglbOLmuRi+T7uvlTGNoUobxO29KwYotsBjQMT2WbFxF
+YEspys6PhmA+PVYhRvZoENAJwZnigiZep0x6QdkhqqkcfDliPN02kz4jUZI+WSC
IHMi+aqHwB18eRwImjdItvQdMJ4sqO1K166esp1XuvD9R5atum1INskbGRrGKuzU
ReESDidSwJbGf+qNfONLNawlnMzF3zjjVmLREpvUvxp5NkhWYiKLbop5TgIbewGM
LcT2fBVx9NbPyBcqDkQG/B4Q7d/9/pLSZYjgzAH5Vjibl3fB/J31s0cm1cAftIzn
0InhQjXdZVQD+DEAR+BkSiF5L2vEOpxjObO+nXuWreBD2D6/VOzECpWo5NTzsF3C
IqN/qLqcCk2wteBfQxIqtGEON+gK6XnLyAi0fyoxDqVtX1XxUBYt2FG3lf/33FOK
QDsNlccm5mVzUygp89AT/MH1TdCX0Mq8TIO3U0AszRCGREOSsUTiiajKaz14KSgr
uBkGwNj3iwj2JvEBWFNkWZ+5WjTVfJDxkRl6PlD7SHkk95CJxH9mmp7lRqve/LBs
0tM3lQP7EPcGM3ITUphhw5iPbmg98RnfYVlXW9uum3LwVeesQLA6uThBxSH9VwWT
nTPYYlPYz0c6ApONr/m0ls7J4eGZGb9//ZEYmC2NGtn5iIpeKaND/uuUOAcp5X2P
t7eN0qFNDtqaY/GX6sQdLiI4NdyRy4/f11WiSxRXr+HaKp4rE82guuBEF3XlSJ2j
JKYC4FE1o4vl8MiYh2kAUVeQy4UG1G/F6Ggqm5DlBkwYv8vTFd+e4qrNM78aOuf/
CDeaNxfQVwXG8z60og3v9WG83/6xYG2YKQ18+/auJpDoF6MjEhoQmpGslMomreGv
05CdrYEqvdiIhN1IsHubU6+GJHIskahxwtqb/Nl+R8EY1YVnTwIlOUwU4UZDczTp
gt1difD0kyTVRRJWqa1FevBDUECj1Mq/H1xfKoAb0qD2kK05f+j+Pn+yTksiqgOO
oHet/z9ZvyWm/TvRuELCBgC7szk37rqEJAsCkFK3ZWtWFk77kDoEcZ8rbLnZZjlh
c+fOCfwI/UfdYMrnx582UkSdGhBguxSP8EwZwQcE8C9YUw81r0t0j3gpyUSvl6sn
WWlCSjzS4iWSeJy247CZkCfVWxOgrGFoVlNrFyLxhz1H6LJ+TPPwsac4QPlnzrqB
+MylINBFTfhPvms/3RWf66m/BBu8joKpH1ZUHQnGiSWFWkaWUxevyFZsbU9jP8qp
+hJoaqrLvXsB2QvAKt0gRWvfdIY5AcKK+mnuqvSAk04PoDXi28EfT5h3VvyshTkx
TPSdx+o+RvsqzCqRkGAY++zBUhV8DoX1BJ8E29jB9ZfESv+KA7TetwErNcksY7hf
Odi3draKXoRsWhmroPy+drf8SOANG2jsh2tuWBJmWAKJ4yivbMbKqYok7kdXhCpM
TrYpwB6tqaaTuapKFwpkD1zviAiaC7vPocNoXvdQgZkajLwYDGsH94O//yLd/1ai
GgJmfKO9H6/MPmSd4zze8QqDU0/rnGLCiefk2DZvq2S23E/FkcXrW5HCmt9uw6+x
wJZZxemsfK9hgdonmzV3TRzHqmeB6DMI/gV+g3uNdFeAllzhVihVmMeBQ6NQi1lv
YXudNKnMrHHoGM+3a2LOxSSQb1AJOe6MVRHJwCjBKibBcT8KOHorqxpW12ut/5WZ
N4tAxCU32fNePZvW5Q5V45KHYfx+G3deRO0VUl46uy33aRneU8+nGcHgSJtKGRJ1
wocixgL+ZKlFb4p4tMcxdkutsBH6yRi3QvXLp+LhnjIdJSNdQvh731gBj+X3tW7S
E1XNkzz7bjH5T2J4TQ437N2KMV/LNYTiUX1MqpUSjAuianfSvQ8Jb75poU7/iCrX
6+BNl3msqTU3NK5L34PBfQrV6gqqUsto+lUILFIYZGLTLI0/2WVbzWGWCzKGztJF
0zkDdl5BQRS475cpWkkEgENMwjWH78S5xBIFrxJEIbG3pjJ7/QbG2E+wnzHOciSe
LP4vO7Zaj8b3ioQUR3RYFZa6esPZq1E1CwmOXOnJ/T3JYsE48+fSJnoBwjJe99d3
jR2PNr3O4tU50LbMV/VfNIMI29G5/qo/5/Cw6rjY3Gb6n3jKsUhPuTE404R6Mn0Q
xTCn/tqEgK4nNMME1091nl61MuVjWfMgWpdF/GROMVBltLby8xJM0OXqoaFHGZhS
sllJ2EWdMp54+j5nL0qi9jDCsZx2ti5BbWPw5rC/mzz1FSOvZlXjne8EcBi2ZIpb
I3QmD9yrqR8ENVqkjnJoAl/7LhaOQnYGnwo1WizqAQ91p44oYrT5XseWzjWyv6YI
NYWkSMHqrMudGB5ioAjK5SZB5yP0cDd0MwwHIGyip+7c6vzlUj84+6a6Vck3qtIG
1uoOulyBbw5VuYi8kb/RZh31wH15jilYDR66ufRvM9rQ6+C4c3Dq3brwjASSPKxE
4739f7VYmzoDPvACVYRnAe9Mxa8tRboldprnT9DSARq6etP8k/1XuDdYoVfcX0Jt
HXNhEjcpVo45cYB16mNJpzNyhOXNj0THpihxvPsDnzEi2SMi8rrC4Om9fx6ioi/r
6bt29j1m5nR6AEwuBykNsCP0REN4oUWKkg8pXAnljftc7le2pyi/CycXPuex39wb
sEWAisRKN2x2Ywhqj1PjG7IPNFgFv+VhwvduRZAMiweq5cea48Ja/UvHMg2fc9aj
//XvVmSQKqWAwduQliAIqTO2cWhu30AWIxwtcEHiwkcYRmOWib380U3q47KXANto
7kDBTegtL12n1EJt/5JTY4uEqQ4RVoUlTP7VnD+x16G5w5KHZ6yW7sxR7WjuIzja
7pRkyMXNDkO3O8AcbmO9X20c9MYJg3wnmeJLADZv4t0QKfbaHYGxuYxtasZemern
VrQ+6Q/2yqHpF3p1Z9+voNL4PXkBzpw5J+yfK8azqJKRyMytb9BoS3+vSWUTgSIn
N1iUWJBz+/pBWGzUe+9ZhiHxnx1Ed2/6mh15FE8SzwYzLUD0/P7UJ0gyMDTC9Y+8
rpsXtEJW3KdNSjW3ZlUYwUiLMnMOZ0gj+blr8C0BNNPNH/CRD0iIibvr/Jfgm8Af
JLx25oJkiRQJerJDGRfBQXNQ9z586PO8rlvtstgK8drPdIohgr4tkes/32TkZxhZ
RxxWB4YuJm32kTizYjRgoG3d5VWIOoSHLyDnsO+9mgzHQW2FPECQYYle7G3wmSST
b/KI47voSujjQ81f9JqJLhQGkrLP8mUs3PnjGyn/ATB2XNn9tCWOjKz9Hjh8J97T
fxigzu76M4yz3MAWIlUI+fsrS1avr3dLlVn1BHKCixyj3fAow6DFG7EGkqc51+Bk
zyevW2yuSm8abqgBKm+UGKJKtCqCzdiOG8TRDwiPkRWeiD7m++V2eHWfg+iSV9/m
ImOI+M/mLR4FVMAE2Hnbkz/ZGLiNrF1/vQyskYpEspyQ6/bkJhge6fKjoOKpoMFF
cDnRwTnZ+twVgeUxXaBvhY4jOYkFWKyd6cgnmaz0P4YV0bd4cDGcltYQ3p2KhIGa
JJxgSs/UDmMpRUcxhK6jvsBXMupurvFK2+DJG4jrIjXfwaxnM1zqMd2NAnRudlWi
E/LxL94PGlwRH1drTJQRyb+nTonapnR9wP2XjK9w2WzNqsPia93VT5T5ytjpXX0I
6fIzjIZYh3stR9tOikFW5LNzW3H5wzqB93XJwYERNXIBemvXRWiBeMomM5xDmYjq
x6+3m6VQ1OiMkXH0yMRuUO26jxyjRL+AkPyFTV5T8ldUqxQXUReIQ2/AyKTnU0Ac
hAW0yxbGuSsmaeURKG0Y/Bz2Agyk6BC6nElAyupQEYb8qj4Jvhr2L8Q4UMEEwpwv
vfjnNlw7PQfiggON3q/D/9U0wqrYpH/IdLy2xEoB75Y35FTD+p1FL5nF9DTIlsE1
U+xcvXywz8dMOQvD3axczERdzhEMZZX+vnQvKNa0+XG+RnERMx2NgEEPWz3US95j
LRtDLjQkHJkOa/+DJmgpvgRK5kOnhmj4vvH7Q7wu52CPmhLjjm1NATbuU5v+lx6o
tqLhZgKNE3r4FGHtLCw9gpQSPAebhgwRttslPzBvskVnuqpBblLH+wVMGl0p3I5d
+J/ar63WgqqQN4WPlHNUyQKPo2EBXqFpfcbR8iu4gW+HlXKmx71VMaa7F6X3czw7
6+4sxQs6rL4KDSTCgTpciAHAxRAeZFn2S1CzbLWcJLT92z0AU+s9vZCrF+tQe6Ko
5UAjnPdc4ErqXQo4fVOXekz2kBEwUti7ZmKX24UevVYB69seb9V/dOTmQcK57dAs
61YSNX4paRQmYXfH+vdsKVCo/OmrnLMX7CHtTC3Dn5e/Z8O42qPaMdEg95/NQ8DS
SKPqq9K4pqA0ysoNE62BlRhtOL4+UaaOyvjbK1LFz6QahMY7usN7jhx8gFqhmlqN
ecBOVPUMGMsQkub7/MA5fro/zg9khuOHkumXCW6mGCeyOyOoo9aB5m5l/qYVNP45
F5K5j/RnOFT6ACIa5bLgyxqUhmDzFYmfweIUuP+L+fUG+Zfa2Bsf6FMTniOTOhwp
fPjjB4VqCwIOviRDi0UxWAwyJQsN2i2oZRQG5PBzrcHfAeyqdCctIXLSLxco0J8E
jefzvF4j/dnD6Occ1jVh6WrGWsvPqlDMjIbXrgAfAYPDShHVwOamRknGNSOXMHz4
xtABoa7Xf4CwtGYSi4TZeic6SCzggLL0FOCnaazwmXrqvP2NwZ0bvr/ruHedPFld
muzQvGTEcqmv2boJKNmMGG1PQfY/L7hg/ZlXEg/DQ2IsgkQbl+/WV5o3WEvuqkNu
PLcME0wSR+Lsc3rPGiv7Q9OWl6eWrwtD55MDdWeyFLAQWQynE/v6L48rQDmnnMTb
mEGTq7Sq+FE4h3q4PRnQXbSa4l0bZOaan780a7Iq2ZA8Otde0Txx2FxrAywTgq/c
3dGgINPOt9MzDMv1uqaAht2KT9I0L6NPIrcxgwR/bDMOIcr2Xv/hHCo297/PtIRO
vsJkmNj6F3sS/5zVtAvdzCFPZObdf907O2sCjWNN6LtozK/dRNs5BRR+617AkTBM
qKqTWIRnR7kSZG/F2++hVi2011JuW+bbntNfvM3EATAEV9h4CyWDVCeBN7NBRAjL
IDjh9G99/SUCVuGQcCN3uWm+/6AobBFZ8bYPdN5YP8r6U1I0RCtGZPzL+j2YqKD7
tuWrS1m2gvApBS6jwtNcEoiEAI5rJlW0tQfly/qjOebQEZOVW8qq3o5KHDYXvnHS
GRGC42VcmVeZ4QlwEg0dtSwKwyF/WAYuH1uGUGRWXtSrHYPpCMjmCIgxnoNMAXnq
v0OGJchHDzOndZks6546zwZ0Hqvz4H4uTjMo1mrFWAbm4C6mP9Q13dWerE3ZJGBX
p8ydl+cIhHFvw7fV40vHl0AtE8s4DR7DX51n7A0zV55QKfrapdeeJW7TUfV/TSc3
PHeZzGvS7zUmDr4Xp9p3khRNYmZi7U+ZGPlu/rBTX2IIu3SZTq3wsBviRrySxo7I
ItfKFmnaUbjeLEN9xXTvB4kAPBlhOs+GrB5/7KPjSeQjikr0BkBdj9hNqavp9xwK
48TcaRZ1InRG7ZXwvNmoOtocHZpvxM5qjSTCNxZDwMmExf3rYPsFMWxYtOeReMjK
KFCOtVUEcDKhN37kFbRghWGz26eSH+4KNNY0BN5wb/Q0/6Wbf9V7K5F6a7MFOknw
bZ6gc05D6gsHQvw+47cEwwIcfp8RgBPyM8dF0Rp/LO7i2/qlY4ExX8UWVy86enpl
wWcnLBAXg5KzBwAt0Sx4r2NBHAfWXHt3D3G8gDQkc57QWt8eHR1nHcZjhZl7WIks
7Q3/ES6RLet8NArFeCfqgI2eL/DbH0ekXruF+uHqQfaZikLq6jqdtXSkIfxy9Uj7
5XxhPNdeLHCmSH6Hat6Ao0vUOCHEMton4ja+53SlHY2FBRoFcWm/bE5QH1MbtHgZ
5+w5x/O9MTqCa4ngjAT7zLiSQ3JiD14bLj1nwgZqSnaoEeqBPcZMnFLIZaRO8uep
C3bmG6P43vvv/AwmeN3inh9OC5H2JAj6TvRrnYGG1oA98d4y7iJ5UZX4X5sQf3fP
aH0VtDlpypoFtvWZd9ONkhYbJcc8v83EvC2H7Wzc+XhLfL70hQYwM4Gcju6i+y1v
HiWrDv7IeEcbzJpmlQCJA6SnWz9he8oFs0VsIx9ln+TkG4Yvn2PPXlQ5y9/BNVeZ
Or46m5mgXvRkoOfJqm27CXPNFxdsyn/7gNcQTZ3WPsqUVDe+la2NrRHlvu8C4B7T
jw3IMv9xYkO5GP3EPg1eJb0wVJ1TPOcuqtdQizLnSzTNY3L2Ua9v3fWARlrcu/qQ
hwDKKMqG4q6sGrk5qljnXsdaLJTxG7C9vZL1WzBZ/x9nOz8Djv/gi9bqLFzZtZiB
tj5nildZ8J3EkUcjXYcjKwwRwklOcbRPHYNiRaKzwhBYeTtijWJPJPzxBgOEoJ/G
ecegkprqLGsdeAqHn18n3Kc3tT07EzY1ojo4fQTN9SAg5xCAgwMY8qZYtYP2vIok
OJJLDkCDUzEpIAVg3bwI2Hafp3J7SJIMYBdM4khbg0mwVbTSmdGW1RlzbZmxS6vP
V2gFxYQY9F1Nh5yBnoDea1TziVNNEA5RkuRN05oWeqye4jMpf8Q43trHoyIT7JTi
GkUirOZD9lFewgbrMyUtSkIXzm9sZlit6nz4/g091NQgCH2slnxbla/nDdLVnBvF
Flv/tAW6T2NjRL8OzleKMtboEQReR87clM/zp2pbVcxq6sCf3y9bTeb7E6zLIukX
cI7U/kKuWjuWwU8uI8mykkitVTHgSKUqIPTqqllJllMbdtchalXgQ0np7y6ekjAu
vZ/u2wg4oKTlc33tpKuwGjQ3aUbDOD7BuUxVCkbS1nrEnzhesefsKLO6QP7019TT
9nyuSRD2FVcxaLQOeU9Yw2DhUWfSnnhHwUPt3zcAbCGVZpTTAvPkkqEF3WahCQ4W
cQTBwmeByzeRAzsLZ+FgJJ7aHkhQRzhp+c42f5o3qeA3Iw8hQM5aBbebrxkJf5Nn
GCfKnYsolpkPLUUdY2L2nG/YwW/ODxKrgX/+5277DP9IKT/0EK8yzSubd/r2zJWy
5iiuWpkPT1JtKmgaKzgdjDof1hgT1cXA+Hxrr6BQBAm0xq/FrJ7FLQflBKbWtZxm
gAogxczvPCra2iVOOtfFV/aX9+5TRZ26edaKJn1PdsRlk5CIiuq0PTenmfWKhXgw
rpAi3eGo9L3/wiysgjjCpwzTj3VO8V1mvKYiiIQdbSqvn07xDxU90/oaPVVngmeG
AuEs4r0SvJxwtaE001KtuOreRn53dYEGwIvAp1hbKIFz4PklUeUdPwU97gvd+3h9
10MeCZ3U5bIXv0Z5Z3Qf2xeBsKPSAV8J1oPafPGjNLNkL09rb5rlK2AcNwKJto86
sEsmrqspBBoIOip8JKe/OakEDKICZEfJGvf2clnhW0DVGoOaVLGqGlEAnGdF7fXB
5RwLNhqkFzBRqeU7BTKkcPmSDOsoARw/vi8WP4PmDjKbKrkkQPgvLlmsaEniM5NN
6IofYcWC7D/8duszXxU3UksGh1MAmo0pjoL58vIYvWeozwdZg/aBK7QUoVZn2MKz
qQDkQHT3iEN2k3iVqZayFe7jAn0RPyDI/vk6bTWvSPWRwk042hP5SmpaiMFTMJyF
CGUgj+B78llMyNBLjIfhboslV9+Mgf9sy84godT2IVgiewMN8avy4SpfwPKXtX6U
pIMCkQzZvp+NKlNOhrjcVtCUWA5wszRKuaz0Jo3rzgkKLfoQt4ppGBmQ5m5EjKbq
yDn5UXbeRrWhzA0FkmEWsMIngZkB7J2ssY1eaJ66+ECkbHUNj/3OHEJ6GPP36m+/
4rzEY08U30lzygdtYi61qhCpGuIEdcFDggyk3BGLyTi27eZIYaMyWPWyFYNadZt+
9F+sZSNQcVPHzvln6VoVcalD3clQqhl9MqhX0vOvt18qOhRbEEuJGTnEQfF6UVlZ
ZuO3IoYBMD6tZ65CDLey2Qs5sgYHW4/4ITxPRHOJfU+uHZrInLxxI2bjjEebh5VW
dmSlw7Er5SYJOxVVNrj8iGLZWib8wR7fgKy5mM8brCpW+YICWlOoVQgFYlvvhRdL
3SptN2mOrt12t1jz67KYn6yHG3hNpqkEprnCvXPiiL1s+LzcGk95iCLgCVWFIKin
MbWU/OujCpzaF0lh8lhCPlblVaP55k0oU7WCtD5Jd89Eu8TUU7dHGwjlVbQmu6DM
M8QgkvT0w7JA0qtQKMnnJypHj4Q2+hOq99J3vCNPqBd9VxIkqpWf2bBfYqOMMe3B
BmhIW7DnHt5nsxOWyVggJQqANzHbNXTTD/889n6g3r6cXIqKLpIip2aFsaSu2Bb8
IKWBKrC/To0WErUsrM+nGIt0qjFVd5VkOVShDaf9dSzK2pO2VzWRQGu2AwMMpbEn
fH1U4LaYZu/5Ynz+3W48cJ6arCqAiSd89ntIIrT3PH3Qgr04m+LLpyODPZurZ5yI
bKCD5CmMGD+Vhk3ORSrB3TjcT2573hJ0UTa89DWmGPrLhuCJrTLTBMDfIFlzQJUd
s//NYaIFXTz/GlKYHGeZNxyacYL5/cs2aufzGvcFPJCCwM42gFdE9M/o1lAksvm4
GjRV4/fDpZpN42G7YDpdl3nAQ+YWTWs3JduC9PjDveqz6bpEzJuJ4dpmVk/N3MM3
nxdxWnWpP86dmH2affBnzYcpW9cRNPVJGyctF4g9lS3G6T1phkAWVFvDJgTMQrWP
oWhycYgZOBGj5v/yJhDGvSyojvOsDeFBnECfMC6vZah5265DbnvVF5uWgiuYt/ZB
v8c/+3M4mD7mxJLIHXNztuAnDowBMOUf9ZOiSL+gWFVwHaPk5sRvKbQgSCbI7RZS
DCqhC/AhsoC6m9sPHoDxJyB7S9EBL7JcY1l9OCoSs+wv+rbnm/kYN4ythgNVd2sP
E1Siue4nqKkxxtM5/uVKZLztkWMDD8/PHpQcMY52y+/k9Q1CWz+YNhJNiXm+vyj9
rWAPbMeRVFr7lwit2VY6YLOgJ61EJGebsm5Vyh0PWSIMq+BPse2eQmELXv3A4j40
pHzMZfiMHhg989PxiOdmkW2wHodn0ou64MdnD393NW0vNz2bmYCdDxxbDPhsG7sv
XX6cwV+eUU+mNKNu+0TI1CbTOB8r9ClWDCIKnnu1Amy/50Prybx5M3dEg3dpOBbU
XN8NThs0x0wBDiJ4X21bOSpuyHijzevAa2ZR9L3U4a8FgJB5h7ByGUGvtqq8u0T0
Gi6K5eKzY/Lxx9xmV/q7PANvrTsvgGsy7A2Bdr2XbZAtJX/g/wiqj2DYnw/xHoH3
98AQxSXh4KCPFPtkewouHZXAF93NTGU+VNFdWcqWgmybTB2i8UJ9ifoVBdh1UVYa
rbqJsBFyVE7sQnr3l1vFvP3W2r7YqRY+MS8zzTVFrgNF82REZFH0vejjOW2+dgIH
yFU5YwL9v2WuasTcJkeLYLAnVGsGzv5/N5dPDSR+/ZhYxjHblCVLkE7vLJnzy6pF
3kYrlhgwnrhUg3ysNtuKkF70Hl2AGG4Its2JCczAuL83dU7jpm+phm5cRlHDulzD
BDgeLUcffMgv9jVHSqXcVH6ev74WJoZ46zlS1UyJ0tYNPuS+oY6ZiaFB7AvkY0k8
ETQFloib90ih7o9lZx5yFdDx6YoAt7WbQ2TSuQWz4F3H2ca5R0QK2ZT+ReiY/aph
D6h8zl9QEGGwNp9YmJHaiuzJqk9cNa9lhpf+OXP7FahZeNsmrxTd65BlcJyk0lSR
rvwUgaM/HnYmbwLyLNNMe1Clr1nw5Xmcgq0z+iZdG6PT6LKYbnWmwxB5tu+1kMJi
Oi7ZOIU6aUHqI/5DHLXt5wDi+g2J17nIXiHNkKxA2YbJB5LAl+HiEEdvXLTNbHAA
QE5yYIab+xhj7VBmvfg8njmoJk/2f7MvWwP17tgC8wmktYPzEOlvbGk5/PoLPAsZ
9/KxQ3tT3kZ4+W+3ONV4Xv2pyKIIDcu5RH2I5c+uJhSWa2uQ/XZEJapmViUisKks
bqpb0DVJ+6GYljxWlctCbG0bQCf4/DjuULxvNQ/yYTX7J9u5RBx60yav2ore0WXR
TZGAojTRmeNsqdeDFwoyBdZY0rd1to6QIUWx276TRQa4He+bPoTXLkM54dzrAA3u
faWlsTf8OQKESX8iikYeP0hp1eFSZovIA7yxhrvCeY1b6f1wTacLc6yx19REudpM
luw5UvJAALHgntndFedXqg4z7/iXXxZZSphh168AaeBz61ckG8YU/nqi/OWTwSTA
IJFhjoR9OgstGtgkDpgQyxt5GhNFvXOi/WaJcRwIAk6cppsUFZCS5nY9ulPPlyWF
7mmrYUZdFu0YUZ644Srwww9fq4lj8lQYHGIczvVLSvaEelo3vDSoPkwdoz9UtmTy
4ccHv9Xd6qc551mdQk4LKiwlfbjrdQCXNBo2igEfhubiCxJBDDBhhY4EkelWuNN9
x+E+mg8BEVswpI4VfKBesq6YGSc3StPza9ENWXr9iDLnYWTl4WUDfgeJY0CazYhM
C7Iz9kiM99TisYGhQOQ8SKlFRzZ/RW3dc3WohnwfUkOhOqAiwHlEqeM63fvt3YVJ
bu4R70HvnlT8D9CpGsdlut5bDFLvNWlghkfpBTHdoLUagv4qgkicrDMRuT7KVKwB
o8VNlZ9A654ZsmBDJflkrOMNvkFJPEdq23/NOMZ3J1ZnZ39JUyGDm2VJzkYOo/kW
KO3hLQ/8EXpzHeyESxGV/Fu0R3LUkNc0grd7OdKXMKLEzIZOOaIZsJbTHo+RRCOO
VCvoBP7fA60EahssA2AHweo+JWhZcj6GY98npoDPDygZ56KdSEElawC+0xhCImkO
/XEQT5uuqSLjcd0nK9cdnyyTvDZxqc/FoqKy3uucq8KN667JDtdqXEHCuWgSlR33
kkjDQecdQ4YYNoA3vYJfyzz/y8zoh9O7eVhNOV1OCUdG8UPBb/MoA9mhN3Likiou
bdiVWBH0fowJmKxhGxQopa0ZkYRXsw6Ti9/EOYtsMBSxW7wS5OUbgBw0koytW/Ld
PhZPtHyi+9ZK7UN1a3xX8rYGB5N5Fhz2cd1xW7Sz13gC9nSQ86Ki+3ChPZor2bUt
pAbdYck+rFf2A9QdgsyYZiYcVibIBndT1PTTZsQ2g3603Ir/LUByLJz4LWFea1TW
UFssnRraqn3JSOaoK3v+jqdLrmhDM0VJGe+sZZOpAEBGea9XSf94YPyeP96k0zbH
fRs1MzqfUB/HgVyZB5mmkp5SqHuooG5YnJnlFXQO2Nooj/lhMF85GWO5AxGAdCuE
xE11wx5xsltqwWXOlxU/4h+FQeASBazGQv6dCN8y1oQuBKR0mt6QlkKkpDmKw25F
8L6aHJbRimUCJBqduDLkBwC/qzsr/afFVkYAGKxHemEoR6VyqChe9KoOSiRBbmZB
PiumUGhCpwcJFi3tPnuriVmtDnHzoa4GpfOALRmjBnuDCp/qtdhfvGIcia/S2f9m
2AR6quqo6ht75TiV/fdt1FlBorl39s73BK+lDswzIt0HEaD5WJZKqAMMRku51B03
QrZij/AF1opLWYti2BSlywAL3qsSsS4RvKvwIpayX8UFhIe4z4fxCboyfeeshUTn
svwms4rl2wwFIPngrC/yvmrd8hM+oxLLkI4lgGhCVSSXNVGxFFwiaC/wGYVqZ+2u
4emdDD533T7YfC3Enj5IwiMXziVX0mRcdFMTHOB7tAaOYSk1nFtr+ZIrflZmZPvJ
PTvd+1QNNQOxzbgpSIMhcjIqv9Id8UeleQ2shqrLm5PfJ/Lp0QUyMrJUv4E9blQ/
iVlw8qvuCFJmrAee8+hnUHNJi7oHO0rnsowwyH+mgmqnK2pUQzZG3e+62fPYo3nr
zKyY9Nz8lnCuqzcRi223HUWjxW9IEWpEGbT3f7E690Wl5DFNnmguzfEKBNCHkvJ9
5KdZEyq1CafgjhVmUAyIIFiPpzzMdiX+CZAgE9OOd5bN2HnhpYmb7Tc/ioFsrFhi
ivI+8wgSl8Ci3i3S87BCDZ81D8GL1fJDRpe53S/9iZ1EG/fF+2cMzRoAWY4HimFv
SlHj6/ZNHf3PjK2Sr3c/Zocg7MpF2LoZegAtT2X5NO71WLJQJl1pPhzHapQ6nGvF
n9s3W6GwMR7H6e6J/5CAyKAnDOOsVAnSrAzpLmuWbc4IHg6Xjncg5CcEQkT06GUS
jLnCZp+slE5VjhVNWth2yY5i1dTrIkHoubHhQw8uoRBRIF+rKJMyd9wt0/1SbMgR
UNInTa95vsB4Pc6gZ8XzCCUfBzZh6eiiYK27gg99iknrwcCURJCHn8JVJ8vM9oIJ
7/Ka0jww/K1o0Xr4df/WL7DjOazVmPC0OBE2lmZoAqkGveAf+GF3RxfzPTZM7eQ8
ZXmpV/HKPdTP3p4LTasgmBlFQHZlA0MOgIIvsGM6cwZrLIkSWAWD6yaDRUcoylnO
MMziHc+LGQcPfVcxbQcyxmZ3qAF+A7fAPvg4qePY1nti/sWuPNzINTwV3v7a3meB
VDw0C7vRYg2fXlgxYV2iyoWihu3pGpk5UkKu4zpk6fv5ein0fsEgrnav3DBLkDf4
ypH6KB2VDLF2MWlmnxLx5y2nZSraMV/PXzASkproYUER0awAVRDvTvWgtsqsx9XT
dMPoZI31MgGhSVH8ZKIlJ4ZAA7T/LLkfx7qhcI/q4A4TUtYvJzoEFYX8RnZ/Af8Q
ijiyWShcLj+dfBrkItKtXN5RYwMRsCgGZ0dgFtIfJIiFgQBc4sE9WZnKOppV0COX
MQbTs4xV1Q09+bpPgD/lslDyw85cHmDDi6nhegKo5ceTAE6cD/2L4DRybZH3LAdo
UqMqhKKInqSfhYBrkcAE1hpnliRXalx8opCuntt8vRHVCOKERKvKcIG788ieor4B
y2zQlOIvRTUFPDhPuIPSygmSUJ9bogDzrmzFVhKD7VZHWGFqPeh7vpZk08NA+AtX
eNfXR/QApMBVjzW7fHpbuSvnv4awbRZdNhERhBYIScvuE/0VFsq5Zxrvb5UpGHIL
RE5NngbROCPL2+2hPW58zB7y4KDCxQXyQU+O6Y+Lt+jS9tQIJSFjJeNZuWodYr5P
ljXhTxiLzzxIiS9PnZLFFo7FdAIyZWGaE7uXyM7XMwS8/TiIKbb9YHpndYVVKdp0
dywufvmxVPPmtEZW+fVqs0yy6ImhJm8jMZpq8x19OmHs5kb5uUbdi4Sihwio3bE/
1E4HzQxTOwe/+xOz7zfNFggoS9bRjuLxo7/uzLNG1q029XpYQvAk4ndRIyAWEv6Z
YlVNIOPrbfddMlKd2+ZDxchNukOVjQHwmtFB6fbdzppzqCwq4xGuRDntHw6nzSnM
97tD57xbjE72abM3giv2ilIQWPTk65tmll2/YPw0VpCTL8uKG2SsQDqYRJOncvgG
SA8o9crr6+n2ZBARZAi7K7UFISBgOIQQzKaCRTAAmkbAmk8uaDestR+4kl8O9NYq
dvqy3eg7Nja6oZxsK7VMXGq91XRWc2o0UQ8njtggO49Tt8196wBLvap+8GWgfOZP
UY4o3rdIwig8O4iZjAhd0LYcBZPBNnfxcQ/3DQev8qQzEXGuGNHpnH5Nb2YTNyYG
iTVel7x0PFxfIYMYODaZIUu6DxQms0vu+ek9kO1B21QQ7CNRN9XsYjhDoZljmrzb
h8j2o1aKSKOV4spYB8mc0euTvlVdWQldMUkj6R+rIJTtAZJyh9fIReFlLl7fphnZ
pshKFX4jNtOd4BOQvllMLy1kVS5GkhFt1IMwzbfwRlAER1p2wZLWH3Ixx5MoJGwt
jdZtKcJAF9FR/o+BM8e49CFL9jMyCSJTQr9NHs5/ubzhRjMCbdGFp3j+iW2Ky+Qb
dehOgXZjQl8cF2n6HPVqbMJDPjinTgIarsiXytt3joT1UBsPTHbsJCkxkjUbDng5
JKAOAYs/KkVCe9Kvvt3PAei6d6WZU+2TaO+mV+dBYxBWMKOVQUYPN6zoVHW3E471
4E9wY1LIOQGDWlNul6E6uxLAecXwue8whVwa5jTOQfB85dUGvqEzl0sHj8UkHexu
TQwugIVx7QO09jvYR1YMOPVnNMUhgleIdQAh+i0pn47gWInr9K1+V5M8B6+M3FJj
x/k3RUzog193gt++kqA4b18IMhgiJMEhTtLXcRHWF6EuhRdqnKpzaeaM1i0aFhPY
lb3it1AAKeFS3iakcRwpvECPXezndSulm5/EqW/pBp72LKw1h6TIsFAaXmdGehqV
8JJFMKK9XYHiyOjylTjvUELepKByF8Ha/QLjhpSWc81qJ/eUT9wJZO5CNJKXaEsA
dWEkfDCd9mQ/DuOp9SFavPQ6s99dfn+JIyeJC0Is918SRk1pIVdRtWjVfWZis9EI
np2Levq1zs/GkweGQc547Wr1oiOnv/5U+8Qc5oKaRfEHwh+d9659zCk4tZNO0iXd
1uNR+Rbt7cIhcwE78egIiL3iI6n0epq9pPGC5MwjSmef4HFJVyaz+vP5VDQfvgsh
ZOVfc+fR98tz6OmYpNmib+EV6bwczJ3hwGNPSxSZu63Ro9Ql64y2ccQCziiYxKib
8Q8yU0/I0AdkvaaXDmlFpeIIeqSGYCwnRtMnnjidu2JiOiovb9xrQ4iknql6ZI+P
QRDrngf1JSPfkkehgsb9CLiMmbbSTbQEM7T3tkuGj3ydnW0AgNuIarRwRs6udZRg
GhLrceXgc3MhO/8CLFArne0BjHt7wTAxL5dn+dZk1NJOeUFOm00hNN3TiY5ti/jv
WemzQ9fs6Q4Q5lHTL0blPTvzwR5ihYdmz/3SXMt8OhBr139BeKe7IyFyv6mCUOmM
NY5kRzr3Hjr6V+CVV0a8RwDULyM+xeATnfIEZCR+EKNi9+GKvQOWSI0xbfiak9c/
OLk3TDieM4KjaPnBSIcGK2xyZmMB04eyr0swzEVYPuUguDntljEhcmhKUg4wzhlh
y6B+fBeG1Hhyu7yZXkbRvtCMqL4QXjUITiuiwJwP8aaBMNh+6EdQITXAFipzeEi/
/kVIni3PifMMlziL/XJhTzxYl8ywovTQZElJnoqNIvtHhsrLKJtW7JlhSXo+NYAX
DchFYSKFf3kDtv/T3IXO/3GXzrsmTpFC5vOnFZSvsbYZOk66g6rngDH+Hmgyc/Ep
XBGMeh24P2TIrRhh2A+pm1EJmyzhIQXVCSTrOkQa77YYws2wXvogJyjNohKjEvFp
OYezQUOtrS1YA0BcgBpf32dt/evlMle0R846h4+5qHP2ClpviW8sg6z6VsZDBRxl
HQHJAcZYDX6WSXc4se770/Nc/FdthKDG/fhm4CJzh/QrO1H4sLa5RSJ+uMdQQusy
SmyBc/324mjrgiBjzlG7cbgRmKhmMTxytt+JizgXAqYrG16rNwqGs5Ow3xliS7m7
WFCMKYRHUrtB9RfXFpYtgoYorkzuu5dlFGAuqae9zwKFssbBFCu/8BI+iuoCJnwc
iT/CqKC6Q1ixapbCNzxGD9BE81Jb+mhw24hEyTrWIyPdL2+pE/mmIMZ3ucx7dabf
Hl9Wwcn8X0uQHCNvD0BDUZ6FBiFYsqiKAjle87utm1XQ3MYauaPaB5zNDraHqtqa
mS3cVwnP9JgAgn6z6NQ5vqc9Jf6RjqIxrCMumsMxuPdzoOGy8vGOSK4YcKP1i49i
fuF1jDt3S3qJgGpQam+Sjb029mblc4v8/6D+3TxZqLfaAyK4r2Gwt/EOxopryV7r
YygxbaTR1R14Lor8m8Qg+O8sxa6CUQh184hZBnEVaxk6WC3fSa7Dq7ZP825swJhP
q+Y38J/rdGTdZ701JJ6vkWlWKxPOJZmRKpIiwwgaimMDfw6GgVELSLn2k2vNgTgm
kD6OGvLBDMXunnSh97ZXrAt5zuH8RVZaIuUXwdvhdUHBh3dT38GeTGXAQKcegjg3
uyQubDf0O4GuqY+3autFr3H3Hgh5cuf+yMi57X1przt3m5VstM3h8T1Ea79f/8J/
LKNmL+Y+gF9CG2nxq1wdKfSAH4EnKRQSAWTzk958LCFSQonfyocczVcyRyUaKP8S
0kbybj0OtAPv71juT6DMQgnLMpea8xKk+164NfGFWNRsLhHPh4i77PrEGp6qMJTv
uf5J1/stT1n1Uznksjkj4cEFk72aJRGlHu/EzqM0JinymoZbUY6W+REM57B2tt8Q
2bT6A4EkuUuO+uUchHrVMf/zeEL5az4XjyF38YbIIWyg+ad4w5B6eg5ueILGpRmY
KpEc66FvNvtOTnJT8xW+iNW1jtzuq+YRQ2oJrWVQ3TiFtwZhSFXSNewk6u6d34Yt
3Qjt9LFKvVs9HwSlXzsxWNKxytzEIjYdcz8RhQZB5wDJR4O3+4Dufiz9hY98Q8+S
SOMhBxZgMhj0CWVQeo/BhIwhXL121Z12vDeCO/FCEjT9z5/b+iuE9aysAJ+QTFfz
E1Nyhl2suJQ/JPgFoz9uOeZMAMoMDTGs+N3Y5w4E6AU75FOYUttIaTRzQ0JeHIe7
dp4oLFITRpsFauaOIA4APkFIJU7jGBcZ9ZG9e+oi43zCW1RKw0HZR/AExWB1dwBd
X2Jvz99SGUCCuVowNxoNsdNqBQ6Ebnzrmc7F+DqdxzWuRRDFY0FGadgsnGXo0a2f
SBoxQorDt85agaMO/MPNY6AJnGH197B1XpWYJaChoIe7g96u6PWw4QAuVh6WfIbY
f82lQ419ZhLwSft5/LeeXxX0/iLl96+A3IZxCc5eVLs+5Q1iBALuPbIZcbaSTcCt
lPy+gDOhaDRedmuAwz5hQC1IMgjifZkNXmfRSwmXOhYnk63cgX7cqR7dlseGBEaC
Q0DkYvmE2dlc8Bvd6LElMW0EiktYCc9RCrQGAeQHmijm3jzqhRA/W88hcEjdcDak
hVpC9IPe/k137bGSvHY3PtcnI3gF/eaMT7R8x10Y3MU314e67OYZvSYtcq83AxmX
s2i3YJkwml6icJNpsRxf/OIUzKupuX5fhdnrOOYOQpbHBeM6BL04ge5OOTvDDEDl
plAkWnrvgKSzwXJmVrJg20ULqZLD8c7dUBeVjdpINBQdagRL7ryjbfKc5sD9J9Fn
mXaHOThN7Jkypp4FMvNsom8mmPCmAaxrW35w2Z0i1OwTvCzgBPml2C3cPJoLDTuA
ds/3iQaeeQ2Jf0Bpzxp1hcRdqUoUaQPQNZAnAkCKp4xCA37KfjWH225pxHmPifBf
I4OLBhRlegg/LZY9SP+qx0t5AHfobYctaNo9kQfbamgxCmWydt7uZ1gvMEJZGltc
l4el3ODKWBe0nozs8cPfHaGBXC0nCFV5Z2/jCSd4RTcYzgICAB8PUQQDtjV1RF7x
RIZ/06lLtVuHhgUny0FQKnd1QHZDTQfRscCrbJ2CYq56TGC5w3Xoye7JaF/ayDjH
z300igRbgEpuhziV+3qxDAOlp/VYbCI6DR1OgKhpFkbv1k2YXohbBf/Cuy52j3PM
rv/4Dspk3EnVa8DK0JerhkrgYRtIM/1fBpTbgvn9S4vA+1bdiQ2FThWqjUeoNxf0
VGka1SE0/lxNB46NuWb5hPF8CqtkOmKheCne+D6inB/EYw4CdvI2EoWEHiG9D3dF
4ItheoHCrfFUtBnnEyesmEmD4dLJ/nsZ60yyvc6llrp/0FvsJeJrHB5EYGR4d2Sd
wAzdv8FeeemmNL4Q8PqLiW2QRtQxXEfGgYXdvNc0xtPjPegkHIzb3r++uZ3Y0Prt
xEqagIMy3GkQV8n7zw3udWBZMylS+aoXD8Ne74QnO4ULsc+pjZjkpYUcAEY/kwDI
MdMVJYFdPRCGCivbhl57hqF+lSnSoq8Ub7yPGO30XM78uTGz2ckpoHItgYm2g45A
W+WGd4I3f+4oC/8ilhlFH0wNtKloTpP8COKNfCLCFRiAYCvUJS5sKWWDwh1/8xbu
RsOALIJ+E19rhzT2nYACcRUMtlDr9aJjqbzpig/h1VaxIuwmyRz0keLJ6YURoRrW
/6cgc/h5lXH1QMBf5o6U5yvEVqq8R3JPrXaQXqIv96bRhzi2v02dAPHbes/HrvYs
mSYeRDZ8P2ZZYuR/UPJ2bBX96XTRcRr3YjcQL0/mkUGfAm2NLmdwGyzAfOEEjOSG
9T9AO/mGRD74mAuHEtg1N06LUUsaKMBSwk9LXLtUL1uicagGeq/9kBP9kNSyvBkG
VbYFlJqUvofhdqwfbzRR3UahXchMPZhk463s2ZgCOK+/ZE4z3TyAldR0LqW2Nre4
wkYrYCg+EM2+PdUdDwGyBWaxzaxmsx7/OqHfepqP17myi/pngsFfhMl2OXSoXD7S
vBfQXbrvR3pgIJmsbfvNcaHMJqnKsWKUdZf1mQPuZJE16KrXMQLtBgleBCJaCk5n
WBSoemy2+CW/PTNn98JniCzl4FEzu/D+wIJbjJpGuxqeO+1bMVEZqzpVOyuAtCGb
QyzLEbVEKOiSNzZVszZxLvCcGQbq2oO/G2DpnRFv+uPDCiuI6sZZ4FSnccknI5Xk
M7cj4577+Fd1F8uKBHiG/BU3rSONU6hfUzlRYUR+V83hOcDYN7I2ziCNX+dYlR5J
CFRujVY8U61e6Z81Zb01cyHDvK2GmnF8+ARNzte1LL+Y+fLyUGDJTEi2Dbq0qnrZ
h16Emst+T5IAAK7jc5syd6OAhTp5RNrIC71BgMLOV7TNebXHgt4fEaAfjmv5j7i6
ZRkSMhFKWpBAO/70P9pB2XwzoXD2koGqcFdAHj6gcmtH6s3Q0yp40qusW4DDtIuX
BYJMtj2ZF0Ckk6SlTBuUMSVDCRCv6y35v3PkEw2mBjiIVLW64gKoKOcDE0KGZET0
VbuvnNWbA1/J0WGYiPUFk3x0VPM3BlW7yWMdMkn3HuDxwymxu6cUQ2bthQz5t00b
b9n3h5m0uMSk8/gtpsF0gvSbd+T2qS4DJ1d5fY4I/WseAqM0LBbo5h0Q+pjyJ6HX
s4ubYnJtd6POi0XipPrw90PqugM9apN69T6TPkuxkFTzER8lYae81D//46HD52t2
jdopd7OuUe8lzK0ATYfdfvJrOuncxCuM8Cm1Y3fPPj4GmT6bXa+6RISItmkSroln
rp3Jmb3nPZvkDek4z1AvGsdNW3oo6086sn2sf6xUBNhII2O/20NrWJTGaLUCStek
uA5zix55p8b1m+qRZUnfo6IOkMx2wRMmZ3vhfIoSoAO0kAvWK3CFdPF30rfteZlw
bSzVlt6Is4I+7byRtf5cdtZZJC7BgVD9sTaQk/dDewT6uvlLe+/bFjjNjjOvhQ53
6HmNOl/smHAHf5BTaDxD8gFipCcF9cvxXdYw/eAtVzIn+bJWSs2bjdyhLreINDLV
oiRC3wIHty439X2fhk7IfV1X85E9O2xD4ARyr8any6mZTMEGDpXgLMCDNbApsNlG
FumHnk7YirFcEfgAJHkWdvzbJ882KaTHbn7KHoS5zZawpcCsfe3KwY+Y1A9vILp/
54D/KtlbLTdbiP9GUlBz19rXZXZkmOHxwjN+eaXguyAt0+0di2Sbg2p+e//yvme5
l+ywGa5qHTNa+k2MAMtI/4a6leEPcG1CDhptuZeXhQ6CRsJ9wmD71TDYIWdbRA4w
3pG8HExKoe8IdphEu8H/EpBiYPt5ObaxBqNve+CTJjkuLlAEdtWKjXjBZTHU+GUY
ju/N2ur/5qIcElVI26lMMDeEHH720L/X6wtZWw4m04qL2m3xrFNyFjWq4uHG2BrM
nSPJ1RTbaXm2LrY6/q+UPiSg7DN1dL4gF4mX3NBXdsCU3lRk9O1iVFxx7OYPlzYL
2xGTPeTJa7kSHhRI2ZK0kAeJtp0ws3lw2fQk72H3+Pz+B1qGj6CrCJqUvmONqUZr
7tYjacPQUWahDWxoGA0p2jAD447JP/i73UkI1Xbl9vmJ0A6jez6QK7zWjPBVFoCg
UehMQHDiFVrs2N0Pcl969h4OyyaMK3VvTvD3lLPaPLMtXl9zCiIdM0x15TvfRray
YEIoYylt7WhhCL6JQ+7JYQap7ZDYvXdqzSWoou8f1O5L4PItnomcWHl82TYjf+cG
3d3tO4vVROc/lQta8JShsrkBLPmkFy7rtuwkrc5sHyX5FCC2HpgPFaQFd8UQcT5u
ubSoPQewLQvkLMZh6oT4VbH0u8/s1F8jB5BLm0rSbXBGFOfAG1XdY5FMVmoDbKf5
GmBNzlW1N7hJeACXB341nW4C7mFZNvpd0SiiMwTCNxAqBajaF847ZFfQeDJ1yOB7
xzqmvmAbOuZLYa5OnKMdersLTbhu5Sr6nkkjxjco5wxAEZcmMlNpzsFI2cF6WJh0
4HZdu6cg52Jm4peq9V98UWWo/4w3fBPJjAbq/HgpufFdxtTA1HBu26sJjJgxefUE
Gf8uZSVcsE6CERbpJMJt241AeeK/QJ5ZXsGu/BxA3MOl7kxdGz6RBeiALxwwqsUi
FgE2SgYRHVBjYr00z2XWN+t6Wm6lIeuN7uDhMhOaZidmbaux145a42HkSZSneDVD
cTnCXbKITUZXWSOikBRpxD3x2lxuWARoiHQFIuITakvRun0Glj2Jgjk1M08jtJVZ
wVRPJaMGinmOOYvGp2MbTkzTsknDKzE/NIQLEoK7pNf/9mpwOgsamH8duDfymlBd
e9M68TTTBgXlKzF/IKelmBKnmBV8zrdnNU6xc9VOp7oy65iVfJsJ/Wh5gJ5mscOL
SpdkXT2r5YWmUX7xHRbRU+ROg9mtVH21voSgIi9A8SHDroqThCAe7vYTjG4/VYNY
r4wizOO4BJ9szgdGZfSeKI5oK1yAT2m8SeYAtrXWMAIE1kavFuy6wGf7XQEH58HF
vqy1KDQ0LvYPOYoT517KMU6swzKzeam5f96lsOJqQnDPJNGSMeaSHW1ISRdMaOu4
xjxF6Fm3sNdw2aZmO+3/06guGNaoHR58GSzBC/bAtSjecrxJJknTxgiN1amy9WEs
zKbMUia44shRlWSBPBLofBRyT6nCptlCQaoUYCsA4QVs4dEdiZTocTRyqumy1ihM
pKnKDWwCLV2IUUnhHV9tIdmHclwIgBh9Z+m5onXqhQ4kR7HEvrNbqQQe8Xw0kh11
67jo6/emNBmNAfIUQanOflyYMiRPwuuivaGwnzWmFxQI/t1Ji9PnEi3WvlgtpCFw
QdTqiAeNHxjdp9GN152Ea9a8U34H+0OPBe3hfYJ+Cjz44eADq2+fdJ23CiNHDxGz
7xzuou5gVeGfr9eTlR6CndPy9sdzGmEGiEZrdapSGTLmMtrSMG9qczfQkoeBUSAy
209jexD7QzL0YfD2rJDrKsALxmOOS465sP8jqyXhwFJlAqBE9u2Gu4JPTTlMwTJ5
/DfZaA8aXU67zRC2z9oz9nIsKn8oyvZsSd6DHn3kLLb7mF/KUxwb+oh/EP2GbZrc
jFpqr8pF6Wd5vr7BdkatnoLoFKw8HASmYENzK46MYcFjfL+kGW5znth/myV1Dkw8
fpMrPqSUJqKulwEf7wRHjDCUPiONywwikoNzxOGyrCXZ8qdHgU1/mBnwNjah6nKm
2pPQSRnbIYmTRVpV5KAJ5w89dmaswaB4G2tMxZ+hGtVpTls1Zr0WiQwFopkJjAvP
N++tCab9SIjDMVtiztPIA9vcz4/zpHDWR08bsKjzct4/+jSqCpPzVSQ3sh6Xvr69
U7V2IfmHfCTFAlm8AmJ7BaL+eH9cURgHKznKOJ8svPFLndHgLamSuIOat6WwP3Hh
5NwrJlol6HuGwP4QtSS0y9HjNwg9V3ZarymwxuGFIiQXU2Vb6SzS07PMwsSsdReY
gwe+lMtVFvR/jUevNQuFFpS7CL7Uvj9+3N4CLgUYHfM05RjCRq68NqjUW+jIIyeO
Y5wHgZKA0uqlciEq7dLnfYw4bqtrdSEzh5uoaGcmW970L7cLqiO9FVmru09eH99S
44z8rFyx3P3JXT7vmMckx0afwravcqeqe+XFAJ8oc1Iub8C52tcUtgNQRi/xX2Gb
YYMXxEUrN+Ja+qfIDIhSupeh1CZG/I8RlXIWK7DRE3IvmTArm7DmlwG8/bTGft+j
rq6EkaqYtTF28+HO8+jUUanQXOCT1L6vQBxK/9dVQ6XJnfCVV4BWk35ye74Cmbgd
tgzOBSxTFLXJckdrEoB3i3P0UMcMEb5PLLMNkhQTmNVD+4sbyA2JHGZ+zam4hwN6
lYOy6DrnNk/8Fu8UUhh06bumUbS/EMY8jDG+h7jmqXVcJ4VQLNsgxJk3POxRn3/S
U4Lx3J9jdmBf04QNgGfY2Wm8U9NzfHN1EGX810d7hJUXUUI0Js/y2jVgXh5h6sp2
GibJu5jzNVxhyFEO7jeL2UuZ9KfEBg7ik65QIpjFEtKnSYVagIbrW+9gF/8PTUEs
bGbGI3TGwi34VrPqS5lBIWG/m/3Hv5QrUN3ZzOaUjOFkZTrs5ukAGyjBJTDyfbza
CxTAwM4pKZrkjrqGhASh76ctYz/l4TNqdvb3Rw7UMWDYSJoj1ec4plv9JbBkY2Yr
M34sFUSk3VK9f7aIDvBVZ9vAY7TFa9EnBjrAT5W/yxgGBj0unyU5yjcoRPXvz0bq
p4FkipnS37RbDlrU10baThk+t3CSEoBLu+7p/gFDM/x53asPKPQ4f1s8QKU+Wc+y
tLpnOFrIEIrkKt1XdEVLDSlIot01oojap239+aA/lO9ul3esY/ps2JnlcMP/rwUz
QbD9Zc3lwYldnAo5qg3UjwBvhmWJF1K2jbinyRyRp1ms1TJscrMo9bpVPMJjo2yu
CLmjtdg0A7fapt9bDQ/m1kwuF5Yt+2TvbCPNz3zpAUU3d411Ui428ImBTzbE5O9f
ntzm0yoqoW+iRP/bAoDwumKUYwkPJRnVOmgocFCCZ2i0V/SAHz3GmXKSTM8TmuTg
h0q3CuevL0pOu2QdgDnORGdIcOBySzbDScj1wgR/6qDMX6VdkOj5L3JvhOjF3ONA
xBWUrsXdVxlAW/pCm0oOQzm8zXvPtXGRYs7aw/00neifkkIWDeab2tsrOCNRmImP
b5Iwms1eBM7FDN3WJ/hwMGYwcaY84L5Siy/PYO/l6R7EFiaqfU2UkF5cDcs9QtLP
TPLZJNnmg1sGYs/H6t98ZeIoe27G9reyVNiSlQ0q9na+bO7OflmdKFXTDAHpw67P
D4yotgu/3w02Miug4HMXiT8fmvWWpkhxbklkdkA3q6nVdkVM2zvK1ec44pa51tL6
BWCAogyFutU5O/ubf7XfKPhvytyjrcNs197G8YDqOcgG37dBYam2G5YMwaIut/U7
O4ssuCqcpirt/8f+tyIXJF92M8woSLfZDnUC8LtzsB531gnws58N+EKFOGzDqYPA
37WhXstl7hfNwdHF0zu0QoURDV1EOw+2ccgGnfUr8v7mvbHUZ9plutwyvZYRI0/u
LqJ9H8ylSCL71A73eiAAfq4moLNsZu8fskCnTiE+35ZRMBpgiLmZ5GfNXJ/r9bcY
AIzI3V8//6zWruK9BXMXcGJq/W7wIg93dys4MxIM4FYCsJCjLT23u4VXAzYz48LC
p/m2bEprl/hjGrJJD1tyLZbEPAvuHcRLNGag4uiejWszDElVZZIQvoO8tk1ThEzJ
KHAwyrkmi4bGJ/4Ez18bJ8LlDZ5MkveItiBqkSRHc9tSSI7+Js6c/NYNB21u9GEL
wAyAZ7tPAXBmwXSHbZmF6lRep1g5ZyqWmsDCZdSoqxJh4NZ7M1blVNrRbFRgV6Ij
5DUNxM5Lpk6EE+DEW0e1iZTVuTDH7w3cAnUqpGyhAYY9bN6Nem9RETEJOlECK0Ra
/cCF6RrFjFCbgzzOdxS/DCxFlMZ53W5n6s7QNfdkPhXKOH4A0ZpbOZCp+gd8yUID
4aoqCT4NCzEzoYwIzvTtOrdBJWzH10t2W9szR0gxq2iEszMkhJMqbMjBV7cIZVia
f9pAD4W1NqGPuOogHxA1PAmHVTxfKP7VH0kKR7ilMYo88wNQKD+fjL8e7DdWSxQe
Myf2e5JL7UN4eRAFxbyg/UUaqSMwl/4BwWpI4L95pU+hKXwd/tTr7HOcCbYBUDGO
ED4sWdno1wfAartbfcVgjK36nKLFoIVVEKaGGO7tZpGTMvx/0iArIfaayfK+eq5G
HNC3SqUv9zJN1j5gspr/NrJnZ7OWpSJNBHheLgukvstZmUVj5xzUwTy8g8eDRXaV
UI1vbf1i6H+8OpfUNY9C4UDOorROFj5uU4sBU8+N4ebGOixCOE6rePaao25ZPIkA
F6JhvPY/P1H34oU9DLIsouYRZO7sOOFuWLAGThlPH/4Y41UAJG42OhTZ2/TGMwyQ
HjCc/epWk35aSDZ+Sr/4tAE+Ut9MqjWI1+Pb+fvg6k71DLqseDhf4LqfbRc+1ILC
68yKdFL2K1GNR4hM6cUrflWv2tsF6mQKhZ5629CtNIfUa4lxfGL1V+B4kB0HkEu0
VF98N4XrdP8IKrK//StZMDaXaHX844lkCEYdWaqbJFexYnsgsKnWPS602D+S6NkE
0EwmezlOQ9bt9AgrPNRSuH8DyHPWKlVuXG+PIWEbDYMvRDMSXKZzRPbR6c7ElvUf
Aa2+fTzu8SzoKoB6/MXhXNdeHgNjNyhb2La5EuY0LPvnoyrZrU3Zs+atf7uaZnl7
zfSh+7UZ1R88QFoMrQM3ZvFVz7+HtW8CAa84noG6e7HJdAanQtvRYCfztpHwfXYm
5E1fyStK5kOYhKaAIeCHfKgfeC74yI3iCoEyAc9rS+cjOPXaoyBdOMbvwmvw4YUS
N/oYSV1oibff4Jx2h1id8DPzvYEHWpxEoyt7t4E9Qao6dBBDuxy4jDpAQMqppQzZ
8+j1SEUn+1oA7n4hIIQL8Zn+ru+kuCAAQMDZFejpypIFX6zKTYzwyyO4lx1e3Var
JBKtMYbAXdAnlGTC7AXa6yw4P9CHvu0yYJYIfxDmnlkRWR/jt5yY6//9yBcPgJHE
BikDyCY8an0fgm0xPwF8pD7VlvLLgW/aHQU/RrjeW0FpU2HAVQe5WHFFHE5GLRud
T69Ya8/Rj4VuBrgsxE062lIq/6siqPmEhTnrpazBCpHxsq/Nfo8h+ewRtkqPylOj
Fr8VHy6DoZJVxck/LMGnSM6UX3yfR7kkwt80leMpZTQCgJ5OUsyo89Szk/FoPzet
pW8Ktt76F/3uVujx2wmcaALDrN5KhG6mgvFv6R/Fyo7HAQGjLnnt0gdWn3GGofCU
qvuX2htCialTbw7tJVNYa7T5OsvyXFOwTMhBBOsgS6LTpKBz7zR1Hr4ZrA9nH++T
CRNg7Ly+zivshsCHTH3AAe0nt2WRj0P3qFjXD8vaidBB2xACksrzGt1D+tD5Inw0
2AuIEm0aWFqr9H9gZp/4t1XSRq6+W6jriIrtElJ9PcE4fji0OVZt+zqN6mnJu4Ol
vD/PLDwY9C3XblMZjwiYhg5I1sNmrPM069nIxalTY0wh2epvMT2aBmtWzY6vWPSr
vk1YR/tYIzGtqSX14aqPE8IpvDmIwhQK6clSScbKwWPdaO/IBqXGGJP0EeL1R7Pc
ZwpG9PbDjO0b+j/FB6GUmCULBmp6GjhwG0gXmIfG56Fs9zQE5sGIgB+lMWM4XuVS
SSRaNnbeE4qavRTbKEphd/K7sXRYYceM2X/1khVzv/1bxRNpxy7WWGOfDRTkklIY
zOpLt04qrP6rUh794feLa2k89qBPiVvRm/Rcq5F3lKHh2WLvs8H+RNqttGI4DPl0
OCadL8JyvboA67Lcnol7fWV6WJaHj/9enHb35uk/3znkqkJAViOdC4W5GCKgDwIQ
ojvYeazWfGJ9eYhsz4+5NySngfXhxTBAYds8G9OLBQyPqQODrzkpN4qWWQkNFMPA
DmyjKukWbTFGIR3++MzkHhfXoR7gorC/LfKs/efrBx3nIUYy6G3ULFV8q3nnkOnZ
QLe9+54Gq0a509fXafKk66zB7GHwCJtQzPIAwN/Q+SUv6qprs23qO0TOk+xWzK4z
+4UhMXAm/iR9gyTHO7Q+STvJbzIsgd9KI+7uAheLAoo/bqc660DOIWBvE5RWRonL
a+1Xub4+WFYr4hlGzWNNDdZQQUEoUO1Xz7ZFqM1xsZOB/UlcveckNK3CM2iJY4hY
Qq61INsesDWMw/7Faqd+cw8VREW+boiXlyEWVE2SZ34D9z4WP4ewcPXewlCibj2S
XUiYq3PFs8MgIV8GFmk2vohs8gXhXDZrvH8vYeXUu+BlObnuxgffplIYHDtuDzHd
fJn6mByCEfksHII2qb6NW30t8W6epbYMo/dHFUviDeG73FRizUb48vVeBOtaY7ip
fb7WT20tkuEyp8fvIQG2EG+0FrqxvWz+9y+pA8hPloDuOkhSp60mlpLR6E9LyFnD
c19Z+ZeXCLO3gUYFQ24gPX1Ak5U1Vwn7ioaAyKuoDxuU7Lvg0vmXsZNITvaOeAjo
932wbonEkeNnZ2+lDbVd67uvCTmoObVKPgrfqEucdH7Lw+wqJbkoosIq9fu+D73c
TF5Yn38Gt6qMMKG5zvfMBhBYbiA7MAUzjcRPDPz1HkRiurIf4UQxrfZxtobpbG5/
FiMFKH07lisCz/87zuPS7hSTGSzeSSk5RqiXxRIYk/e57ZsWqTI/4oI00WWdUfQh
+KSeEkwrd8xXsrh/V6yNsmVzTUFB8KAqSUQR9DW1FOm2JeYXXXJijUdNrxFCC8+F
BU5SF5civYUBttBETsLUWu1oTKtNGQ4+dGyC84sj7ljuR0SXcDUM7boWST4kq4Bf
TWRFte0HcwYlTpb8hWg0kviTP+7Yt1Zq++ROo6MY0IbNIPyndlGEFQM409wrqeV+
c24Z4vR/XJBxCjW+abhWNOHouiEa5W2mJVGY6j9Mub6+/kxfIKP1rRbD9UZfeqO3
BK8yblKZA+ckopdpAea1R8G2COXzFya29ncXa8AErCX9Nn21EgCd29q2pNuKilWT
QBoanN1OqqvR7OvrZiSU4tdKieXhEnLgC0AWqtwrfb6w4qvs4YBos8KxtZfKwhLR
RYYnZEoLf1+JD9XE+hkKv1Gfcsw8TAe0+ut/j2xqOZwzCT/t17dKbvpMOq+cNRWJ
EUsXQ6/8LEj4ErMcpfuqOIE1S7ClYz5G7UMnPd3h89P9cXT2Ty4OIN2A9yNaZj5u
NLSE8mWXpg2gZWgyMlCffp8mBv9Kp7dHcNMw4pnSQFes9tL+9iK2Ih6OXPCt4c30
5KxYYFRVGsYBuVe3GKvPJj+ED933J/MkRMfiEGrrMqB0/RhHzzCEugmJ9REO8VCx
WR/Db3/8IEnj9m1qaMKYuyIX9+z268hqYrzHCPtZSAC8Ar8KnTPOcgiAxQihhgt1
KuCjAV5j3bm7zbD92f2/sLnIrBsMaFgrQrq4wDfCNqudwDd5vaLKLH4bLeTZFbiJ
cAO7Qq4RUsW4JDMYA+FeKShnOdTkM12UeBuFNm3t+Wdyyj1uI3LlxKaUFFrB9xwH
GwaQdeRD89FpXRpnMo+6QAeyYei3lKHBoB/PEtKqr8lq4T5Fogl8r5xzGMCpTBTN
5hQTHZDcLr6PIFobrhVIcK+3PS3UvZbKfv/ww7v/R9Yyav0HbJPRLCzuMZGs7LjV
gvpRhLEn1t0c8075uDgOn0Km3ueVA7Gl0eiOGt3Gf4Rmr/VWJ53LSbLxgkk9ypbu
XuPoLfcgsf2AuJaoNgoMnERJCOGSgc0k6VXsRnC4AZtEbxNelRlwvf82zj4jMYTD
6BvxcGgvb+hzD7S3Hc69wb1ELfwIFADo2llC7gNlknPxazptwop+XUEwR2kJ2oIC
x5C1NUrD+WS4bJPjREQw0ygTePrpsA62wQdAczj92KQP0N7lZnZAgJA037zn6DeG
8rJFCu0ObdTWtKLkU4EIrHyZP+2EX+qs4bZnKiOTWCu+x4Cc+MY2Gr4kLCIavLpc
aCu0b2SVCARv7tnqj3YH5v8T8/pdgsJMtBhI1kiYArL55hgKd3pxtTF1XE9KDrNp
psGdnamze2tzidcFRkH9ywI0M4DwjrodZYtUDNg+BfbFwwYmeVX7KOKuFBS3SuWz
CX34h3ifhIqwM0K8Wvwq4qBcKbmyA8MLcu0LfCdPtK89V2dWfET9scCZwq/vcJ/w
0v0C+f/5xW0oxa0U+ay/snB1DDFRjjkS8nUp79+2pecb75YX6QfkRBbuRS1QuVsN
PwFiFVbIiPG6NDqGtIqw7ZOKLtgeqef+n+jD4uhp1f8jkd/ekYoC8Ofe2Dgtua0+
FAesovv74Mpv8x9K1YotKPx8uQw2ERnNuGXxJXv8ex7dtlnwMdBUmYTtqv1GKE66
xw1r9VuYWc9nfml6KuP63HM/PD0eEMHuOUXcTvd584MsDWvlx/YMqW2Dordi16Li
H63Tg7aTcnr7+kaOv8YCigFke5zg9YXyRpLfvoza+CBro9NXE0o8Rvy8EyNNyPa5
3Jhkn3SSaEgH0sinrfc4kxmP6QPdBQVbN00Skyb8BwdDBJI0FVEdsWZfNCmw+pwg
E8p2M1iHk7WxQjYzTqjwBya7C9wAN7wI4SYqXj38fclFmZ32CsF7Vm+48xRbz7Tk
kBxQjRqIyuict+G+lsbU/9hIadeNpBZsT9ItBxkMzrN/K4qvoE2Qf/sQnI5e628v
4ghSNrx3hw0OpDBB+PfXMlkRG9s9213lihV9J11Na89zDmEBnFSN+Omn1zMvAfQz
8eNWlNB7GUq4LQMppO0RTmN/KA32yaEE/2UBQfzDw3VD5Y3I1SPuHkMTiIgDrP+p
JGSWKKmz6KWp5LED4NJgl9Kuex9zPAwql7wQQfnuiVhtU2onhibxi8toYtuJdtnS
/euTPv6Nastf5lNk9BLp7eUV/ZqTbjpkSNyaHosz06xoDGnTz0vShIaHP/HhPUQT
Ya9NkBm4OJlJZUkHdvMeEQ5ij9e0sViRal/LSz4QvKLCWWq3eSlhoog9Wl0eO8Nk
msqc4pdFlP9mG9iDa3fdlOuyW+vZ+b02jN3w80aVrYrwKxkup2EhuKGUDPS0L2o0
jymalwGGng1CC+kNSMD40yBya3iUmGeOBKwrB583pfDGwBttqWf+rP+/2cQ5Hsi3
SUW+em2mclt9kDVZ5fS2T94RZCcjccBdKPvTe0JU7UINZVA1GXyxxf31W4VpP4gL
LrywrqpEIsVKJ2G/63tiwyMD7Pv565AUIMoR/9pd9Wye8e/FmFH9RzhbsPVTdSx6
NmPkwZl7LXlgxwGW5qmegMIy9wQsrNaThMxfen/iWdBqJhd23BR+mPddkkcWphGC
vvfEwqghz5AYYBE3F/YrSRxRyI+U0O1fhIZfQOhtMj6iUoVvjBN/EaEGDtbankmb
wAimTpgsGP7uj3cebStgwb3l2+QzFJRlxhZpjJ98riudtoN2L5ZrQx2QWWmN3uVo
ccAHC0a5P9qcnkVE8KFimdLmmvcDVwnQMop1E5WpTHZUJhhPso6XuBIywDN/63Fp
n8I8IJ50vInhhEuobFxutQ8nEnp9uPA5JeBPigl+3uUuu6BcvB79MuWaGuE0VIwA
coxQDjHiM1BL3IEiTwF+tdt6HSjLtAfhAUJMQXuOI6F4QvUwj9yaptGR4lepTGis
Y2ieL5mSnvMsXObnQUAOskMvwY6RdDrGBLNFpbCE4VaNhUg9c2IzzS1PgEajwDR6
HNn/FJsE3Fi09aBJfdRnOBjY1vXIMYrBDBDI1kMc2+QeFyzEv+rqSSZSxKniDnQA
tM5ptMza+RAjWcvEosObtfqVhObIJAvOHR4mznysWtwumsZAdzZcqZsEh8XHztBu
aqecgD7jeMR4YsDGGKSlJmxvxUZjFObRuCS1CK3qSsKX+aqj0DC08n+h8ZBy/afy
PA3erOJECszgtcBgnpaPScldyjtoluRMmPIuu+7hcQVjLB5EFJIMTupABEjQt7sw
yzkx4RdO9dLjNLCqrOQIAcxny9CI9D19KKWpgAtTjWmqw289pjGnUxb7rALfN8hU
/whf2JuH+6ys2E1X+3XnBMZWJJVkWlsFB0euE7nO+wlaT+I13wx4D6RcHmVLqqXW
tnfZPSGKh9fWcgyNt+a+dw27Cr+s6LPJmHwZDJouj37fz0rkvRBaf+Tr+To6LuJU
iiyt/Aqt0Vi9Ox8HubB3kQ0ftFwdsbLsD0AfMrIMvFs7RuvtlLRGXczhY7mdpT0x
c/PRdDPexBzL4ReIzxH5beSflxJBzTLH8Ur4rtOwwijnVvEA/xy2igjzHEQ99ZKV
EEQOfAhV8yodpywWp8S9NLgLj+l5dl9gYuFkgjCe/IrrX+0cdDcJ6ZS8BgeErmjF
6sk09QujR86WP+M1IMcU9JDHXNbxL1YVCxK8Kz7lm0jhlE32F6CRwjCuF/u4w3Ja
KxGGnx2AATYrW3YwCNKlQ3FMchy+cDJY7blz02UElxYibpz6lA9CzBZy6mcL8TRG
YNWTAV6NWeBd43IwiSzlzba08f+RifWdpyDu5uLcjphLtgfNYXCyFYIBYRuKZjm5
QUMytjP8Zsc2TMC/EDEj+yh7kdK6+PYrfOQ2ZeOWwSrmSiLyj/tHysT35XTrpI8Q
uFT1JqYP/2wFwJ0Mn+//OobnVmZT6wyLuNFcaFQTP1MFVHv3wHFWcxWnCGTHr4a0
XzuqOxZkzjeHrah8brG7jQlajdkVHFnxV3VFN8dnsRNKEpdTSFVL7ue6Cu3binPZ
kbJnp+54M1uxPPlBV/3j8PM5+BNLEozKaJZfMXIMklD2qrt38DYrOYolmIBns5HR
7OeYRrZYsuSbBv3vD2/vCEr+r3Kl+Q4Fdfb3DxHrJVs2SDkmRvZm9O8ScpVk/i48
gMEyP4i/bcxGByIUg/VaqLedT0v5LBdSBkRKu7rqOAXfyLXUZ7PeFwqPIo+oHnqJ
l8KN83iIMwuhdqZbe8kTpXTN8rRjUc1+QjNh5DEI3N674JeggR9nUUpUDwoyNKRX
ImYulv0FvHyPtb7tzCKK0XFBfVnqs5fkGsJOYLkNj2HPTGRSyHbMf/Jwvcu/KmHS
kHuZo8PxwgVauTkzNkTGSxz7AdD3PBkxMRuPzmtR2f73L2qbo266yqHRlYZKXTZi
wY0P+uUmxZCB5xs4tjd0VISTyoAtDuUKE1dC1hbTc5K0vdPQjsmJT4Ucp3Qevna7
SIiXJLTZRv6+0P8NeXJsBYsQ7HVLv6ATP5Eh8a2g2oaOfywCN4FA0Jv5NzL+smgE
t0lkIFULM5s1NRdgxZABMWMzFmbo9MzLdNOgPDaldDCYlgrg95drNSy52maiuA86
R83Ry7rmaOVpZKr9MqbAuyXLj++VrPuWXRCCaYs4Z2ZonpCr9GM6vW6gH9eR1uHp
i9gZKarDBl6D+6LCO9jRfKj0ZpHyJBp0Sq8/fIGLDs1t9NnGmdTciH/v22uY5ffV
JPw/N2XA7KrnRy9rvcL/cHqZ5WZaoBJc74xj81JNu0j6GTgF1wl38mS4YQlbs9+h
JD7/Rfh97u6PMtyLFdzIvSfa6W+kp0gTZDtH37X0u5aCVbI7ta2GgSSfNvevpU3l
wS/VEZz+EySrG6jp66m9rSEBrIxCRmU3rN+fzfwp4//bZgXzt6G4LtZaKG9OH9ac
Urn0eJLYRKb9mEOB2TPe5BtCaFMMkdDiRycjf4yd+y+D8aq1XCr/2aNmNY1mcpEk
bUMIi7GpE+akIEqF0aBl5Rb6wbL6w9noTzF/sL8YE12GzEO8Q7u7yWKCGl/Om18U
wnIyNfj2cYV/b6vBZOHe5olrAiA4bUXq8OUldQ//xRUahkh56OFCygiUP55MNYso
X1E7QQ9c7UqsZSw6pE35Vw+b7MjWp7Q63GTzonbswboLvNHlB48IzD0ciNjDn+fP
fBqN1Ai0U3Ktu+GKcDQdYCvO37fKFMGXwJAtZIyCbYEf4Y6exXqsAQv32R9AXq2V
KR1RzpgFHye6pkbSwS9xOEybjt+dkDUG/CZiZKav0UtWytgRYOViXb/tvntLDZqH
QlW5P8altsxv2JrJCTH80dCiBGtpejadLetn+iw9KgHaZXXI9TcE5vPpu4ihk07C
D1CrBmDyJFCY5mRwrY4XN89PU0pUdhAaGndIwsTan2aQWyeX+j0whiFv++FVdJqV
FE2O9Cwn+1qVa6GWJCfxDRKiOkT41RmPZX63+warSk9is194I9ltK3bMEXW+aWLd
ftxhEaAXButv+mHXhXU+uZjG+K+1Wv/VLmMfrP+9N8CicbflikhHKqAaHEwzR4pe
eFuXzGFRwvFZOWDwVHT0pBnbSZmcinYxCHoVV6ut1bJIsckAIVkXrPf6VqxuEjhn
SfPcgqhOOhcAo+g2dC22r/gx9YGpNuiOS6laUdfsA0rjpP8y/G7mVUkX2VOVj6Pr
sUZ0xZWdY57+ls7ydqonGEvwrzUUrYAXOaQgdRD0rgQz9nfWYeX/NPzXCzNT7SfO
kMLHIyN9NA0nIEJU3SBHFfEGH6xW3KmB8qZybG0DaZUeo0fZne3WtU2qlufvdHkm
w8GEoDNGIf7HfR8QWWzw9qc+8ukjkGREM3v0ewncegpcls+661+V49SpBr3mdRRe
5o+VhBiKcSJzdr5dZxcH4AfAjRwnXXMGeXeQFwRZ2sLRgT1wk7WupL8B1h6FXkqX
DPxr/HPXMsox266wF9VamQKvILyf6Yb/lQIXDcFYH0M9lyMGgKfpNnp/0SjsAKyu
DSpBVCKwY5o/w5XS1a3c1n5Cg2gcAGIYe78Tc60bkcbG9pkIEMdsxsRew6M/KqLm
Rl67Nxr2HJtd9RL+GdbBNp57TC0lw8P+7D/4Aujsr+XecHNt4N3UNht569u0AU5a
YAqZU0SnXn9TF2qPjpGAMcAWet8GR0V1alI9PsNDqUJQi4LsYlco7ndOtZXbVYJs
ePmd7c9gdUsXVrEq+TYAMuwsJnMWvRTsmHHXgwy75L0T5+z6bH36xRA8UgHF1jmk
A6jjEurBDjLilxPI5Rt/A53+3JQmd4B+a4NDN/Tp04EHB/XXUo5pt7EmV7nBRCG8
7Vjp2n0T4/sSme19q37pVZJ/ohiUY3uj4+/su5o1wJLHF0rpr9mYQxbby0X7U5/x
eMcvP6K/U5ldlBp93O0tW5YglCEeSpm3f0P0lIAoY5aL7WUTZ4ot1zBcnWFCGNAw
6s+1gwKk/LFJKhczNMIziVbIQeJWyh8JiN8Erd3GzMzMpPnnFngeB5xl039Rc9zx
PhIOfju6r0ZALHFvzJW7nFpDAHAfunXEmqwwfUGtXLTsIdw1lsDvIdZZQuWbEKFd
e0EOL/QgCNZVO4MhAHBN6Abb536RVw9E2mgIHIg2CRVduQRP3kCBov9ePprvd2Yo
MOdPtGZRwHuc+nTy6eLEwRdvc7gSBTXlTu3PhJQbq+Cuf0IF4lyTuU729zXOcwGB
MzGakvVdr5sECD/aI8cAKoI8w7Vae8OSjns3CkWCY7ha4OkSrDzyvftoCje1Jy93
ZQh/WwS0UHrhKkbgcN+G4x5t7ZrHYt7Fysu1NphYLSLfiXlCO7dDso52fwCWzmsw
/ueTxdA+ccgnTWWB01CPYZnGTiqyeGDTfwwfLw9zMCSZ6aXAaeklQ+UU5Oyjao2z
fCe3jklgDc3GtUqyjN1ihdIN6PKwHvj+gGQsq45KYrLPUf6rt5IHSgg1OJoiV2fL
gOaN+Oop+AYDAN9sO5UB5921WTVNcrXwVA7azuh6+k7W8aesf4pFQ6sLJdIf4lcx
YQsVclkMB6ce/ccTx5bYpLNJOM/9TpFnaUn4s7LLPL9494w5/OG84eVrtlq/qu+3
lXyB7DRmX8t60qGdsl6PYHpSZD3FJHv9dqWGvTXc9C9NBQbIMkLoFZrl068eUaln
OOq6kRC5DkjorvWO4UzyjAfAO6kdLDPMgfFQ/aKqLwPCvxSzG9eyC2XVNT05r5co
yI5stw+dHsk/uOIziKl3kvhA4mY8iIZOsexcP9qvhV+w5zTOr4ULeQ00Gkjw+pSI
wBxeieiU7DBzlhxzLtFoZ8qtfMOaA7vyljS4TL9iHIYVz13QjMscJrv/0JV0QtNK
oTwEvqehDUhA7NYQ3gz63SY/O1TiAC30TQJ0vqID9i7ZFSxSjNqcxGtk8iqlymZz
rH6Sk+vUp2dr4y+25mVI3T7EFFxjjCBt3AdGi3fAX5r+DYhgMHEGxFAm+iBN9Y6z
6vvlSGc3sLw2PEAey0s0vqhmiQJ8dXiqC8Oy+rRK8VMRNeDonM1tvzRRvAXIHar/
IYIEtHVytx6gcO1f3aFvr8k23CsTXKATmPx0PV3pL637VnoEZbie13U/xlH1s1dz
4dfDmP2/Jt2FNo/Jb7SAqXXd7YGQxNJe8kQVV/hEmfugx3r7jl9GhXLNjALYk4NY
uP+bK0fFx9nGcLQp48jj2khO4BgmfhBcIPJPC5iDPRRbyhc3qcJewS7hZqFLQY44
DR3/WQNcNYqcolcXjaleEiTo5+j7ms+RfQJx+Ap9gRixM9S7D/miYXeMltdoHpCS
/Y6pTJEc8RSdWq70Ki/1BH3mIjU8ICr024f6GLAG1QXWctfeEZj4Whvup1PE49LO
i/wV642e0vWYIqK+kdJr7S6RL2yNBJTArm7ahY7WSvVnHEoegnW6NmFL98vJzsTQ
yfStLX54VBs25503H0v47cPgPSXccOqyR6TmaqDxVseP+GON2xakCxRbFjlbP4fz
wafryKwSWquqqQB+8TU3hkJEYw60TPOVNZnNbPUdwxqYoVmJsU0rp7LWYdMqEFyW
koDxMmwDBH2NXLLIfXnWX+w+Fuu63F50yWH79HZHATeRKOZ0MMBZLQcJgC4PaGX+
ph99D8ZGAQPjVwTAEXeqxuoJkEHkLzCK91cdnirJsBwCrH51H7AIQxgA2ejDeKpZ
GIrCx5EyQXvC9P3rLrHj7PDcD5gLUYvfiZppXiwrdi2OcJm8m7Q0/6RE7CkbGUiK
McvmMi6jDmb49uL/bGKyZoGRImXoV6UZ9mj8dhJlHYxH78D+zIHcbyJ0U7f1mvF9
Qaxwus/6m6iELNtNQD2pLfnvH6vTvzdCWJlGCpVcKjMyd1wNgI+lvh3+UaSCyxKw
jLqu+NBZrDTwjSYzcm5SPb8c82xEFLn5L4VXui4dWJ/7MNY78OeZygvgMwibgb1o
vqx8nRRyz9/CGBlGfXZ/AA56qgA3dw1yi/BNvwsSrowQWoG8UuW6gPED8MUwOsIQ
3KTpyvCijGzlXO6CTh9e/LOj1ZPO8OY9iH8rsyLGnnsKMuy+xLewczagNwfGPGlm
+F/k66V0KdqX4OJ/p18W7E5WmqxITQUC2zr6RTuoc0KfJ/Gu4TeiLcoqxe8XW1C6
Vq7pD1T/EH0KRQJODkyGcrbsPONw6gePYusg4ntFdLPaGYVtP/o2yyxHwipu/4/E
pmMIe9TvxqLdIgPEA2AaKAFBu0+KStUhd5yVpXL5IzcILwzJZEuxtwn4mDNYycgs
mpwERuFe560YkDLM1jtvU0yoJBNlMyAkeI8HENgnTpjuBIX8wEkzEiZrRy+O+3pb
7cD/5EssMTdAQ7EzWilnaTeOWjEw1ACnOcUF2b1JbNhhfZjxZR9pAQWEL4PQQcnz
pC9Xu8fltxQQbu/O/jzMnRLAMc+wqnHZOOWeYgT2/mauYsJXFK4cjdXs+VgTTBO3
6pQBW+EilIMhZDDnKQzbAWfS13e1NWvpw8ZH1m3GJLnepiprpnopVFeirhmcr376
qyMfDSkXXJcdL0TH9PJpt1XCLU/aqiXfP+p2lIzjyPjJWc4sHFvMPTm2D1P5HWvf
7OijNx9pCGPmybYYGp9UN9ZAbOnAgbREB0jJymU87Ta2j2krGji2sg+o615StUu0
XGacsXAVDplNhBMsrPMy7w+Fmn3vuNCrKKtc5LUj32lqS1y3cXlrA5hW+fXHX1gO
x/BcXFZX1zlBwyBn9HXXRLFwvS6jRj4eoLve08ndFwmhbPtuptqNlgNEHkHoQFPE
llA2xa6g3DtCPGzFA4BNza70bO/pg23d24OLvvN49iGfSV3n+C4NzB+BdVEAr+Pn
g6+3merc5ISrjltEM5nrPHrvDcyTQoEoU+eF/UwmHBjr6lkbIv0wtqVYpJsNXs6r
B1HQZZpakPjK7F6JHpqHrrKhpaKoBGou98pNjvY66V1FjMKH4LEZcxrlL6Eo+lO2
b0TFq20fRJjMAvBe4qa8TurZyKi8DMkqpTwqYhR6JL5k9DSCtHvitYUtZPCvwRFz
sI9wSav2zckRZe2Bw3g1MzZ/z7laBpwzMKBGGbKOJ80Qngg4ob8+mcVs8XcMu5qu
cwQ0f8AMZ/GfAi1E55ddDIzStIH7p8T+wB+cQJC7Cy7q/+vAnIIN4VOwPAAsD8Nf
aYtLmERORBfA6+G+h+nN7EEZ1gRpW14eNINtbhmiHcNizHbHmjod54Jh0WY/bCmR
Pkl6YhqnHqCsWNtCElOiWOZxLItPl86PxWWeUKy5iVJXSy38xjoLZqF5Hje+vJ9v
h8EmB83AlATF5ILIe0tztnGu/xAiBp8sMenHlxvzzrmKum1jXC1RyuBTkl8yciGc
kqFGA+CJd/kjW6HmJA6xiYC+790PkeX0eiSsQpMAtie2DnGCKXjQj71Ur7mxRl0f
FfV4LtFVxEnrsuXegd4cPe3OQMMTLS8RE6P41s3V+TjRPWqXs+zOmygLlQyq0WbR
qk3a+oJexAlGRuc0I9gdT/B5ee7Z8Hga7lQG2pSLBADxiBIV1a5w9BSCQoCWe0Lq
stl32/WHSWiQqukztNyg2XPC4gHoPKBnMwj5PjnbFwFkBKLNMR1nK3ldc5kpfJRt
+vfx6ezqAPJ8dNtpcP3/mdMZH8U5KYGKF1Y699p35IcGs9YH9/2aUs3/fUW1Jsmk
hO2La6RgdQcROocIiyMGWLDBR0E7TFOKtZhi1Hw/YcGl10dR4bAIXC91B6utVLgn
s6DJCG54XanAfQ3JWA61HH3MOqPXvwd6RbC5IgqP1xhaNi45RpEbDYNHXKpBTJEZ
BxSEI6ESHIhIB9b+6l0mbLqZICLDhEzm6oXdPTaOIE4tUBhWZFIglz6m/eXKF7kX
uYstFXNLckrmZ//XIj5dLESe3uSsnsSAOS0QDXEpT4OQoO0Llo0yMQOdhXNqoga/
erxexsw5NmZ0DXGbRX2U57TrD+RS+l79JgiYG8PMUr9fyN7+k1NP8YZmnFss7SAk
XwJNcHyXFScuAb2/ILM9XEc8RUF0hhjJBMjWJUB7+ly0MHAjsIp53wHUYSDmWmUy
2A4Qog5GJKnjj0sLrEselESA5SBsTCw9HGOMxyjPCqc6UmwXgz18rhIA0ClKMf1U
Y69xXE4/+gN8qgFM8oUQvgYKGlZ20/ptpABD4/EBZjb8B5+30j7udvibBWrCXhUb
KM4F/UqQKYom3hwgSWWbzEwsm8DgHr4GlUDwgOCLJ5q03GKgYKh8hGShs4XRzcs0
pqtd7Zzby+vOYyL25+fYzcXiA8Lm1G+peK80DLfR2wHT0lkTgaRQsnlX9SqMG93Q
xNRbd3ZPFQdQ36xdMhz903AWkBGfOJItLJwSO5EZX248SYcfzGWIP6LJoGDa4ChU
1I2NPaAAz46fbmE44tS/wG5nVOYPQ5pAJ5S+r13y11eEFGQ1YXzsMt8TM9kAi331
7dxmzYcdrt8Z7uML0iTouJ58qTTDKrmSQ2Nb9+DhBXvgoxa6i/cmRgiwOeG1f7qR
dFQnZlt2eGB/6k1fpNO9YeTjJ/eW1u47SB/3j3yLm7q0sUY+FAgM6LSDA/DGL/KD
69sBKJSHFY3zVWdgKsYFWzoXED0aJqJBWLgyFTZPz2Bm72Yo1HlwQSP2NUW1FcRZ
PZQMmNmo69UKYxVnZsKPIXFQOvzpsJKdZmVOELdWrFq6X++OymoMqm6kCbhN00zo
U+8HWksUJswSWv10L/VFoCWrNptuD75zwtmj7sd7W1XQ7gu1pMrTsI71PtGSRvod
UMLmqzTlQFqQ++3AsgPCq2bpmMGsbu5vxD+DeliaKN++vHhxX8wYW0wm4wYiRGzB
/r7wyUJzz318qfZxq0DWw582VDV9SRt6nvcrX5BPbHp54hfXZYfVaXmcqBD6pht5
aGB1i/H2X27shAAl7mOag8jPYfyUqnr3gQyUU8sklnIibR03iyHX0O3hxpFsa3xC
tsxPmFoPUr7EKzFAbv1joMqE8lr6RUtmlQ6ZWwixQbJUsawMeyzZfANnkuA5NHdn
2pLTVJWb/rwUe3SAUK5z2vcESO9rjZ8TDCsN4dCUV/XCAcy8g6QDYuMY5PyExsiH
zLE9iNcHprec1Y4AgIldU9b8Rosh4nHBDsOWOVbbepk/EusjLYbOvYVw5SU3LeWa
KTu/Wf6JR+dbq/wyNRw4TLI8DNT0ybUJoVBdwHTehcX8JO4xFrnvM9qhMbuZ59EP
bR+c1QZ0kbio2Ny+R5nA15+QgnpQMP8zlEhrWTBQ9QBwsmANQB6WrYJ3RJfl+A8y
5N8ezdBWetXvrJ6R+qL5nT6i7liu1B9a/Itu0Rv58G00Q3zV2HujxjgRSuYV5bNA
PpfKjULsDI/6KtCyBR0IHqC/GT/o+DA5UBrsiQ+ScWpKms3WOj/c1pWR77TO+KLN
ZF92L9gYJZ9JERIjAV8igpqwmuRsreSdURJ2ifnhiav2/VXJ7VwpY5p7S0qbvb4m
nUMHxuko1ESrio8CpuBZc+5VXQJnIAtxpjJBCYhrnYo8O+zh22g6pUnYLFuji3IJ
WT8Y8C6FDh7g3AxN12Eu6i8Ra5Ha3xuC9u3blSmXamkpeuYyqt7KtAEMWWT7zxwX
6n2bnFS7ExneAhEakY4gcI32k/1fL9cU6vLfM+FUcRpQ1wOQROf052B6CHrbqYw3
aYylcRsr84Sf0bMJBPvXqZTgQfXPGrok8dvZBLbEMGsPBtn64YaiWee2QKQF8VUf
s7ESZWu88TkR0AiPPKw4ZZu/M5WEbt1voEwOHLHRAYfRlxAYv6hJAoYHTRDKfdQz
vEON4H6eqauV7vvztSBo4aEWsFwJ/AuxNTlDx/qMR6bB2YmlTj/XVZlcZ9XQDeoa
zAyaJNICoclKnXjvIS/JdfgP8nvLXQNSICDqQSbDsmq4kXGOZJ+FBLdf6pfwj2c6
Dt0I1wJg8t60Y1Jy4GdPnQlpw+nrcTRazU4toSQ6dSfBWTMmbOq8pRMjAzRS8jQD
vRzghxP816wkM6ShEvTBIdBdQmPhH2HYDNosYFp5hxaTjYbBz+XNU0bO6X8swM/G
FiDM5H5EdRt0wdisVO/wt94/Py9eJyuvPFFwI2brVipgqMlO1vtH7hTkRziQASDR
gCxDPbmT1padjBXc2zQcgcqrZULk68o6zSlKhgEHSffdBvIDfNn7uBaXi2IbbkJZ
3eSnNUKnImeqVgcR5fTJAt3fnMorTYSTttKyC8Z1W3I/MEQrDwIxrN/BKlUret1F
REwx6TF/UtN6MtSQRT3JLzjlCOsB+2f/ktNXu8Ln5VfurtIstGbFJu2E3Wzhcqjh
uDjBUqJ28y6YSUZ74u6+histvrxNP8En9A+hqBhpHLfIkD13/skyQxlO8dthSfwe
0/RqjlM4vvSvJJZwaYm7HqBDkfnnM7rqPzHMIIFXB8+8emeAuVcI2/bmWU49uTr3
HuxVSoVlT4KKgedKzz4ygYzbGGTNy0L7Av1ITRpvB9Y959Lwi1sMgxwEAZZIsAXx
e2yJzEaY7BYoEJnYMzgLmQorBG8I/Zi6Mo/OHpTGRtpaWB+ojhNC5d3XFoiVRnHT
zcTZuqbv+HdkcCSwrH3zQrT/QkDJPi2NpNcLKnygOrxnlnCn2fYkhXNZU+K2DDBm
vHoJX0j86SLiN1heuat7xymxqHNsgxqGLgupnC3T5yghUvKgAkb+G6q1PCtEeDoi
04HddgX/l1SawkdD3d/3fne8fksvy+tHVTqRCECGjQTdZN1OEzzGRMJra+qDkrJ2
MRh3qG/uBNctT/Th+sbZqRkj89Z5Gxnjm8rlHOJpJCxvowHYeTEuMBh8lv/0QxhH
EETI2Lr0auUdVyq1cjqVhw+JoRV2wCjitPa+GqGeNvAjcDoQV/7q9LY3kCr/+5s1
6d9CRYUMY858NmPcSLFPiS7lpZiZwxBbPU8mAV+GTrlTJYXaZ8IAF+P81A6ZYpnH
W/7ze7O5apQwTa8Sa64+CEE9HwZi2avOk52mMb7A7CE7qk0Vkp8p31t39eKy3jxu
e+1UfjXQYQTzbzpuznujBqVn1Jpg8EoIFtXQOGFZ7dwsG8W1ReO9ZK6SR7//z8jV
Aw8VamV9UOB/KwV/W5xNDBYfnbPGGS1D9CnGY4TH6/JP5OW888EmecindAQGZuhY
o223XodHxq8RbKFtCoGveS5vFvTodH8zaT0K+GKs8iGfBHci0cqhvizAstr9mw/T
6jb/RlYWlNWbLAEeiBK2JcrC0malVLEWxG82AT/lzCAudZYJUHwg+5hv8Wf7zJhX
jvB/Lj07S6CUIWc3Sla+ehqpHH0DDdT7hQKWEkKFS1S9YajBzb15St0eNUtaIBXI
zoYMtqvfjG51M9NxPJMlLorucK6Ot8aM1vkTC3RwPRCpq/G/28VCeuRDhW2bFHZH
qgDNuT8Z9DABnsAdjsweq2r45tiRgcVGXja4F7Lx5K3vQT95Vigd4XxMD3t3QE7P
XSxZyXEd1oxdf4t5DPTJqpo1e9gY0vVZrXcrIqufwL9xmVvWi+2PplswjmQjllkN
SvdaGgqbOHiR6EOTCj1VeRW6F1YXR8j9GoORc883VRxZtszCsiFU6evxYivdxVsF
flcx2/hggH1ynCk+TW6SOijSKr1ZPekjoQUcPyx+Wt4/5aovAj0QwHf92xCpE2LQ
eIxCPDnI+LkwuXr9i3/ZiGCDJ6uqjqTMB/yKtHLguZpWpueIYG2WQE9nRT7WSzaU
IHmjrDnpzuDLET2nbSbAMhe4dLD8UuZNDvxxzuGzO7j+A7WygIZDpq9B1WaQGnOO
njSGZ11ahhrN4LgKE6WynvzVdoxzaOSO5s9sO1RoN3Mkzu3UloXB0vCLaIfze4qo
z0Rirkz+O1G2Y3YKNZoFtw747lEVeO9OG7lHRoCQ2HOf4kCa2jJkKWbdBZM7fM75
ncI0q/tn0wnYp2u1XF4ODr+LsB8toO07/GCkRMI+JTllKxH38EqlH7v+fec0EY1d
ecry742StI+GVBs/y/Dwo6V1BnT0FX0FrOtCfghPgQh9UkUpLdKPoe+a4dDY/uR9
YtnpC8PjPoCQ4rmUKfmotodWkdGKi+Etltho9h7f66suf8aHg2A6cRdL77xtkjsp
fZL6wqKZXavHfy1v/sXRI6GVtT7jlMuWx1nlipRMvOily6DnqI5txRFWdjaW16zz
qRrTluYS3lRTdzfI4z88JzPXyyTCfRak9sBtnud0pyRIOBbD+HjUGM8Mvlvxmf4I
dDljH4hjRwbrHGqIuWgT40IFib5P6Fdmw2xeLPu8F9xIHjmIHYTig8Rpvnxlvdag
54UgcBlwqCsu2YW/3vHF2EzqKTdjh3QHTN8XK96gvCBS1WhJ1txmPw/KgjZXJNgO
UBO1xkhuhFuOh+YqCbF2xAr1iqpHHFFCF62q4rkT9vpHBnqAi58klsV4CvhCjyne
cP1ChjTsDGaLqIz2ieIocoAsB/SiV+b4pFaNwIq4fVBrKEQmixZ8f+dLUTe14TJU
nYywHoOC08eo62chXN+MWnjClq+0OLnYJqKeuzjU4H+SyIutivyJu+Hvaka1C4iy
b1Nm1Mol/UMtdVbYIDpnGFkTgm9W5SpNcv9TQYWijSeFXvlQbkXtXnN1+8J6gsRJ
n07fwuGghJf19iMAlig1Zq4M1DLRwJvbWxETvM8PgugGjdKGhKThAlceziBTeR+Q
fD9h488H5ZuIs8jwDnSn/t0RzN2x1ZkkYAJbMT9T0m+cwuyWOMszoJ8ML6O9WLHt
4mr8dnie3e47J2jGuxH1x0bm88FgoU9alpcTodfmgK+C3oFqmB+GKjyflKtn1Lbj
umbKiY/DHDvYKyX4Q+U88mirHsuiNFxdofWQAr2lB5sLoVeUf0K47bRXffYz1Zwt
n44RXBkR9brmMn29VBYs32w6PdOixfutgXph/QKm4HXCk9kdhgAYk8vSmVqyEOtI
PuAnnhIrMwKQle3Unyy4tdX9qO8XqkNaRkiP8y3ULS0i6T8B/qdqIggLUqYo2dwo
bjBd27KR5PwidHQFWnS8Fhq1FuVY71xylvB66WjeBBPEk99/R35lJnEu/Ei38qiE
dooWvyIq6o6F+GKRWcWWPgbjTKcfkwtlbr1rn8MyWwzgtw4rVCaIs/khDDEiAAMz
BfsSmJqAgcpENUSXg9zrHZlSwZhI2nFL02gMuDgLVud2artW4LfZLx3ARoW/2Cjg
w6EZSkom7g17bMYE0bWWf/HyJOkrJ3NWSaAdouMJcTKzasCDwYGxgKLcAl5VAZv7
ZKwUq26nLzv8anXhbJpt5FHhZ49aeyWR0WHUc5SQNHeljlRNKfEwZq+oOAlykYwC
imGRJf4Am8GJm1USvmxoqfEe+PqkWFUQIqxXftHhAoNV0jrJOOI0K0gSBAbUR3DS
fmbqbuoc/GHBjSS456Nuf8FslrPdpJDKu+mXqbhrZJd6kMHnG6q1ypLZiJGW/Fir
MJN5wAxL+VBt8ZXeipm9eN2l4Zcn+bIm6n0PP10MtWW6vF3M+1P4sg1SoHGVWNO1
sUUYZVDVQurOZy33lTcDz9EJREJHMB8Qi57G2iWwKEzWu/GeyajdojZjdTXvEpPw
XzS/4cBbjjMuJ6zx9XdQ2IpIG/Nh29BcovK76TvbYXjN85EiTZ0JSXbSAj1ZIZul
3MjPxqMnciVUUC2ERr0Y3TZdFnnsOmCPEiaH873iBFRLU/t+2woqM640pml5fCiM
euMW+G+DAWtUipwyUb4WZdCOnUs3sEu3TA1+AJGHq9kWNODTlEUH+WRY2tdm0TPa
yCFwg1ge1gVqHsLNV1mccBVGn4KwrEc86ibj6JCqrT6CE9o0NthYM8fP3XB3jYbg
BSzjxnBEug2t/12CQyyspJjF5/IZIAdI2m3w/eEkR1gm1SUauOCCbDv3aRSzCr2E
w6DNRS67gLvQe/9eQTHaQqqkYWLQSuIz9npObpAzuSf7s28DwZ7hvLCEo1MP5pMw
cPgaCrGKsJzTx+09mcaq4LB4hWMXO/yCMUvw7VpBBaBUfPOvIefGHR0pPBUMNw9z
R1hOGgE/BxVFl3+7YMQrBQtrj06lzJcWdzSk/f7O/y2wVqZBGvPMNvTnqHXBcm7R
eVrhkoaKjyUgEC02yc9XanrvCYUItJ+0RxdDp3/KY30w72y1OoVF4LmbEfRZYa6z
TlX2l/FJyo6ykhSjWgjxkBA5mook3MIu/XVl5wEfILMqJvfbmAfQZRc8GOsTUFe4
U1/48ovaOx7Oqkyihc+dNBrUovGezYycdcxV26R4nK2pm+e5R515LmmOY54ODXVw
tyhwZZr60KIpVTV/ueL26V8naTw6l5IWSmiigfJXZW9v5GOpsIrWssYid47gFANM
ejqT3SyTczkgdXsXkVw80b6Jwe+BzjIAUspH9Nyj5bgZoEFP8zkvfym7JlqSSfKJ
9pGdvgbMouX0WFJK2qS7xaozSyYqVVmI4vXBtC6fcRGdVOJ6fvOUNZcXPbebN7l0
hdMQxvaEPt2sy8jlDp8sGyLvYQXylSWFXE7czH5wn2ghtGeTXhXYmJ2vzH7uMET8
G2f3B0jekgoG1py03AJzPyIRso3GKeHkCs74ka3gQ9ieNUEEUQXW5lO5ZcT32BHx
SlFEjEggwcSxbNNyW5wrtliI8VvpBUpVBc256koLaf0LA8hzCztVSJEuv1bVUmAb
f/jeL7apsUgotqrbnQ87E7Ee4k/D+RGQep34BsyRxf1fRkc1qMIR18xesi7DkSV0
TnJ9fFz2Dcx9QyI5WEvasDUZZ2GBeIn+tea+uhNpJ205/EVIeT9D5AaEx+D4tDc7
WqUHvUTFXgGiTaRi8ZTYluXbkHzFcWFYzsSOft83Ndt89lcRxzJrZs/bV/Z4Gbso
MOexSSJVANxtHdeTryexIJKbYD/gPBX7RuMCDo5tiRsv5x5WtBRgYHPGPxJ5hDqY
pI3gVQ1j3s+UqGtdbksXC2qsywbE0xK2VlupPHDEUoveXr68GNrbbtRldYBLOnRd
2UNeWuVjKYdifBp0CqpUQIcBdeSwEXs2OP5yUfbT4bxUyDbUZn7KlV7qF/XR1vHS
6vVE0ezeqURy2Ewo4haVI3fbdhNkDJ9aS2sHV8jWVNp+T8vyyUlv/r0AFAbyZmrm
8g1Hc/10XPCVO6pCYEB9jDx6xd0NFYCDTrE3VLedVYkqxdJkGwf1tPF5CaSjcJTL
JyPHcbZ9CMF9lb5wAQx28Kf6XP1VsMEctWXVXqYn2UyQ0Aloe/MLlL6xH/myw040
aL6bgSBfxTJV2UNVfoZQFeHXZf3VfIXXzvhyznebAdPEg4nbkbVPE9ujk0R1sDFq
l0m/wBHanjGuyJiUR99ZD6mMzHQkJlQWzzXnO8gLJ+y4IAy5oHlpAR08OCYuTVXW
1hoZ/vlnemKj7svXD0hv2iZxeEPSkDIAkrCyNBOwMrXHJIoW8CoWYI8sIReFLDsI
dCqrIPfmNg8XcE2SVXX+4pZTDJ0UU0tEanUfOV+51rz8tGfLqaJaQkDzQvZJWB3Q
R05rdrLSG2dJx54mo2ZS/XeSBP9FAo7+3fjmZt4Ne1chjbxsiZ29PWd+mo+i24Sq
irdx3YKBHYJuCJtONoVkATgeomS0Af4prjnWeGXefPSqSlVCGCNbmirp38vDAbwY
9tN92e2wrCrnSuIMQaQfV83Sg6Qd/gwI3NJLb5+lD8kdum5wmBV0biNFHzHh8mkh
gvFRzIuoXIYUQyn/E0eZv55fk5m1jKgInk2swj2mEhtSJPQHMKepSAKndiipCWO9
273VXglmNjhUSAj+fvkThawyaqk6PB5pfeHIZ5wMZz6SbEKD5ioTuXDD5cY85qvo
8HwRAwScO0pS67j/tCliicQbNIw9vRE1oz+BDsPOP+I/ALo6sgYB7E5jY8B72DB3
pl8HhTHRu0cY4o6uj+JpPQEb5GQ14tPpDBBrdHJtZGNoVB1CJR9XS4Yudsd6V49o
wrr1MtXLr8SMIFJNWAX9QuxicvXbsfEpoD8PXXV9JRNzQekk83AwNgDkD4R5NgX7
370U8KJ69m5ECKAVmtke3RtFbwlCOMxpMY/LGJ9rMlHVauyjRxYNIbWSFX4P9G3G
wWi0rNDIw+SAuPG+l9mg5Wqa5bN2Mz46k4XkMjsZt+CwpHu40K3n6SHJLtHDCbJA
EKvYoCAGI0M25t0AJMLlpsKsLSwwukyqVRzcbeLuerWaO0jcT3dzh3UKwnezKEP9
1teAnu85J0vsIMoGg/7PBYgJuF+HnlmzkmvcZ/DaqepU8ROfzGKv7+Kx10ZyTxah
7/adjY/QKD+H/oqa64DX85plV+tlFiVSieuZwT42PwSrnFXsmurDgPQug317bLqD
zscvbyx9PQDrh5khX/TXLl6RE0gefGQ8qKhhsIjkPrw1kPCZPl6JT9167mH4LJ1j
T+4W6xV1pTVtFL9S6EpyNyhzbL1p9EMNxEvcs7IpTFXK1wJg+4KCY5SSuVU2nHWp
BQfAk72zIUYeM2kMONkAza4bdJsbLy1GV1EAnvgLSiiQgl1UztTsoUJTpBXrPxkA
qzZKE79OW1GNCv9+Rms5pPACWhxYBR8BIsNZdTs6nLiIEn70XS39aAAa+44lJxGq
LClacZcUqqbe6NBRPEUDgD3TCfSH47WSF8J207AhJx1JlOVhiQd50IReihdTpq3i
V4PK7ORphOebyI3qRznm7KD1OyJHdtYKhtxiZmmMlvYaeaUgw6xHFQCxUuIeXpK+
9gZV5yen4/I1gUBfjiw0evzzEOQ0Na+dIUr8Mb+MsrsAGT4cs8z6Xq8A0zKvLhYQ
/KMnhE+H9JmZeuPPW29OBM6UiZ2F8mJ2P6tC0vRaHtl7H80xbfP5RKjllKSHMbX2
qojVuoUE+8snLsrBIeIKqxfLCiR9NdoDieo/I3VxSH/oxnY0OQa+HfrNcJek+dU3
dWHAX3KVo9kOhNbQJ0u3TM576W6kbIao4rWHT8ZoGH83Jpmrz3pyDGyymEuBfvwN
KFUnM6z4bPquzad3dXAq8/VQv8CCpw3GTKa4c8ZaAlipPvvi9KviU9GDBwi9XUjY
7hbKTzo1eVhE4e3Lb4XS0OxDIozXg/QPp9nmcPhf1zMddFLE/M1eSdWKg6Xvxr8z
wZ561JXEfDoicBU7kRBSvS94/IXoM8Vm0pNb0ojs7yB7Bls7nwazaG5edT9ck/fr
stIwW1o94yGdUUmdn1+wXE6rtOmrAof+sng2pX/JEWzsLjGiZ4yUBUyczfeGamLt
eR9ZS7Zwbj4NRZPk6CU3jKbP6uJwk8+7IpwfcCYwCurVfyaO9/mlWZf0Zxwq8aVA
W+a2ul1IgRQwigj3qy/xNHim2NBQuhZCmOwSnevAkqjKrCdTYHNZNx2ODG1ZnBfm
c7egkp32c6+Zf6E29phn5G/AsEzCdQRkgom5pbhVNK0CSJ6g3BpjOR9+2Jw+eGNu
bUpIEISeo+AhXeTMoLsFh2UCoaY7L1Ba1TiA6NXL1PHRzaP5KL/RPpw1tZxHfHFK
2jgO3VQYnUjKUFmZtUzG8NmCYROl5YBROGIpoXSXcnRwV75etpa5PWobYpkl2qnY
hthkCk+1UTyI4Q0ERUFkJg5kSZAaBbs0kSK01JR71+NNjTXKHCo1T8Cn/QnfcYgn
sO7qzOKrcs9AuR+ElCL+s/2CBS5mT3QXD9mORqMQWjt74OXcusOe91qElgqmwCKY
g1q/e5Tkh0tJ8iR4bMinJxkoH0RLJCmVAa+fFC/3whFyiTvbb6p1xgh61FwqrzT6
7h1UTfRI7YzfL677s86/SLGIB+F9qjKJmzIg7LJHt2zD0HSyQpWYxhTxVlEOTl4y
gofRSZoYNiXszSPf/NomVMfN1EfxyPjM66wZa/YytFkv/jk5eoZRW2h6hO67YbnF
WC0yRkQ9+MbLcfYC+OT56dg0LfUq8RUYtwNDg5ZFf2ribCZop73dTksc5bYKwEZ6
C+JaxQgH1pP43LUowR5QFfgQuBLV7B8fqKikKI3gKcK6MX5lFmte2uC4vAA15uJp
NFjKP+GB+Fe2d5WPO7vA9rvg46pJeQq985I4deFft49JP6RgjZNIh8hj4/pQ79JS
ZdiQ9O6MT5t7ffkWV4taEo7w+8Q76hq7zWLJY5Tx7+ckMlyWPuKI3WdZYAYaWUsr
OMRGgQ+yCsL74N1zX6jNZlDAxvtDXIzLTjjgy7I0kKa9pSUFLBnOkvnj7SzUpm3d
/bLmZ707OvHRRM2OIkTI6xb4K8zv9YU+v8nGZYduGYASLi/36BmqAl5iIZCB/I4p
InNo+aAeOJ+CTUJ4RzYuJA7e996bQtQWvtAibDbeqj/Xy6+LxddUQT3nKWdqLO0s
YZvnRDVocwzDvTB/JrnPRryonV4FuH+7bdXNKUBZWAmnvKFjTvhauKcASa4JqNRc
7s/6ktVY2OJ+kxmDc172KweiG6DluTNC2KfUNj6K4ogMXSM/Pmwnd41RB+FmV/2f
jqNiIMv1YglqniLpKXc3jKImqD3zhRxesa7G7AOTCvGsaVfouxUxSsgJm3CAY37g
NvKxNLERrDmvvrTLCihFidx2hYWBLwDBJH+FiHHjkw5MoXrTC9ZjByN6blN45Z3L
VmjV4DCAwieagXm4628wCgq5eio7TOLs4RGS8DJCBufo8/cogTYadESpjWF+7YmJ
0Tv8c7I/afloQ681x6SAvxamkpU/uobpZl6JdMZSlGWcl2BKTWDgViPOlZbJf7r4
l6N6Hw31LEjaU6/KE5z9Cms6KBq+cRhvUgq6diqQHPJ7HRhDHp7FsoWyvj+r4po2
3FQHKjlGZZ9xfsgtCUy0iV9UV6Q9qpLtGR6AgcGq+warn66KiLDJ0jKLqdmfuhLV
DMUETri6N7v8yeMc3ecfoBvbQb2UTgg9lFpCMiUhf7C3gH8221ZGJ4DLYvtzTibS
xneeGSv2Mon93gOF/o/7S1FafIcUW6y7Izsz18gE4MQxVhnuk9kIxvgUnCZ+0Hli
LFQA1NjE2uE6b1aHB0vyKw3AUpm+7X2Q/StYnsuom+x1kgihmnex+Er8osd69i26
elW+kuYsgknO7WKeQeazFWHC4cSxHQ5WsjQjDD1OKFdrCnemaN4oLGiCIb3Jm8sv
u83tf7viaBbGWeCytzfLVVfmFP/ipzryU2pbTn6noU6qY+PhwwxPYKtyV+aFX92z
fZroiid+7rwBJMz3+HfqUEX8wGbHH2jQg+GT5+lzSt6Xs0n2ZnFQdALdZQ5PBmDP
wRpDBgvHAEosV5zaj3fkX33AJZMCMoRH0qNrJoYcJLkvjqgTOXCr+NKTULPppCHQ
OergNYZ7kNt72Q8FKdHGAEtRlM2mPXK8zX+85+jCx94nBl1i61S/DCojx5fdibiB
czyaUv0nwEaQ9B5ttElHvWi9Cj0+/cnEWW8tuSKQQErp83YrmEL28A81jNx+eFJV
WzFcyzZ/DJ2Fvc5j9ddW4t+Sr/oOdvKgh4GvOxQGKQjrFQPTRq2CKwprPZ218s1G
OKty5vt2YQqlBeh6mGQ682DZ9z+j7a6S5DWr0ksxiHXIBrP4QnXU0M8cArtT3oaa
GUnIXIKFj1uBCi9bvyyOATFCDCxdBRg/A129PYITLpwnlHuv6kjTJxcKn2O1PilC
TOTi7vQq0ZZSDP7o8GiULVPkI03l0ApFKQVOUEqjGrdHl9vRvUp7qbuRxcgv8D/Q
N2THWPr9jvJbiCK5OEiTAs4mUUAiJKzq8odq6VKoyOPi5/2XlVD6oJ1up1oBCUVg
TYVKedNPrL5N7gzUasWqtcPKcn8PK8EujoNxR2IssouTM0ZFLB3hs9mfHIPk6av0
f50j+vXiUu43n0Nd9eQtxTUtjVXfZ+iYPzENhP7UtvDOFzm9UrCDnxhyumJRM1BO
9sT/HaPzJv62sTS8Rz/tLOsWJfxM2Gf3nTk98Yjtw4gjqvWSzefPMhbB6innDaBS
y/jQK5LFhBBz3C47ZdTvArBi/2fvfymEEd1ByHF+MyE17uHiCHX6aHcFtuoGx2Er
CHZIQI8/qL1LpHWXp3b091eArXEe1tTgLGfATqFEc31370G2hwt/HotaBXcqEE6g
m5zewdD8RyeVaLFkjoPdocu0hw6yimzwO31VZkVfOtrUVQa/RFuhYlXil41uogSl
dh3GAANJ5QsTtn6Ul2u53rWfA3fjdu2wLcWa9qFiWtqIvBOq15MdenRvAxDY3Rbq
wJshiPfwN5ZGWnpsunk6tBRSs17jeDgQmUThPfW92mfAx8cpsVwrXfrbQQ6e6Lp9
SKhxECU0gKa7lk2c4/21LEcMQ1rMPfzuCdUmE+yVWWITJZThNPd0jzPDWYje8rrW
Dtoi2aBxOT9Kdd0XOAIzFnG7MOtpsEKZ6SHlMMU1GVswXAPzWv9NhLL2BF6vPkUi
mAUhQ3c+A6l+twtJNThVp13+Yi5SF5fnuK9DkN8fLV5KrFDUOw3DHoQo3TAg/FXt
U8+3Xw7aY25FmJkkP1JHxTfhkXFsRF5F/QHlxPzS6Jg6hjWr4ojIyJ5Hi32CJGhM
YDaFgWEMLCCCZJtqleYc/mSkz6VfIV7zYtQKT/1DS+ZN6/ludJ/ePN06MIG1RMGx
Jw8aeQeG74zqd0+QNUMboO9VLo571oDa+e56K3DsEnz0FSjAQ5xSfr6ubiYGH6Ud
jqmMo922j4UTs1crju/stOHZD8XIAc4kwAFto1uA3MQOrbgAsUXRa3EPiXPop2qm
MReb+fHEWakckVRyeHCnJGbyeVfZgnBsxDsQbYAMWkNrFljvdb/JsDh12qdPhQLs
Oyzz+bDe4x6ipzUoyHgLRXD09H7tPkFb6gjs0W5uBjvQbu1ARv3TUUKSPbqdAVZJ
EpQ5IYckiIy2JcuD090HHWXcJr2L3HteXYOD4c0lY2dVV0eG3+QolyTLDHCEEK1z
tPHmgLUdSFm0enlCdKPZJ8I6m1arepD4pjdSe6VsQtFpTwAAuhq0e5kVXUZuKxpO
08Tn2yJy0tQkxYdvRl8PtdZ7YrobZEhJZZ6CiTJSzZjS0K2TBXxvE/TuK6g0QFXr
YS4QQdkC33nNy2xs53ADFLRlnzhaVUfVxTbtR3iy46y0hExRhIH2MOAwB8LQZ8up
TfEB62fTT5Iq6RdDzif1GKhiwO4CO9f7sQQqcRi9hinydHiZNVQwp0/9VDO+Vu1M
0Ind3iSE0es9xP/g5pHIXasnbWoIUXQrd/UQz2/KTeyWwf7voqymm6N6YXdOogA4
UtHllaM/NaWRf0VyjEDzzenx3gb+Q4UHTZVa908Kpf9/dmAt1EUha8l5hVpm9MrC
d3MzmP5CP/BftNsYJxcozWgFRIpdyJ/Gjd5kn2MeV3QDyA8DlnxobHNueGfcNQ/l
QD3+T6Zn27m/bc6NqaIYk2ej9Oy6g3G7byso8QpMiowXrXv0GKLRRZG9Im5vh8+V
mNjt/gD07qx2yxHobcrcSy5EVjHG4uJTY3jKNdmIU5/h8KIvlnG8hLy140mClv25
NL0FqPX1GeK7VpsKkMHxm64H3bWRscwuzl9g7+G2t46Yp3C9sJR21VhYrFIZPUkv
ixYR9AjF048qy/WXKWFeml5v8ldbNj0aH5Zr3g+hh0WWqt7Z/jEjhe16SO1mOeKH
GU9K//KlrFu/WOhVtj5acvyw0ym4340APGx9qitekAZTQORgh+9m++SgIOa1H8OG
wXqRZIkc8ORAEMJ1W84a4bfuZs4RwSQPG0X2oPJ9LYrtwdGMHjvP4UaSppOh1fPo
TLimp1/qQawKvijs5NSbpQ+W3o/jcLcq8a3yi6a1yGAHK05MJn1t5p3fhubw2ZVw
xXYRT+vwPNiCKd8FrCH59BedKt3z8B87IWlzRgLttUJSDs+RLTlrvPke/Y+hzw0K
LTWSdahoPJTMPLtZPzCmZo9Epnd2KprvaXwqR+drFPaYy7wzNlYSDtGXvSPQh699
wgyoMDzODiCmn7C/qYj/7rKPOww8K79lcoKVobIoi9yRfpt2oQRg0W6LHTs9eyfX
vNeiNGE5jPYBqtyNHKniZfnIfDcOifcenP7kthE97yMqqv97dr5iyuunuThoLSBE
rGTEcGVVoXoRmde4PFhm0Rsq4UEZta8IPz8ArNJ+GFAhF6+NfIQ3gGkVWye0MAEk
Haw6fRIqLXZQLFI0SmposVN0yIrmMkoO6n9HM9FJc2k0Q4BtsdYeoSqdaTRKy/LN
6erJbHPFvBW0J7NFhqcb6x3W5kA0GlapFv+Mr/Hia/DKXZtc+jq0ZTIWhJWPk6qQ
EjngBfK0VfmPBEXtl3JHdXv+DtjkbOlVZthYEZEIaPGwEcqXh8rvF92jNUA4ZF9e
fABubQSNUHPZdzjmalBw7EQ13MH5d8tWWyscfaSmVETaZedjPukIgWLahj5VjwwA
5C8oxCOCgfDq+/MLpVGrEF5P7vioNwqPf2ZJBiu3nUTucaVxc5j9VpS6lEvA3HlQ
lufIaXwfi60tUcNaVqfMBtHNUxe3mnLBfGbpLnXzthq0A7EsCyCDDDjRNayq9vor
JNsDDrlm/iAZhThYtPSkXlz0yjdon53ODBRxnrn+FBuvE6UrNYaKQZ/Wuf79Ed2i
AYflWuX21K/tc9a57h5x0Uk3al0Ixj3wRBD5JvyfooJv7PLwvPVLCAUeT4IT+R99
/gPRc0+KB4xFwhXLlQBfe6Xrohq3rCB5mBN2pbQ8G8y1wtLuALPJOTBOqKR1Mkr5
Cqre8LesmPRnMu82XuU3BI+f1icGDHgxk0h7uybzDp10H4qeobj/s2aMtgxaCmw1
QfQxQLsmHO48yE18Ut/dutud0FVUNf1sMc4jI3ZRs3+smufdfrrSySMpkttOCeG6
qjP9Dqm1idXMT5puJoraMFjqwnYU13Kc6ApthvVlzBO5XRMMbvZmb99Cm7y8PBB1
AteiCXnZT0FeAGOgePN8IAVA/8cTCXqQxTcOVZmjDIqqTr3U9x5sk7afS5kKmyBb
aH9wU+8DPhKySZITqnH3SA9zKSR1jahsNQ1Ne0jMULRF8gmw2O4mVHwqOUqvQOcz
An4UPDNPPFgegxx0w0mjDW3A0EovQOHgwoQIdxYx0MRVN9CBZC/dAkuxiE6I2QSw
4RpzxcLakNdZuqsBhbq2Jnta59Ue9FEH1U3Ee9SMRWYRIRnhfr0IZoLy4MRpWHNj
/Skc5waoqhSHxZ7ge9nqGBqZgVVgFo7zStfoeod2XEP4waOEZLXx/1W7NS62dwDu
gHTlG5ZWqLf4RuEUnqFMv6y6T8JIerAgoDGbIIIP9BGa9VKdUV3vm5yz/aqbH6y8
QU+pyxAQggHaMRdfNGmCyJeYv13IPdcSJ2cZOzpuzJ7hXQbRamIzwYVjjpf/4v7M
3j3UM4fd8qsQVR5X6qN4alZAixar7CxWDmZde6zq/m/AUVTOJQQpJf7bIP0VZ/15
92UjkkKk5amXhASM2gwK6/0et1uY7QxzN5Yd8lCy/eua6wLq8/Ny4My09MC1ylyi
T/8uKWNV3Mvy6ntoIA+IDT4GF1ja3D8f+bMm4x7nr9M7ogBEiQs61TJYDS83sgcF
Q7exQEh1sOYHDC/x1YP5nRN7HnwF5A194Z5Ovhq2hgveIYcwIjLqVSdusx7Crkcj
K6sDNAlHopW5oszD5gFEEJ8R+CJDOE0ZtFV4dajkS44mSaEymSzTfprFmhdg/89L
mIYe9pB0rc9/eutkOvBIim8mX82kX2nt0ZrUTX6+G+cY93NF3Eajui/mtpxgcwcE
wEehaUvhOSo6I9rwKDjzCRuyf6xIH8Lx/oflS20gPX7VefGuisrjIMx98gue/I4n
6G+4eulTPQF8dqp4WASW5w1d8Fd+AX3AD+XQvd2PdOOuBmgm6Hq1Bl1DqYm/T+vc
w2HHJIxcPlo7dKm5Q440b/xg6BInzv70DCJjNE/whknv+PSWHRyEVegLtr5mw2tp
mhssLa3py5TudoNpZJTVjOKGZQnveWF1wZkdZpx3oRhYCmtcIhHllRNsLKDBPJEn
xodN3xUUs7FTnAZEmmRALubdBVJskUwZIKi5xrkzSnc6cx1mnsW70aSSIwIAe70u
OftE/ng25ZjmFbq/5ud3ZISnuW4lMg13lh3H0Vk6P0Z6xNBQu9YwNBr3OsTroiuZ
f0PySvgtohstg/Gy0ZBsAufG/z7uasPzuG5Cri8VfRhBd3zomDk6qoM7z+QpwN8w
6PM54s2tVmU4qW1rkFI49HuDSzu4hYJWSwxnBzk/Ep374+1PhNH/pSOQWDHoZ91G
becUn5El1pJ6lOhVncsYddY+8zle4fTncp99ksaimu3VfToIbsUIGnr3j+eN6pTH
pqNkpiAY3WampXcNjQvgpX842CBkYmC8cT/MMSTS9JZ5Cnc00HWGFsVLPSRvS/8M
9nErJ1CHrdLHgVvcVds4rM7YgN6RED6hK86cpaG5U8PZTuoiy9elsdDFHmPka6kG
sIM4W9Jygu09YnkOOofW0FPK/HRHpwtm8Ls6VraWo5+OKjMHhWzzbJjerzz4AJrF
BqdxmKudWwkCG2+qp9Mby4a21nF5mQHgNiL8L59l5gOYkGmlRI/rXE+Uda7HX6xv
pyFJkPM2axnHhO/7G6NBkEJ3ZYpHYJCEy0fMdRAtszJcFuvsGJqmpJcjWD49yXql
0PmolY7LVsxktw1ggJ+3KZJozKfj7UrZvW0RfaDiJcCub1O1axoN08zdbbOU7BXl
c0KnDRTsd0M/fhIOn4h9E4H6ggSSvGRC4JX4L80LnQBP3ET5+fdsmUfm2JIC0gpg
ossct8IOLMYcyHWEGHFtp1b0icOHFVv79Khbroj9FrfkpvG4Xos4hhkZsu5NVtS5
gEG/qhKAWr/sOidqOxhPtCsEW6E4gZmnds10L0GD1qVPoQxlBk1aH/q0tMxMv0ph
VQ4xEfCoR2z+qOMolQmxDLZ4mBcHxlWlhiO6r0okIiYhxRQdj1Je2jbirpVH5V95
4YpLHWF7rMK91lKyp4ACspiWj7i3j2Tm4z8So0gBv2R+6nw3ZJMVLTtzHDRudQku
nVh6JQJDW8fZgCQbFUg6QKXQwxY+ficZYalxijcs73f4f1aTnqdjVVxxYu4FN2aM
IJf3YLAilK4SL8e674bPI9zgefBvFCoo5ldbRiZhFjSaFMyyxYfZzXrKL2nVMfC4
DQyoGshR8Pmas2C3IKH61ATPUsAoMGiQP9RS81VekqhFTv7PoSXRSpkGRUdNJaeZ
oDu3iTJ3ISBa5oF2k50PEPZdjUdX+r+akK3L6omFBCreFYdrHZHvkWjr5bASr9he
D7N4CF6zPkdL3GdKT8S72q4TTevQlaXvFZc7b0uzacYs/mx9czd5m9egDBoTHUPj
wbght8uF/LhoccnoEj6WVSQ6fgh+O2CHKN/UkpKvZGnBCO83upJgTQtexRC0DS3s
yqWZK/G5ThcrmzUh6ITvJ4uFAhVwPqw6nDIBCDg0sMUtDFRDkVM0FRhJUeeUliki
ZrHifhD0KYo9UjDsu8syxxOlxm4Jmo7xnX+x0JYfRRciPKX3+v6RsLNwcGNf3OTP
imWSkgq4JC3YjToroSb1PTlfJ1acmpwcFE2QGUKHMvwmKzPLFLhuyACffiAndyCD
f2GyEC7lqbP2zv+B9r1ezkFWfZtdS8roDWUQAVsOv8wTSAaRTyAAIizybIXWSq1z
VOhIVNnWImaD1+uetSMZ0n0Xj6RlL/nCn1oebWQiC67eLbtQysMbxMPL1958FAC1
S4n4NjWU7E2h1XA73YKOA7ZG7C0f3Sc3JPVznkf+g8ESkHV4bP7Wqv1J1Uxmiec+
0AQxcdhLcpIWsrpnyWYiTweLV0diU6i+83X41yCitwZan4bJfio1RONxOZlsh3N2
V1V7QZgqQvuY2SbB26DSLpv1FHtz8OhRg5h2/vcMvsDb6Cg0tJHY8//ncMIOqhJb
WmZ2eIAM3FxWeDkjhV2amyQR9iyCAkUYeKbpWuvQ/h0iIcV9m/ohV56j/0wydPES
uAcYgPa2SFjJ6RL17GWBdbx90P0IjySqNBmZoOFLia0Vr/Iz3Hi4X2UDEd3TjbLa
W+KfSemkTvRc5SUt38eCi22yVqn17HWi025nw8BG1+Kn8Rqqu7n5R2qiRyAcgfvU
yx2FJMyZgt38yVCaImmK0R3X67A4rjYx6fn+2N8sZ035g2b9o+bxCvo+Dtyn5667
RVrhhTkDBKZWSNtOO/UZWNmFG2/GnTly3It+J8USDoNxC3Hq8BDKN5IeJZRsRcSV
Y546cd3CvjiXBmERFf5PsRZdH/+B2HnsEgX56ML29TdwNtWWTiC3F4ayrGsiHQCb
koT5AaP/nk7wSO87YKmCsCejFGPjqgJ0zwMjmNs+NbLAgVqwaeb1hk7/zFz6Jioh
kYplSQXE8V9+X0QMbjnevUDpFasKqnUABR/+Nv047Ia0eXaG9XAyGWqLZrpxTTeM
JgDxp1E4f1FIjc57meJhfcDu1luBsqF4m1AZXhWJgR16O7iSQwJV7xmqihTbIWP5
1qfp/j+8e3dWtJi/frI7gZLsKpQ4Cmx+2BdCk1oR/MAcZoIj55yR4F1iLqS5LYZy
1y7A0VAVn/T9mfpmUv7wpNyOdEeaGb3VxdLITc5/qgPfdPtT8NVd+7eWApD5YP/P
s/s/v0d9UWBcl9DHUkyTBVSxR+Jk4/NPgo5d2rGXFIYt31/GdTX3eurEib9eqVDX
jWKNfiNzHAHSYVOOm61s0v+VC73A0Qv/dZEMzIYqSjOYVhog88lJqAkRtCb8bpQ4
1nhyJWtEzhXud/XgrOcm2aHTNXYi/vEkb3qNrDUL6VKoeyuaZVhdRNu9o0ybsBF3
2o1C2HCnCNqUJUlvTWKSnYG4VKdbskajvI/9zcXEVOSNpSDr0AVRAC5gyojp2P4O
MGW9AJHGj/YNN7TuDxi3N06aYcnAnB1dEXbL3J1PYOG2XzSvsxShU66Azgf2FPkh
bGGLsPUpAVhaAUaA3jXV4dha7yDDPaG+Fu4pLZrytUArvtCaFpQIGMCimIf/l4mC
RZmtVFm5NW997c8zQuFFlbqe1oPG8daQGeEQwwkGeSljl0k4EUZohlzIfONqu7dw
3c/vdaXZc9O1mjjd3v6veWBhBFUlzREOHslfJfsFT9Pz1FcVKPsATQeSb/zml8oc
ynmJYV7Hit+o+NZIqZGywILtMHPzLSWP6l2H+eweuWwt8J15uKuyz3tM9P53U5fX
hB1sdoBhaYEhzDV8riW5HFiKAzjCMI8INaQuSrZCVR/7Ek1o8VACm/MppobpReZN
KVkLHc2/BkFwTIKuTQ1PPKOMq21cPCZIlr5rhoZir4vGvqSQdat/Wp47ZeRMAf3M
3A/3m/ojMyqFrQiEPVMfgnM7u6Jnid9JiB2Q2wkJpUh5ST9zj7t54PSVnYdT41yj
JpL+Qy/UD+zeNK45XALOHMGS81z7WN8o5mURnP2zklKAdC1GjwNyfoJyRSxOLmdu
L9GhXdN/iIb4yWpnVHBZ1juB/tpBf8IqMRq6jpAlIgH0U0o9DHrNpCdoq3Q8c6ik
fLcDREWkaQUWm9ooN7WfDQZ4ZejVj0f3GpPjAY75nem+jZX9dYiDhb1VHlGKPDur
fvZgxbdlWrujFw8t8KohdDbo2jGidluxMB1m67OGOYAIha43wXJ3cI9jTiioxaep
j2tM/SvoGoNaMhmGbi0thiJG3xkRTADj+bl8ctuK5c4pHIe0puo7T0R11CbVjmgv
bREdMJXhwsnpikwm11D/w7hXkI3ahoc7tcY3NTHWBFMtX7QrGH3BprtGebZMwyKv
clAhu+lXG25Uji5XStsJ1G2WUMGjCaifrU18FfaNxBSiTCqwcbZ30tDWT8VR2ViW
cA9lp+af+NP9FpIn6e2g+hKjD3rz/ACzLsRFWd2UQxM7C2ok0Asp4yvCULcgYjNe
pvn0QSU3XG/B6a76pLzWqTe0eFNgCmMGczFymHCdQoxaKi7DiCQ3NTzI/E8xV5Ci
c3UpbOBZ5l2vZeYOoF43M26eG6jIC3Rh4adnou1/OBCoynxSBwtNW4IuRH7F33nZ
wXlOqZlGBdKIBcaDI+ezSIYgxyg9EhhNgGm8tDnqdc6EAjKc9bBX3a7mYLWUM0rf
wB/tLPz1nhDP1YMPXWrpzQXISxM1IdVu4BmD2CtmSSEBO2hiMWAgqbVvGf6ylLfW
H5/dKjwsHzj+M2Orm0F47bf5+qyw+QzFyxkbGFfd8qkWCcpBbWw37lO6LxnRFGhA
zrU4v6ZKjwE6CzTfhDrteoB2Y4pZ2Qh9GIAz2ARZv9mh4Eae8RpYxYw773sWzWs5
8DX7qXAjhV/v0W1t/KVQMePNGGHHq/Yztv711oQZpES6AT6ejrmrQTC17qXctKuo
fH/7js02aWC3rQpstgSfDIHjUSz44hFQCZ62h124wmte29IGIna64AdIJeMgGFTw
JEKcAfVwZhXHxK/eyhS0onnDH/2Pcsb3Fx+YafHvLX180ZrQRVlpjaJC4YTcFNjr
9DbgWpMk5uTKTo8+k8sgaz0W89an0Ne03nM/kruwWW6RXa5UO5Q8ZCxnnt31jo40
aNwGh0IdjlZbdHnLSB344K2UbSysEDycJKtF5DCo3wAc+EPSkEWWs+2avqFlmf5Z
m//0l7gszHuCkDlojllePi2KBpEHwnEFAK7JFEon8sIYsG7a/hy7epjy6LUQ2MSB
5YpIpi2/5plcuS/FnQ5gtQfjmopVuPm4GaDIgW6Vpptv/+J9TS2r/cZMT3OHrbdu
y2Su2l9/HRVDMDwtp54hMgo7kR/O1JYO4iGfz18udIn0U1RRP/4yUc0dHGcFdOBI
h+3HYzlSm6UcLoFHA7/c8dwGqHaNfNhjNCR/SuTNXXlLRUEM5cCjMIMwjq87lUml
pFsQdQdYwwmXRP7dwjBXp1lNTAziEw4Z1VWcSEUeSbTXo5bWaErE2XwGbdO3cbJR
gqzfHogJOmWMTqygfmneVq3u+4hQmKh4Br0f2KweehsMwlURqLm7AdmTRJJugRYt
bfJ0UelwQZba/3MvsP0IwPR0JCOKdN8w1+psh5hiVTwQsg8nSBHShEeehmSZH+59
owiUcRNAlj1fCDeWFsDbBRZ6woyjyRzS65Jf/gV2euuvptW0mw1aPHmohrXK7dxa
ma61+rSBGmM3gsVQgTuG2matBRI0rpCvV31uBnkFMHGXy6POhXH8Zs6TxaQs0yUa
86TMSW0IbFUprl1+T6VX1DeFkBaB8tYMG8dHh5sCdcbga2c5zltmwx2lddHq0j5/
SrdNKqgqdFq+PIvflqklBvGbGKwgBJ5Y21R6AlUiyTCfnb5xvl0egEPHBhy1Dof1
B6ybfmq9DhoSEeRgI1FzErphqNna4gQLuMbYWb5D40fc9yeFoQhpRBZz3IJBjyGe
1wdU2LU1XAoav/VYQcO+g05YU/hXTJNgRUerCIxGtf1yun2LMyH3D8maaylDSS1a
vm41zmcb2JmzE7kTSon8iGCpUBiip/5hMv70nwGHqZyS7tBdKV0ej9T/eTn2RWgM
ErIL6ettU0SXXpmskknGXteSpewi3uMj9breS5yf8COe7vb+x+zLNdmjNIt6LuLP
qEhBt3iLGTbHw3pv9D4fCjNxtAgJ+dEjs84VC7EexdYPkB3qwP3Wu1/T25++3iqH
2sGQO5J3tNqCJxYuXe8oYYaYEEGFkyhQd5AzyWFNG8h4D+fgju1kpu47K2q/3oIT
e7UEWkW10yZZRqLddm99U4ihzSY1spweaRdo9cvRW9F8XjOuJNlU737/zpANUo+k
p3TuNwIuRCI3j99/hhhAom2sgbvlyEQKvsCKAag/FNj5BdMKQFZxaU8hmA9UMIjT
7mO/pt4NKVyf1e8blnbVVs2Guk5RGh+RnwwBJWCSfmPtJwXHOiR79oJ8nHxlYRMC
YaVhNwQIPkBcsH6A5XCMg1+NRiCAN7V/0s4wMxKQ8CaWDvL9vi+0Y6W7uyipCegZ
jB4g7djV+qo//zsV2Eel2W7ph25I5Vu/7MTkS4dSUERKXje5CVBgNNeQ22poTPb5
OJo+JztYQ28HBn5YXHctGfd/47cblAFLF6uFfg9VXs5gsapGbf22cn0sAALxLHRS
DRZ3XPr8rmw8mmbrK2Myg7RlpC1oiHUTY+REb29a7ZkpyMEsFRkvdQ7M6btPY+6k
yr2JOcrz7R6fFHloL2eJxaMCf56R1MannMBFARr4BhV9O35lxWe4VM7dsNwmvE90
yxOFY7knE2pslpK2VtlMtm8Ahac2apSuAcsL3c476lgrb4n+eH97Af+auLNuWHmf
jE6//c10m1MGtYZ+jRVagVdcoBgIbs6WmcOqBUNIZNcj3HAp2DG9q7fjEbF4q7pw
8pYRyYlWx+Du5RLbEBalZF+/qNpNhat2F0HP538PCdS9S7lOy5W6aMEi/wTW0Kpy
QvpPDK4Cbg70zVQiCWcxXtFTUaR3X4SXtP4oStgZD6QqT8RoN9CVjsqZ/jQDu5Da
FLoD1rl9HD05QBm2CPVVASBu8zqY33Y8MjmFZSEUhUM3U1miMsLuK1ep3narmYgP
QqQz038WurwAyrQAQ37GoMz1oEEJdyerrbhd3eS6UJcAIhY6fFF5LuzOOf1D03L1
PbCROwbxkVRLcosgy8t0uiwtVD9FGmqWx5aNG5bzmiiIUNi4e/XeVcYxx9YlQcOP
mhEfEya5qVFPfx2QKSrl1vdC1fHcQJPI/OIGTHv2AAzRsbXxvOs18khLz4LQM/iV
CTPVOTqeISQkrfLYy25OXXxCQtFeBuOB0zDNIeZ4Olc9gf459V6Z8YpUshFukRUd
EZVmuW1XnBr0CYbwVwghf1u13WLx/Af0SF59U1+M/Ehf5xO7JHrV4KxMEz0TAwSW
88ehPjGU97ykpZlwlFvtQfRAxhdNqJZAwKLYsOineF0hteRje5B/Mjk2c2x8LvKM
erPK1KCejqQBwkM163lF9w2yeHulYZcRcjuB43kE162mAQXi0v1RbetAmlApjthP
srCa4nvZ1VbPVG62iONV8oxyWML8UtnSd4/uWynBGK4/VU7KKjKFaW29L8jMBsDR
YT0ypxHN8dg1kLO1HdDICu0KCy4Lla8EaRuapP6BkMCUlE3xU4qPkEF3ALShNjcv
tB0pNyfrAVt/3RWmnTMvdz6Dk/mv1aEKfGanojew5FyQDzb7e2EdmgbboDg5cu5h
/1gdSvbdPKNE51FisIcgjf7gnREAY+iarWWcwtaFiP8viohwr51NocZnrBDbKoS5
0iPFm2Q2JMyVdC5mPvUog9ZKNtzTDEKVuk9HErVGsL+w3NjsMzwqbQYHQ5CIBYG3
zB6CkyAlux4WANuMF64zYE7GzfqriDeDTIHi/jxJDrCgsjwOGc/qbxmgakhJmGjT
RY7TaJcKGz4MxbVu4DmK3/PbcyjeB/NthGDib3SIWkG7iEzld8Le4cL4w+iB3L5k
l5PauCVn95KdLn2yG2mwIaBX34jwF9zWsusxIQe69Jj+kh0FjjFrh8u09za/ILkT
uiSyc9zFQBFeJuXHtMuYJKq9hXEFr6X1iFT5X7TO5Vn7bbXYTgAIWVvqkwzJ3jJk
cUAIcwXDv84Q+oARZIk/s8fpVBr0Bbb+AiQbeTzLpxusDDD1tvyUOCCgOTpNdV7c
w93TnPWyMRw04KktvFTqU0QnLXlLhxlGD+FVlvaqNzTpOeMpcfZRdc9NtuUCg6z+
toO7SgjTtUBk+x5xVAt4O4vSDYtsEzpZQ7RX2Zhsp65OZeczzsBwwSPa7TRvt1Bi
UlKGa8m7blNBi30TG79Ks3NYTCVfR3y8pGyWHwUWYAyMQ2XMCBZaaoW0UQG8PAFZ
CbXL+VFTmr7i0P1lRQXJHqNXxC/qFg+hr3I5rQwCvXjxnApaTVNN8HHWy+NpkFen
Hs1YHO/URxcvZ6/B0DhSrawxt2r2BiD46MMXNKRv500x93SFPSPaAFSmESja6FiY
Awz6AczhiYwVOM9SvF4DulReYCN0rQQ7Uovp3bnd6OKIFIJ5dARq7Xy9TmOzD67e
xRrdocZicShIzoGc3ZvZTiZh/3Yh7LWa9jEHwDAMOlKtgXL71Dxm8Rz3oYlOQ4Ye
kaXTzk1Cx0Xj9+WY+R0E12n52slJvCnLwlb0k1AisU/4TthfD1MmFr/xlO5dPeP4
wWa4KY3Dmq6XN6riqMf+Vyuhtgd/ZGxXqfnupbSD73dWbiWywtgqK3j3YJnQPVBo
rPnMEX8TLU2qIyALulzZ5woYXPh4YUvZLbtyNYgkH+oR8ZwcH8BlQsIUYRYon552
nxEzjAepX3q9qdmsNKJtYfgElFsSplcCe0x/Dk7itOHPaExrdtUd1bhcIJnBSbMy
5oSgOOw378nvL4CXrFSoIXLfvlFBPljliOMBmREjOfkn3GWwpBc59IXhtwJcZdBf
nRKiChm5GSIMw0+2ZIeFp3hBhjHuYsHGF3c21WhmxRxNQMB1FkMTmKcFM0RHom3X
6fjSq6t4RScXiAJ6uzXk+KvB2qLNV+FG/7/XydPOyE9u/sKnvWHMkXkocivzNMQw
shrzkmQjbsSvRk4wWNVQHhGx8p/F8tKJGkB9GZ9A854cPvcTajYcaeazGSGg1dKw
bxv1Z+UlQaY1kb+TLryl9tXiMh4Mvg7l9mxTf14kqOrci58OSOtIX8NyDRjLhmmN
PeqMlBuNP4DN2VzR/IqttsmLqyDPIDYjxmvyZ+8tbLhoPHM0Em74LSee8v629eix
br/BQ5V2aJas8+EjfxN6ePyL9sgAuYGNjPkHiDpAK9kSi4uscPBijPnAAjAICne7
bGM7J3eqyLZYG/BVrCrQLob50K19WoOrWzRFoelM94Hlvr52PaqHSBZwgfL8DEiW
NfMgXTjo+ge0Mcr0KtNNYE0ZO2IzUjVy7ebp2XsAYelLKQvuha9wNy8LEYskyIh7
kEe3y6k8Jlz4J0cVKi4uShxtRLCOSeR0t89QsFoiXBL7CTQbW1DxiPUZecDJyQCl
bf1oaj7od1ihQ53hFgKXPqAHEurbQx3Pixpqs3BEFAeBm9XGMMWYaAM0YhlU/ptD
FUtiqWBHB9oO2VD/7d+CbpNPcmQhXjRGDn7V6PI9Jcjv26kBfmUcRhFcRAJ+XSHI
fkYMWCpkbcegORL/gRNVeRUAlj48qKJF6KVJAB4WZYIOotovrij8FsLHUwb+NHbT
xbCW8Ik3ogrwBiKCdtSONPZmqKlr/coSd3UWxqszHXVUuag96NllSwQwr7OsMSKL
Kq+V79GOnAoNFLByMw0VvQwbayOpqG8+rbk4TEZmTSsyXBhb42bX2B6+KazkMjpo
6RO4V9xOMSH34ZZfFmt8+shKpeQGvnsaOyUuL6H4t5XrRU/3FkI/IMZuqdToLvCL
VhNtyMiOPRwKuZtwo0bLXxiGGVb2/ah/JaY7h5U/mRCvR8aFUnROPhmp+ffUy31w
fs0AaoCY9b/v0Hm1272UiZd/FdhbhrKqYTUlBGf1Y7CwKu2qfeknol2hNM0JM5pq
tV9cZKfa2JmbXnlLs1lxdntScWEXgjFj/GgJVO/YOPZ+WkMRIC8ZANPtW1mhn3Rz
h8G37Gh/WOKDlbj9mjfjDImVGQ+pm3gCpt0tphanS2QO2Q1fOKpG9g+2olQjUyMF
htrFwR9n8Hq2u2xccBVzbivprY+ho13/l1dQewgb7vtjs5pIHHCKwXId2rd+E9at
QEY2/Ed/LeXjID+AN3zwOy33s4Er7qUKn9k3bqRw1XilOzFxy86hV/AtW9izhP3g
zokRYBNLpH7pfrumdRAXR6U+rLE0WE27XwGVxb61DbNLCzu/+T1rhT1X+xFSC2J3
+ukhkMbumBpUMHOzPLdDsZZ/1nO7Z20WNYNVxBlV21U=
`pragma protect end_protected
