// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:21:30 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lgCGa29P6a8MvrjARup9oN8Vqf9t9gqOsvC7v7fkXjAf6bfq73c31qsoma5rA5Av
jW5Uygc6jdvEag6Ul8BIQqr66Yh6l8tmHD9r4MUAdPh4XYPgxjXHY7IpotA3CwDm
O3c2R4drt2W9Ap9rZwWSK93uaIRwqbNssyYeclaN7xQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 3456)
UcFYSeyB/hpLv6FAcyeg9go6OYUyv/PaAQUdFjzl1fUpY0H1t8kSXCj+tHksr1pN
eyCE7uAfb6oSgY1y0WaYIirocs/hWDrONc0WBgw6nr1rR1WzGMtZcJmG6jYaqmSm
IIfwF+HD/8dn95UxmWLGmCkSpG7ITVpzXyP2NjW+Qed0wdQco7vkPAAnq4C5DVvO
5NJudGTBUr4YboLWpWOLohX8HNX35oQoWKf1bCRL45upE2Y3a/OBt0pqVFkyQrmw
svxrYL1nAUQu9KXYVKcV4DSS8NjhWDHTDAIFmHD4X9epovzjhSv/tLumVvU3t5ny
LvHopLQCEZ1753kymKC7K3aoHeLJqeOaGyFNgMfWK1yhFUvuZtpK7LfRab7gQe7M
Q07hFV3oee0pnUx8/O8m/fR73Z1Y+OM3+3AksovPqO53Y6Ed6DNHqDkWA189NwXk
0oJEscBQ4mtdbbhL89fL6gvjTEgff5FKXKB4Fuh6k8BSJ4oxx9O/2jRGr/nQR4kl
ea+b850lgsgTg96QDItjX7UNi2gZyX7e60BP02GzGvKz+uo1+ruEJGRxLTBIBzBw
cpadey/1AmC6pt0gqQAm9WIAYv43IV3h8l4zLN6zmS6kRfTljoDcM3Xbha6XnwD5
799O5nTEmMBXQR2cRFX8+uAiA9sFW64Hrrq6JcLW6Cy9PjeZ0rD1SB8v8mRDVq4+
yK2zx/9431jKQqjDKArcn8MlRwkl8eVwsG7TvcahGZR+zi6n2LHjdGQfkKcnAcak
0p0rJqpX/rnTl9q2Z5nLzAriHBaUPoKObPvKW42CMip5ghB0+hrJ+s3ZMJi78ez5
IfYJyGTM00XSVP0Pe9t11fS8Y+koAsoW83jntB8lJzDwOvrL5IBDfCGn4yKwq1i+
8fnzCJcySZp6zKfmAyAvurxgygHeAIxSbBn4Su9BF3p8MPfGzLzvQgBKdJIzJGtK
2+64uRpjWkRnOOC7nrqhcFn6feow3eWwI5e987C59swzx5tfj8JIl4UZHXay1Ion
liM4nJ3LhO+IyfbEEoM2m19i9rwMRNHBOJpTwhQnB9HuDoddPuz8s+pFXqpm/9NC
pxY50CPRif3TjCZDCY/kjmYc6/ofhCS78OA+LN/MeF2T7d/l1TUI5DJ/S/LbI5oB
cqLbuix0poQmtIqfJBc54WIFARSC+1NG6Ns1mRoIsIkwHSbTAjcSfEu4NhZilPdo
weecbZLGsgYcUF2jqSRcx4SBDeJmTDSoNUV7eugl7Nd5S4yx3XWoTOVZIbjkQUGb
IrwEVQTJ9A395PFBg9YXSkn3lw9/hWaRudMPL57cT4tw5Rk1QhRF9vO9msWxb+cQ
C1Lz61xq56FH8M/RKkHj//cCVaJBg3K20yNpNwdYvwoqOGEMDTgX/VsaamuNNmuG
Kh6Ai39ZH7IsRRmqYTyu57tF9ejBOP1giCgZ64B5OPNxTgJAHggGam46r/SxBU4h
uIEj0oEXx9GuQOOjFQ4GGec/ClTTgKIx4XqCwiv1INy8+ZyRVDXN+/ddtzm35hdF
iWHT8AY9R4sCKaTa1MdtF4rPyztiioioVFmdNaOcHXSVjn07+NGM8MwLm2g7Xab3
OCiwL9vIT+682q3CjcTDr+HKzTbn90WEhZvmBtI4+Vqs/d4SBI6ARAQN00D5scOV
5aWm+Ooed2A3/czn4L2kTcXyGFoZBrio7ABtWRD1o8oTLtm6CC6pZAn6ymz1YJh6
bcmGmYoGjevetuvw6hWfYlU8NKtn6UxWkyNqQ3MkPAKnD58LkjxnzTwBb8r9xFmo
KeP1wOCGWszsQvsM49UZMEwiSC7PXt4epQwxUz5HOf308DD5hUPOdSK9F5mEKRD0
pdIn14jrAaGIyS+sFYQtjkBi/n2nnVauPTQKjfNAHz6qQGg+jDbFjjRv9Zp5uLGK
fhiCZDUn69YJPL1GR8d+q8avrkcylmvkp2u2sARxoTDkrxWPk7jdBRESpTCPYqhq
3gYoKeEvbueAwDLg/UqojVIHOE10eNTCpbl94Cwa0HDZx7RuWmuMOS5w8nuishkg
uZ6o9U2K3m8kyA5+as7Rf/v0sJCJ2z0EnrjPCvdYIDZ22HnI0jnmI6X3YguL1mjy
FPin4OQVBb23vzKkQTgWZc5vRXGwSTo8bJa8cK4qi2c8WB1VXQ3WHoZM+5ddHYeD
36484VGHiNVjqn7upw4I0tZ5ax8w8KwlcVqwFaZ/8SNRZcbiIPt9Li24mzvEuI7M
2ut48FuKbEmrxitKIzR2V97VyI3OtJyZK+8zdjzOXpU/qO3h0IJtbih5platcESu
6LJHQUtu8GhO8ecftnhZH1bSaJTGsYSGRJsHRQrW5MySfwrgr8g2SWQqhG4EgWTy
hI4GesuGrc43TkTv9IFWltgKzVT/uyE9j3TJs8b0DwnVgupWKoP5dQZY5aMW2Ow9
xeTGM5Ylh7MxjGRg97L7eKyOTZPidKcF7tWovf4w5GOQ7pPfy36Ax1I7c2gbRZnF
/eM+d36NQrDE+/Tyy0Zm+GNgfSJ9ZEu60tPgBOtEUuZjc1ZOS8uG3xFwAToiGoj5
7z2X1ZM9SqKfZmp+VPF63Pr4HxkjKwd5jNHAV7jtDa53tgfvT1EYKuF/owOACvsA
tOu7I0dWv3kbWH/MNpsbM74AlPXFm68aSfJ9nUrYnweE69uIsJVM4FPPD5JOMcgT
PtCxoCX/iLdnWyJpyEUgawLu4oCCsROYOPV3b66T5d5NJLMGOPBZRm56u8XnRJeN
TFsCDscLZz8g/7HFfoRA/eDAUXcsibOnG+FDAM0mESzsEOrhrYlEVpbx2ReVX5Y6
fmAvClIXMl7q1L81JyFIPs8+dCbKFf+5ucQSd0aKtz3T07CCPXoRP9pc0ZMAN3Pd
p1k556FatYdRi51jQh71/ZHmtIKGuwtTum8qtzcs4wusV4a/gjD+sbJujR2GfQCO
O3yedENGhT4zz9QpnFtfY8YF4ZF/GcPFadWDUzH0gYJDNHS/pic5CpdP/vUcyFY2
9xetyJHCgcwQILtfWRe5VqltRpmrjwRknuJsjAJ5gkU5XuOYkMFR6sUWIOJM4uSg
y30NlGSEQvO2ug9PNmtd80WJZNucRQZzuAck5z06WqrMIFWAC8+DlKS3vD07VLyL
nvBSTYLI8ufv9sI9FNp84HElylPfE1o5c8dWjuNLSkhPvy0x9aRMI9Zp6xJpLpLh
Ozn0TG7xW9fcvkLyUamM1DJYozPn0z0AIYpoxmyWc1beBe/ktTsHCjxLUJQ9mEc2
X9zjgzvemJh1PeFLYJ4GHsVtoanq25WCB4MKbaaCl5zsh/OWSmYvoAJ4SbLE0iYi
+JrNGnwg/WuXWl++Coo/1UdKe7oHE6aAWaNfncq3/aEiF8gYjfMg/O92/3w1s8h/
XvRdIvx4sA4uzYBEZZkos5k/03UJ7Am2Y/x4iHe/WmR9m1WHNNh/W0uT8w1AyRFh
+fw3UYg4gXwSODN/4cl/8ONXV87zMsPwNsa4GwQOQ1aC0AYh+b8berHdGG3SEkTk
BxJA4j/PO3OfaU5q8RZ0JQ79IG89Vh1+pLbpwIhaSFNhvqQkYvkgTD/IbdzYOs4G
GLfyhrF+fOYARW2crG62bUyiDKbjWSNCh0U5LaUo/Y1aAHaMXyenx/kZo19xY1GX
0N5dHuh0aAkoYtqLFz02KmXad5mzIE2ziaX+170PpMK1Wglj4+SnFTA5upTo6psD
cBdhdC+UUmbHK6CAIIir+F1/ppq46NkDqKbl7I5MNN6CdkfGh2DMJcNI723t5WyP
Zb1F+JsK+KkCJZwYoUlZbGhxyj5b73eobkG2hx5opatCIzP9LrUyH7V438T+muX2
JVnPyHrrBe8fLRmKH5idiD9RxvbM7xzfxisLzqVCWZN+pwqXfRXgwWrsxJOsow9a
CMQqpfOEp1h9TsMv6yY4Ow9z4w2/B2MUjGbHt7ItXFKMUerpSA7juPP7seqkja5e
crCX/tiYVYEhCwVTWL5kbwcN0Z17stU+RCOUy/ZwZOi/mOZs/mLgJ81hz9H4FREQ
dJ8/hlkLWGLwlzRWrnJ7bmMSJDosiSzT1lzTIE2NraUOaBPj+1GZm2SFfGPZwi1S
tpukUQfY3rigMuSOdQhcQiHlx0Bu/rIIAdvrhzU3lpNITSf+PicgIgtfs6+4HZvO
reWT43S4kirERPrVh259Mc9i2TcXtE7Iyb4X9zbZ+cR//yg2gJIcoXWtTxxb7SyP
chJik/fiPovKM1gyQBkmmTwcQDKX+ca8S3J3qCHDihRFUdctGZ6FWNjLQvOyp8KE
g6eQgt7Uy/oOD5alvQ6iUoXOSQgeawwj6kYxxeVPWLITePyHmpcgRjq5K6/87oAr
xeshv6BvUvYImf216r5KM7ZitCxwnL0Ocv5Sh/hsUVdKgcM6ag6gcv57qvFZpa7c
+0O0ilVF24sXA6TbN7OX50npCUhjFtF8HUwRwkTx9+axTH719EEtMpMV1ZGOWCeM
bwx/C1z1sQ61IJS2n8/P2piNTfoAYZbS9gpe7SKC92H02CU3Sjzamt9eJKk58DGC
DDntwDKYfSaLVq5tH4zQAYB11ZsPwCpKw16qY0UB+d0YYxXUsJXoDkuiWuYVbfJB
`pragma protect end_protected
