// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
u5YmxHEWC72StA13Ivc85ZXlL43xf05nld1gCiUbGhLxSkifQNazoJhW8NsXCyYBLV3ob9gu6UFN
g6KaPoDP7d3gDdnPzqs6GB/70+TaU2eZQKle2aTeqpP9gWLmb0GD08b55cwHT5N3i6O3SnY5S3wS
lafPEm4NQZeOBaUv2E8eDl8Kj83HKiql6c7s/qLImchpRa5KYzlSnxWvSbms5BpznLueeaa8R2L5
ztRy/ivJty7yw0IAEFbKVaIBjttM60VIOzML9S+XLJXk0W9qfH3LKlbRYaHYRGVpuERW9rWWPUB0
oqwS1Dnx4mrSja1CyYYGy4Qb1E7LbzhSIYNRTw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 37136)
NL96d3ioka4zXv+kaZEVhfHk7c1u91tJFxTIJxZH1Lw07eumn/OneDNIjXZixuMPouxr0e+nlnO7
Z81XTfGsXBDrAt1guodl14vQMEDotx9QrwPZLyP70qnJEOGvRG6ZO6BeMYMd0odEd42KR2kFxCGV
FUE4Si0Z/pJo/yHBYFJ4Orwm2gkwktd5dlDoDsTx/3vi7ydEyJF0xO5yrk23NGwg2TJ/tPLeX+Nk
+mDicAOrgt5OKENrqFWph0HPKKJRebg1MSGqF4gOaGy/0VIQ0IPZtHDY9aOhzqfBM5ss7o3UI9QO
AIt3mbUKjZc5+C7vYbVkiUM2j1nr833uGZtvKiQmdxnAo3+algG7uh/RWxrpz4CJCTiaUKNFjy29
MPfdwxkvXMxvgJlCzX6rTCXDcAbEBGhJBasRhsGv2vzffyt05ACvf0wj4YaGTP118HYSfQiHC3PE
cD43Qow5QWtpt85V+ckEiwgL/BsBLuvwozfZoFZmZjzfuTsyrrooB9L4yDWkisiZqfZo61IZAA+/
lLDDJ96YtR7HuYwo/s9ZoqltImvoUOKjUMSZLsQ3BcxyMghpEEo+nvAPali5/mXW5/wCRvqK2FXU
p6SswPJroGGKX4cN8aoMcf2/VvEVgECMx+zzp7om1TArOgxavBHSUD2HBvDJpYhg7cbHxnHl7mTx
rDBcSVfJfws5xxOurOGxdBfHe1/wk9j0UE0F78UzoRQyXbJYWpeZm8LMQjc5r6v4CDjDu/W3226/
vj+4WZq52QhfHAvSGRgDoDW8Wron4ulf0tozJM/u/IvuLaLYr9csSeWJPdiLd+6GIB14zEf9Ohq+
jRCG4Z2Re+fTNaRJX1IDWzH4IicOCwkk4gLqAzRYEwkFBlsLu+9kWhSFWYmiZG1UobxuaXPqW66g
tHQL8Dkc/uocI5xPjeoU0TTvqWfz6PlLFE1khPPVj7Q9NarS600eqX469YH4BTlkyOMYaoQaL3p7
B3oLpQp/P0Bw/DZvcS01xEUMPH+usPoo7ba50Hzo+JrJPQpBGbw8Akq/4jb/TFjVW9xM0u9VOIHg
hfU2Ox1wavXJBTFc7fhBKSPtOy9CthXpY3nNGMO/Ey+F8cTbgutp+6Ya0cFGZwFeLM9WZC0wsOn9
spopjPJR36lP3JhPkX9hcDyUdP7Cyso2yZGguFG7HuQUE5IYzYuJZS5piSaXJv3XmcyMvGYZjXbY
d9+7IvlObJG6hbkYoBBQErdPaf2ZnjX6d8RfRs0NygqrpT1PYYxkBrFuOfUFq6wHuDsjkl0SmLwI
cG82qt0IUlfnkIJYRtS/dYxnGx3V77xScAxw/TkbU/A3NbaXUVCVzIBRQGV2aK4sosnEVYjCBu69
h3g1uA/JLscXnyD2DVvbJP5q7WFtLDAeMI8BeVMptH5pSilaXIM/mp5c0HfcLhftUveUUmBayCB6
BiaC8gc6NUy10JyTNkS5KFqOA06xfFTdA31Yh6YLDOQqekDqN0KKawfzcOEVJRwZgzkl/hyiA9QN
d7nxPgqBX7Xq3n9o2qnUkSi+kNSu3HAJCThtrjfVS7FbccNuYBws7s8Yjb7Cl8yYrljLnzOvXBIz
tJIaHfz451R58znRX6G5SuJbEooGeEV+XmloPo0Mq0OqfdGFKYpY6pFZmXpGs+vozNB8WA5L4nwO
7yQAfcAIQ1aKIJsZus5/NBpinbAbpTObsQ/Wuw/RXMjT2Cv7+CckXqDmDr6j8RpDcXabQqyfZAG4
7mnIForp7DMRhWR/nSGwmTQEm6A0T7PRZVtTMi03wusdxy90gooILgrgGafIli+n9lU6DX8ezu+I
rufiOQ8FijKbbcT+eBgsaRrUbp3YFikojVm+MytFvd4isrrfusX5Z5yxcxqDTHDYHGNKbPlYptu7
Om6oJRwrqmxleEi2DdbI9AQbgV/o9el3HSxBCk/SEnTWRedoOvSPt0zGLVheWLg6CzRtKTintBF6
gpEN2cHTrfBn7JiRVVbuD7+/pfipUwitfD5mOWF6IXdmTCjYhrvi1jSXJL08/3b/TIsgDsbpYyZQ
cbNHUeXDIgYazdNuDmiycEFCP0CbD4B3L0lAvDdEwIsTZ0L0N67NeyX8GJYGHCiRF/6bEIfyz/7a
Zd+VAkC1r/+tOBRz5sZ1ebzOgSh9cGZD+vEfAVNU8972K+ow/cjF1Fzq5Ctwt6ffleSjMFpYO9er
aw4skAf5brGIpNbWbKKFCErbgV4RNp5BwH7wyajzNHPGK77KKq/Phafv1tTrZ+LvqJpmXlguudbL
D+dVgNPjGHXFU6NjcCFg0e3f5RIDRLGdBUOc5LIaWJ7bMhWC/zFXHU9IDPTXvYmBVzdjKLKjw+Rq
eECoPqxVjoMWRAk8gYuWxLob9e81DHFRdDPlnfOsfCg8adVmV308+CESe+ASAVqaRC/K688e/yO2
65kP8MGKCPFIqEb4Cm5a0ravI/g474Oe4cRH75L8ow2GDxSD3SbXdaAmr1wXXn9gkIVT/RTYiP6Z
8ruF/oYFF7gQLsj4JQwuXcftbQbfecbGpj5kSGI0ADH6xartH6T4j/drTpqjOWmQ44gtthF1frYD
HMq7bf0/hrrcNVkncMAD9UG17TlGviNIZH2w0YbJ9j59t09oXJ0jwPy5vKq9niZPnT8K42JWpWII
Y9k3w2LmdXehPIoNpHMKUmgXS5afydB7S2x7sYmDhJO8Lyjlw71ImmlKf3WvCRkl7W9csaxIPvhz
ojFFLd8Obk+Wfw217d0x8+zSgefDxy7A/qYpeojKjgGQc94ePUzrRJokccFYhMaSSLrPU5ixOEgP
H+gf4rhYvNThozoNVQs+wD02CmiheCo/2mX53mu4mBSqtwdw7P2lncapCCheW0YwzwLj3hGGwcVv
Bw7e+A9ZAUFk/zV2GJGre8nHTzxZsmYnv6BIr0ixEqui8JsigUjB/MpICuoYiqO3vx7Mx829SmVV
N6NEiwVya6LWiHRjim5msXuogKdf0XzshZj80zP5JrYB5+Af3Gg27pJa+eoNGg5hZDm/B69UbDdU
JOd9TElnUtBIfDKguKqfNQSYzQN1xG3V5XLFt4MLpM8EdI2D1HcGPdveu3qeeWvRnPJkb5+AJaQ/
mIcjAd9e1NCn8LeE+c1mTe3mzZ4XCryedgHID+EMh3liioYktgoOty5683epjU8rGiqANgle6MCW
GtgiIZA0JuzuosQX1og9wTfMFPvvNjwFKScMhr/Ek4pIepFvOIIoZ2fX1mGaA+O3LTGQ62KwbE9W
h0BQn7PA2/QOqj+6Jfk/nPxqAmEQyuKRxFafM05raatkAwhm5lSW8SgfxNEZUWxjp4AKDFzXY4CM
TFEQE1Ynjb1iR4eLCDn/3pn1uM+UOOiuw1XM6UxJaMhD7FIW3FRODtPTuccO40CCsg0kJvCkSB55
9e0Od8DOOhW7j5Js91QNKxB42jkBZDN1Bf1y13ZJ1o72A5VrT41hy+F9RYZEl5RFDZsEQMrXeZE7
fwlArQGAUKgiAw6NSdRMXNHqlbnmWbtQGH5UfvIdafBw3QOPums3zclGVuX21blbGxTTi1kXkaOQ
NH9D1nCHxZ/ffkXAWbeVRwlJx9CFYgKomr4AH3I8njTrgHgZNYAXFC9lxVjeauQ/6AYCJa4bDd2H
S8Rt0/LtnH4TxpcGXGcAhPg+dWjqlW7I8oT+jVIDf2+YodMF0P1dW6Z2UNZRsfO07Wy3I5+MPvDM
BadxGK6wrBSn6LBClhgxj76MF3VyRh9Y0dMPwm9OCjLS86nr4ciTMuGFMJGo9/0NZwl/rX0vGim/
fkecf3v8YuB9za6uqgfH48xrrx5AQennZMJ00wU9PeTnlskxHshBDoRj1FEZD8//ftWoXjITm5Jg
S5ynDjj49n1cjgMSKO5YmJY8og95CLxr6UuUQU/RHzmaow6HN/iq5StN7SuKPyaof4BRizyeAqwi
WnjovhkBhrbaBQwMn7+gzcqye1AUFzc4pMg6uUiC0xf1aQP0DvxdfnMx8sxQ86fWnDnBDK1wAMz6
Zjg7zpdFiYnlbFCbXSk8KnCantOjkVaNXBr9LYAHSbBGsF1h/HNynvRulpacsxtc7N7wOM4Sjhqb
L14rwM31SjaU9Xbj8865Ae1jezk+Wmea+X642B4DtlrZ1d1RGRHa8xO6A6BegaUUBf8g9moULEIt
yO0DH7O8PICexXPR9O8dt2F/y7o1+QGOMc6XJfsBXO42FPmeogHbvAjfcS5VmlAePzZChRiQzh1x
tGmvnWEwq6WotJBNnBI4HY/oq7ccU/M9SF3KZM0s+lpRUtov9KfsXxbQs9LYIsNs+Cf8cpAuIRwW
fVsHeCx6L9NqpaX7zqohi0Eo+0AibhN7AgDjNmQPoW67NKnaNuXMW2eUqxzjuo2T0vkpR5JcNbaO
efPipgDTMqys1FVej6LMWrV6iH2qFhWsvV315EUaOTDc3dmZ5kKQLZXZvw5RnD9V8QZQsIB9gJCG
2notXJiWc3bzfqLL4rkqMeSA8HNEP69gplf4c+1vZnhmn1dVg5Z2hvh82td4xNbekmOIZk6wh3wn
QcWZusbZQ5TTqmlumTNdeE+MT/zV9ioPz09+Zau+K/NaRkhk2Gl/Mm4PPdjKHfnVgw1kolLHwPYC
Ua8KFU9IW41eqZvz9GNOA/5AkWIiTrcIY4xOC9NzohSEusDXZOCuJ5oX9H6nJfP+5tcXH7GMXgYg
2/hjc+lTaAPJ4oSRXODmV0cIzyREgLy83rRfdCGKHNj5Tut984r91Tsl4CiXbs2Bv4bI0vcvxGES
rZvkLLHcJRlVfYG/AlQ3KhoppnEM5jwroEzYmpJhzydIJPoTUos8IO9odlcdxJEGCBHLNaBFAnvD
XYOo13rmsCfelP9y4RcJtKvWvDp3zOYOce2PtjZJxo2ly6sJwaW5bSCPgwuSVOrD90nZOldCblGJ
9Tznn3yPCdrllDK2xHHShcQ3nFKcICs/V9mV5jFEVnFUTZqoAHHacc6e1Ag7BgBQ2L3wH/0cOXS1
nrPOL9SDbAEwZ4D4hH54vYTe0Lp38tI8nZ5oJWXJDV7oRBJJpB4hGflpDEMS/uGwLdfy4AleBAtR
o7m5yVunEsL16sQhQMHE+FUASYXJA8IlyeCIRyBegrDoPR85C9rqOk4EnX3Y/oJQdk7L4wWZ2zA0
VKLGsFKcCXVHn+XgraeI+bVFn8Fx//oZh52OWwQqpDbmCPshWmVLOCuOqSjlj7o0NcG5UpjfZAZz
pkRRbi5JUsFvRGV3bFpbq6wpXn1xCqCYBz37vsgH3FWNcI1fBPvd4iCb+zu/QCuIkd+px5Y1SJfA
dxTgwpUGf9muCnSinGMgsUzJJgf75h0qgwjfASzuicow5OkrztBWi6/k+6KFYxjszAWf8RuVSsdZ
5Qnpnv8ysHNTz4yriSDsF0nXyJaos/gSSdpaae7xwT/DJi/tpKf9dRUXMTgqT5ftkhkADoabKvfH
gmS5ee50KFo0BtTCdOghh+FntxYqkCzsZO/pfYQw9OttcYSzf2Np2jdLbskkwHeCIgOaQ120Pn+g
NSinM6J9pqktUbY28M5nO9DXBRXFfEcsumnn+QbvMMngzKO5Qw2cFT52NwAcS32G4ObCElmQWIvq
Suv0Xm/ojdV5ZsVdx4XYobmKvLKsoRFzAHCtfxnLPokD3DlxwUDzID3zVOqT3CkA+qJHSa/BfwKk
uhypoyHoECJxbqF7e1RcVF5sRy7cK+NngLcoeybdNsM0bJU3/uOfXxnK53DekZG2pFusSwyXahij
uc8jbVXVmFxffFYfk2+y/2/rDKEga7w5CWgyPE0q06NMOvmOBWdnQzxj16sTP6CE/Tb6ic0jTke4
LTwL5/OQhXkUqkRycMRRzzJBxysmpOaPqX+4itI3DAqrxzmfWwugCa7qeGaEjtZ/8oj7Gny57KSu
soUS7dRE/4Dr5iWCP6zuZObQ8LORZMhXWVCU44Z0dlc8Bilfk4TQ5Rp7slnYTqZWVxv15sIIC1Bc
tyx8IrKLffASojZAyMznHaxF6N3wGlk0ZtS+9XZHTAsTN+ed0zrcde/s4T/Hkc4PMPR37Q0vg3Rr
3MVN4xiuP75Ciq5PtyYe9nSkUize9FjEu6KSMHEBvxKxDbIgdw/LkUH0HGFyRdUvm1TEIX3fRyDM
wYKsLi2zTHOdO2nPomrWyhmtrLOpSxJR9Y+6OUTzjEEcnJX5D8wqQLNw4/hm1k2ETWexAst+/LTi
fVfIxetg8+pugtfOig6FJtQHtcmX8qU0ZGagEiVxsjplQO9JVE69ag3H4FmlBe7Mv4BcB61LyVcu
47lpPhqNIu2e8ZsiW69cel5BhRg0v5fSWofkK0BFA3Y//vF3yFd42XiMcR2kIIekQj7M8m0Ywh6j
kqj4Sh3wBxB/HYXb5DcU7X9mKZ5pEkpNlM+IFJ9n3XbOdeEMk8dtfxitjrpxMfgqG5ViuZ4Iokmf
0sqTa+tvLJNJ4Br/k7exnpj4jq1P3x/okOoeaKr0BWgPWMmztknM/YAX+n58bn+XmKxxbYu4LuaI
7h5pPqiOFeBKkSaCGvuZMfb4OOldhK0GOrjjaCn/I9zAPTtsZZT375RMju6Y9ZIt65JEkVXXXWu0
HNMIeeR5GQCt88JpF32tM16DkiYT3FaCelr9u9YcZvtv7uZQNAQSsDL4edcq2rLqMhu7hsJri6TK
JRs4fZaSHVDYFpG7eH98JNmK3RDUZm+1PkLH8luKZ+QZ/sazqKimPkvaTAjRpVR+imhRoMzyW5pV
I5ZysleDlUw90B/Ssf6BbZmvNc6eArWrdFp/IWO+CBuwu1O6iJk6hAyvpgICH2guu3eXqTPLglG5
N/OsJd1nRxXg8GZAJP541eqTn2fesiIpnEXXQP7z+Bo1RkWKptpuVA52AecXo6Qx7KKcr1Ctc7+a
aU7BURLpapWCJbnDJnjPw7KCCZMppCwpH69bjJT4ZssvDon0CEiFMb2E/ciW2q54w78X1N4WqEmq
2cJdai5QvBM6D58BZXAv4NIZ49ciJMXwQnn7xiT1EA6nsVjpGJaxKS2fTuqDB4qXYtFEG+BaO1Bb
KlzhqwjMlxN7pmRPKFtcnza3Su5V/I5kNm/SXXdBo3tiQRL/wzLUldw5SPFgnp62RCpG7DAwm8zq
vQWXSBrOxP+JiIiavAmnnvp3OV8lpPSjD3V1G09EVm7kXDSXaFijErE435gBY+jkSjuHf9ovbfbN
iHhPS9mBW+LXsNn9hoEueMBW7pC8pUGwKnclaN12OUeT5cl7ZDi3/vBnoEbUf5EPxRvlKEqX8MMM
W/jVGKc/R8RPryV4bVLQMQhLhR3RISpU70fFvAmXZvvvBiDBlID8sbeOueqG+6LNxrhPHZr2E8GN
z3bKzGjhJH+aUm9RjAhjjv5VARk0/Dsjy+WOwWuGPRthu/0GbUYr28tl7gDhEJMK58wf8fMlPWUu
PmxpDe5YUiY7gVozMX/BRwe7r1jCGfEa6pJwjbg1QtzhOH3n4oAsXQbQKEmtmROkoKUQ4KT7QNme
O7gmeOXycOU14hHuHHhP7Iww4hh2tPciJnMLZVoIRfWCV5PzoqVlHCilTzX50uOgLarq7i1BZIjp
qFmPsrYAsVZiDKPMxMTc681+9go8qS/d+Mbzhnj0Vhflt9bZy8O6f+5fPq8AmVqe4cYE6P/lf46j
dxF/xNZNgQgMGEWrc/Wl1Zdh4EFW5ydpP3iaqUvUOhLF9Ob4ibZ51KNYwW6hj/yAlWo1sf0BGK8W
5PEjU8xBpxjk7revIGudLEzqBoOfB7AAoSkKRTqrk7da558navktVfZcSrHclKe2PtYI6jaseC8n
a78FB7wAxFsIqONnEwoH0s7sSkrvwbXU9Lcq5XsCnuav+4rhHuB2EaE7Pte74FQf9RvgJvuXj/GS
4uvoZXgMtN31RsSL/ziY/Og1QhU4nFH2C5zp/1UHzIb/4uxZwkjo67gGB2fWxiO8btzi0My9jTAm
Qnhr1YOwElVnkv3NIJIEeo7VTNdCTqvexU5oy+2JPVBFZpQDdUrQr3rrhLfyYqJTgFd8/HzKikhK
0mqe6pvPfv66wChcOHjD7KeDGuccG23mi1bybF/jz0F3cM5Z3y8bEYMU8W4Yn9G65r2Czk0Z5K6i
1y0eeUFBLRAHHto4l+rkhgVeiI8aoVQD6o+76YU5znU2HvYkufpIksebiYky9ToKiBgsQQvEJLSi
cTCucSq3OrgmQ651z1RarPGUt2JgXR9apOTULHeWyP3kSngDB1aL0sQDZULZroKR7+/VT7ZFnE1l
kHvwPbxj4FRxCcHYlxR0RS2TQNBzFt8HTVORtVnFgK7Igy2Chdv4y+8KvxUlGjV+9FgMU/GzgxKi
7XPKhxW5kovBn8pDQ1ljpMKcGkGO4Y4T21FVPSGLCpfyq8ybwS+03DsFuuyKfutLyQevhCa4xREW
hmsC+h6d2sVGf9LwbnkWvcD4c+gF0+uXTBh9mkt8coB/WXgJ6m4gN1o3oXmNAiC7ADliwZQ8MCct
MW1/BhKUPhBFv4aTBeGVIpjN2sI38advGREhyONBYy0m23C61iup2zQolcku1BbEBbeTn3Qqqs/p
cvCzFJ2vcRf10zpka2dUgXSXxYOri3Fve3Ce4sr99Vau0low6eAWhtD6qW62xt8ZC+ZJz8loGowv
vOj/+OccO0imx0JSYbmc72bBU2MCOrkSLnwWZsN59j/pAeSVVYv+G4Tc+EatqKggKMPO26TVyH0U
sixd2lU2OgxgxIgpBookg4SE8xaVIISjkkq/bDfUrXa2W7N/uY6kFg0DuueREfxql6YPFU9gN2+k
wWdiuAB6TXl8sk7Rj+OxGgj85HzjAdFzU7/mbKoYm2gp+a+q0ctAtb/VxCSMsG/Z3RU/S6RKUmjD
p0WfEmVpM3YOOuR2jl7sp2B+PtRPHnLewx7ebGey7h+k+coIT8O8NlW4G2vgLamBcymoqQacZSLc
JGobs5E10Hb79/VdGL6Ou5y4+sE3VG8Op/NKNaywvBrZiJYFkug8TrwZ4NO/tlQKKGlNF0zAMtj9
CSrYVwtB4z77jzfPzZ1GPAtPCpJNNSJxLzCJ/kE6alL4JrD8k/66WLDa/Cl5gqPQ03CCh1xdQr/o
Hz05xe0MSv98ncZbBGweuDCNlRKiOKl3jgxBHxxfJKsZ3fiVS3oBtYFYEAtNAKr7ExvCOZQ9YsLo
FBFtqr9ZEPfhkJ+YwGvS0sFfnpdkFiTU1zEWbB4AkzSuM/8CRYAJG2c3TDWGBHz1GfauFI06c2xL
S0Fb+WTK51chyK7SiDiFih2Pwomub6PEIc6ZGaS8z/7VM1G+4ks3j4ir/39lBVBVhzugUY9/Yf91
6c3YNFfu3nQgtMYSU30WvjDDe0NRUqTmI9iYijONHeaQkWu3RGzP/XmPfOQFZuYEhPlUUAylx+h/
2x9+ZVgvFnaNzD5b0L51qgXGfenqrOXc8aylC+csl0h+LEt7IspSvG5JY9+MeERiLM2l4+LHQqvu
/u5B6DnvHXWz+xUj8458g/3pdI3UGux18MuKqC18+LlNQyC23G9cjgVjOP9IoOALLT2fVYPDlAvA
WA/IDE2reGzHaJg8dFEI/BjmWfRqmLArFV/TTFJKfE3XrOy+273qhJjrQBK73IDYwCN+LpoxKu70
BUybunMijJLuBHuF5gdnJ5b2HJqqcMBpmY2rVzPMURdWUwHOTUsMX+oiMOFpoAYRQfmkZf2063zN
Cxik96eTbZCBKhFuadag4ZKgKfFZshhUqgHMSGVg3bDKHtOftg2DZ1Gapq4seEK2MOVlgd/NJFjA
XfsfyYk17Z6U+SwALxEawRROElyLClY3AInAyz+QQQ9N49a/o3fJpdXTFLyFm2udgnMILDjfdQlr
1VH15sRSj3WG8mSrNILzPz0Y3aclRhzKIAagyEhX3dcRbDM4/5T1QUM+Tl6JKsnUW9vqJr4IDIgA
3zIC8GFn6KKwrPlQOow7KqT//tU1O11vj9x9yDFlFtwUWvrzE4XJXB2TdGcH5my3spVWyI1y1JLo
W0b0fKikfk5WMajS9UeEONke5QggjlMyMlfQBtl8A+808CzBNg1Y2eKM0sSgJVXNsVG/BzAt5AfP
4tEwtXQnLDsi5tO4TkkKcmFF2D3IwBKgFAjcZelk4Sdnj0XMdd9eXOM03xSkJShV3cJY1KDU66NW
XfN7M3tNv5BhXSGNVpoV9CrHQ9fJx48uotds5I9P2O3V5nqlFHNq0GIYWnTFX3dMGbHI5+1xBwa5
6kvArKbMxB+iF1gDC5IpHaCb9WCnQx0OxfHXE096jrmfclQK9i0vS52li1TKAnkNzO2oS8GZITkm
iSh/qJ1NJTSdZsH6xSX1gswt6L3aokkz7JTP02JuwFZ5NX/Vi6fF0ECUE8EO6CXo3b+ACf47ZF8p
FxiLVGXg1ZnmGZA/ViSMgLnxGYSzwNUM3rk3XeJGkeUbPG1BHi96W7Z0FAIjierJ2uLZU5g0JGsr
1mn0vihpsz4CqFLYZ+Ip0uN9s86NpNY6szm5hZwuiukyGhaaYF+i5TJRZeVCQcTgWZhIIm0wJQZg
vQdwtEg6VsmAaGxNosTrbaBCATzRSqbsErc1IoQP7/lDhNxlZCVC1T92w3YzjRxCB3IdpvPc1E5R
1S2JprS29x5TBjdcOZxLCR9QlstK/7OfthjeDIbpAEUBeCT3oXFeTdz4s7/hm84sXL382bzdws2i
32NRNXPZbtY0MRvvKAv+cld64gxVdM+7rGp7dQwuJR1qnlqZqc8E25s0mgjdLYzVawJPx9PArtf9
9INPkccZmtnQYMaMDvkBuL94pNY54O9Z60cMLkl/umqdXRzs1TtvsDyzK7Kgalg5e5WfwZVaRlNW
Zw93R80YWvLq6sNICOyboP6/jYnlOWU99iRv77SMI/syBJ01uBveIxvRjZZbyUlkzA+A3maw24JH
YKiUBLuIk6Y57X3m3Yx36hKwoSi6F0NlY4qOxgVrEsPaRyrQU5qGU/cYqPqKdcgFwBk+Bov2pNVU
lgltli56nH/Z4HNjD9NPyFT4+s3MMQQqLYEkaF1+Bj3YKpuHJmV289KSM+HQBZdhKQh99+deuYB5
BJhZQXgyZSlCbttL9d/Ak5uG02O1xI/gSIMklfttxEGYXcQzY+jWguUks8uzS8GnvtQvqIH7T2G+
yyegwxYCxBuJ//4wioN79mLHp4AY3MFLkZ0XdFVfOMjLcm2Q7Y6eZZ4E4LTPaK/ic+lMbcvnyJWV
Tw/6yT+4scCBZr79LEeZK3PmKLam2GNG8AF5VoehCdsKwJMPN6ZFp7GK1SAPdKek/XpfrH7l2tPr
LEelxIQmQRdMz47dVQU5rNyXQWjX2FB5uQiY2p1MnXHddSMlf4S0IcL0RAnYylRSpDya+JENSPgJ
mlAnwX5us5DgHC8CMg/BrCl7g6ommwFy+DB3eTjHo+T17BapFf21v0gC0U/O6LGjW3g0xKCHyibo
KpcdtjWfx4QiSlcpTO+Frdq/Nrjlaup6GBsZBEpnGWV3wymk/+++6WYENyWiXvSdEdUG8yXWJaDs
JkhHYoP5KPe/ZCpnweVqmgQiagAzQrcHl2kyNSmyfoo2F607CmnnBFenk5xbJbptIRWVSREuXQAA
ENBFxu4MQhmQMgLQiRotRGxU5ayspHNr8bv1X8+53+GmijzNY4hCnoRwJCRsEszFry9no/fawv5X
kViTTty5ih7c2fTOVwkLZHERRg3Y0rjvS3pd26p47mOZ6SraU0TVT5/8kHHoIEXKdZkC0uGHStlC
lJUjF4D7ltytxtdRznk3rH6Ez+R9/tjXfU52akK8Ld6iybJ0B3mMwbqpVzxg89QXd+6uNwL+LJWI
jKY/Y5F/yW7ORhpm8Ve+tb1uVZbqCnF4iTQBwQGliaHjPqukJzsGGns1i0zkCrIHI35abYSGiMRJ
CKECOei9fQVvo2lH/MKUTbT2kki22/RXDuN1UxOcF0OZ+eAKjO0eXPyIfLcmx0BxsCnjSx49ONW3
ksf9/eF1prPzDq0uufM4Y0HDtQXuhzY4NzSTUpywxF+9bNkavamG6DofAzNtST0y/4sW+DDxNIpY
X39UkGHlBptA7FBwWFCH8lFKa9NGn8AyjRtpUuysH2tFEnuDNvnGgG1eN0rfmnr7v2qUa+K5IDYf
J7cD3N4SyfBdw4LIJQ0pW1/gdNZ+kCQg4wagiMdK8kk4n/d+TVQYE774p96rd3NkAk96G9t2ohZL
6hmgdxHGNxIpxVZZO+8qWWMwYlCVMSfvwc2WFqH1K7WfNa5qZTrKdz5F5rf+gmauL9zqRfsmO0Xr
bLJGxlrm8cIch6bj2CEsbEAbDBFf5nP8cyld3udXnl5h7hJPJ8ObIMoxquPW92TTmxDiS5whiTCN
fIpepBhbyRn5vHOjbzlLA/lvBtteDBXmHF5dFjRdL0QP0hwlPZ8ue6zpTCpQTgvxkhkBRE0qv25S
PfQ49oqZzkY4TV6n8xTxI0UlZaXNubuRt9+pwPjZ4TgaSQuQAo+MuhL2nygxNP8GdyFUXAxD7T5G
RyNagCdaCUoRXdVKQaarQGCppeKUQ2iKK2tLWCFIQLqIsxbRWY9Z19+khqrAMeny9rAEfjyhFuK3
pKXl4lLmKkMi9eKQKU+XDYQN+drdtCFbO2wn1YL4VYcaqaD3stg0lEFDKLhj8w968ttRuxmNCRpM
0CohuojK//H7oHaPwvLMDVc+HDw3RonAAYdj6cJtH03rLp3hd+CHNXqemJeOWusyYeQ8xSnzMGob
ugcTYwdBMIZLeflRwnZkDCyVhml7roKR+0Neboy7aeFr+c74hFMTpb9PtmCCLkwrP9/JhPX1XAE6
wQdF3eJU0l4xcS5CKWOHzTBDC69/ByXcE/7kAsBUT/+q/BEEarPqqgXu16xEk62rqiR2XWYDpxnW
7mDcj8Q2xKd/rETw/C+Jwa4mk5/sdA4AkJClHCQQdch9iGqAHi6Psi1aF4K6yv+Dgtr9OsJ4s+WC
+Kg5DOJ+l3LJ0pp3Rz+2khBcPwoghor97kUULcet2GLktsqY7GJDUTBJc2rniuAyxo2bLn/TaViY
+oflKwqt9h1ZWWt82hmG19kKJdbQlOFXBXw2C3/orewWQbpX5+EhpeAIRwRq3iZsdh7N52SX4KAh
HWKieCQZ59o+FcKf8A9y1fcGchg7INQP8qsRh3/QzO9xbLuTZH2TG6mh7bkL46lkiwqK6wVtQrQc
QKi5GqOjSNBYWvXjCC28rqCxqQ0VtVB8lJbFytG+9uvxnclXzSyFvdxgM7Qc24fdl7nDjAGY3EPL
atmbks+bm0xDlqQzdi3tO7FwVe8L58fzv6MTbmJFmVVCwtM+eYL86y30ZjAs08DQrXbDDxKVhi4c
xglsHdnHYnExc2BPQ5+lYLwfSD52Zh9uFAWxAlQzhh1h9bdAthZSRTLPwlHIXcBBZS1pQ8M4n+KR
gb5bK5DNHoTGXlNC2SxqCxhVN51SKyU3fkwX02JC94pHQXZR4ImQKrcCi3jD9Lfhv4cYAE+/txS2
Q+pXtTzOdPqpsjvpKtrtchWbIVOFSxrFQHY0BRP3O0FrvDDWIJQoGd5vA1eA/Kvuo2IKZc4sVPT2
0jbdaSg5zEBKFVLkrdBB0JEeWGu//i5m1FvI2QeRLEbBQuaeR4vJM+kIjQcBxbgaKbP3sBbo2hF2
I+Nn9KI37AlTt08F9zqUDA5fQ4H1reeebaFOTupL0IOhLQkvBYvtjptjjsw7R/ULXyn+TX4QSME8
LV0BaXk+DSJIRBhRjt9MAgw5BEzTW6BR5P7tZifbCZPR8DmcPB3r3V8/dG3XGpIGgMKlNP4k8Gsr
6WfsKnINAkmTd32pxtSyEYfMok5IhENEpKbHj1eMzts7kA1A6RYjPc5k2pnTaG/lX65RtwT6X23+
2o6gmpc0K56D8IQe9eH5KllDi6eRJ9B60tZdPUHbtwwsV3o4evjq9hNr/ZdYfFlKEctVHZBaiYGr
V58DX8tjlNeayf4NC4nLR+KRHiI7k9l0X50BVzolqlmDWh4Xmfyb3Aa3R3sctTxsQ/gE/92k1uW9
8J3fXaSg7YcvGisaZ1pMH0NPqGZJqUNQkMAG7dv55kVHoFZXTm/HvRvjuAwXG78tKoX7zD8mcCJ+
8e4nPd89pt7UR3MLD1ErBycOoHnvlvnHFyd42pZ6YP/L0kv1ha83zRWJU71rcRN4tZSHfVJhuUA5
X+0MFUdJ/6cprTwuMehWgxKOxqzKQihBWSW/n1TYEbFZt+UzzGmJDkP5SwwUmIRR2DAqxnknCg+t
6iZse/CGASyWYEZtxFr3axJjrPzsDcN9g7SfQpREESaV1A1xroHMP4cvbJXfsB18As5sEDEZCgkN
bREgwI3Vlx/26MbxcP1K2AEOtKNGr5jSxtnd6VLt1hIl0AwIR8Heg+w7CNDWmBS9oPVeNlXy7LkN
oJl9cHAk3Rh99wrCkk2hXj1z/zyIyE1ZaRAhsKMhAF/oJjjaZE5Te+9ZVSBjIyC+elfp9m4l1nhJ
wpfdW9IIMd1AAqSfOs+/x+Nl89rje2TJBtQdKYkode+QhODtA3YDCyvY9vj0yctXz5aSutmeMzL1
w9QOYRUEhEjQro3pvUb7i+RufVGPfUwOfedUCVf1mS2RDTj9/k7GgE8nJemPgJMy69yOvumW0pcU
HXVqVfOOJ1vDS6ZWYHybjmv/QgntIMd71nWHQsZNd5I+DOLwjfgqycVV3dos88DCQOgn3hhO6vNK
5ll7/HHhtQ2sdDo7c3btYIgq+A/8Dc7YiadkYHSGfqLd65nuRmgAsLfRlxsxonxiJkAXxVfpYL0U
hD817sclAmN50e++3AQaiOu08NUIcQl2WQ18bAqTlDzi7EkCoAHdVUXFNFB90+zl2FmEk2FR3F6t
/p1jd3SXI4Y41WAl8xTgyuE3tyygAGlMuIIUXuKGdFBU0gNz/pKD22FJxIJ01vd0FuG4GBXwebP5
11u2NGQPsqmCcDeSh15jUGxHt3kYCxLRVQkuY3iM2dzB8WNLvrDiOwTzIq2/rNZkijFfYwzXDZiF
Nh2i2x0RmGTmgVpqkltTPzd8uXaRtYA0aAhxHdlNBt/f11CNTdwTvdZLwVFXSd0AH/fZWFS40MPv
8uZVBZ+3OEFV0ii7wAeGjONTKZPnk/JKGLdM0B/lBFSeSis8lu1YsWpEGrD6F/9ElsqqBLZ0bYi+
6OecXZIN3lmOCceu+BZ/+0BgaWb4ue69CXKNcPhQ2QkGayk8vrUyS2/j1ApyJRfsSmcTW85M1Ajp
eYvuInGoeRCqX3/xdaBvqI9OHRZ0kPipXuVDiRprZzQVpv7Unl4V7XZOxo1/sha5E9AuH2MX5Xeh
Az4fvM4gI8B4mb33FKY3AnP/cgaGKpbEn+kZCLszKO5bw4Ekm7/lW3Kzi7l2sZ6gJwfp/9iejNxR
nZoF6pbAwH8HrpZbY4QrmHr/Tdd9oomGs5RAtL0LArJqa3L/OqTUZwZqzZX+DW3S52B/SWEZnDJO
Mdob9mQ/lw9XzkdekaBSRmAHVV742X/U3e7qiBO0osflJi8TDt8JL3H6UWmnBPxGnMNhEY9JV4zw
gx+7T+O4zmoTpuI1Oe6dkTkf5CB1/lDC/3hDEoyCDe4BQ9dOYLrPvVj9fgOupARJSMMKGp0o9dYZ
w1lnCipGr5+R+kMhPaaJkowIqbUPNy2k+cu0Tj6ts43vSMANYZNgR2YOSM53XWsLZA45p0LHpogP
FoGusF5KZjfha/j1Nj+cZomJVyhTbVsSCAF2A9c+GSdOH/WLr/RfVZdkUEVVobQiOMDIkrf7uQOI
zkqRlMGpEZ32OgoeaQ8U3dZyZ8XWuMRyIA0WgHs2JFX99+FQUw4bHuztDr0SCjdfuL9em/zgX66S
JTXuMDUpLDImOsV1XzSxHWSxsswYgADMLcLYwFk2+XPojX1SUF3S3OvdwNLFXUctY6tB3kMMpuUy
vHcaangsQpknb+4kh0wDSE2UzIjEXdGa8GtP0fn5Wym+0SgA42eXNDzk1H962FuKly8RIBFAdDLn
AveAXsDRcCJ8t85GI52Pj7q168EEHeqPua1gWEgpTx/7mgZKIQDGbC9aG2KOAIsqlgapSBQy0fp2
EbOd0OEp1G1sip9OyeMJkiYYBOvqtCu6Bd00E6SQu+ZNpqEq80rV6lRxkUQWp1tPFdRjWaam6Vii
44WtR+pJMTHZLwCecvhit63lF79Nb6lnBR1JMn30RiQ6CaRu3LtmLQAtO7s/cKXJt1NtDOPbRN6A
yLUgeHYFsyfNVbsYhgIkHlS4qWs0c4J7ckajjx3XhXrgI8tVCVwaKKsUW7rIlbpibzXKAeZrq5Vg
uqtnGsVpbts/gh2YeCDLy1hcv2cgSxYh7scsMEx1lrXAmPIZyhFzjsmgBXYOgObU9T9yq4OKMiww
nTTEymlH2DXzmM/j6RB/5IjomyE74/L2i+DS5Zb5f6WUNvtilU1Tdg+mBa+M7VZh6wAO7F784zSf
TnZc7o7fI8X443DhEybgf9AJ424qbRuEsZiudZKR9M4fGy2Pa1fjdeqZSzAW5ZdhPht8RI2zUdGk
YGFzBTgFpByzBA2f+XcieG+wrswOhIHsCBmAItM6Bisaww2CBsIkQy+OXtEV6ASYOSq68JK8i+dZ
eX//01fZRsMDPhpm+MWPHTuU3gZ9V1P2tHK2++M1oVRmQZ27B+gHNw+jNL5QeKkehrBHV5hHefhH
+2h2qolIdUf+r+xzwmbOROnse1nqvGCgjkpCfLLUiv6xis36+QOKPmNvDy1XBPGKDDjKg2iJXXbr
zzqeCxjDvrMgm9y2P24uh18upi6EiLAEKmMBALEO7cWM73yfbMRFn/gRitpGZ5NCwN+0L8qpmuZS
uY0K6BwWtfIcZkVXrrMHHL3rV0zw+fzVEXXdCmdCUhA1Z3APj7aLkwpgKA3L5liDFpEB0+0knBpd
+1TgBF7bf6ar3Rmi2fwBFxQojVI3UvNJ/1rACLmtFtWvKGgmTfgbFOKoEfjziR6+bArTBH6XDCXm
aM6wlImo7dhCbcZ7X1TU5GWxxAc7CxGV2UYUqz6EgiuR2VPcUTTTbdMp/8soBvahpMZbXHAFee/i
Cbhbq9f7/XBx49A6KH1hPAppTNkODXbBwJBj8HnUigRr5mc1gamZse3H4Ot8jYM7veaKZs/CVw+Y
ABmIhTiR582aWvpfrG8eLKQw8v3NzIZPNyjWmIq/WQUjm7Fy/URKBvRbML/COxqrg0NY2Et66La5
etxVN3gK65cNECPapqx/sYc1wh1AQWjSARg3V1ouQbJEWt0aGorMeiFj3NGTH+GXGXfw3Kag9LiT
mQKKsGkyP94Yosgw8PPht6kbp8uymIAtmsjhy+Cr5+gYbhLZisYlFFVTtnRlnItS8TCFV8Y8is+h
RMubjDHb+aoRZJf95h86I/hDVcfxDsNQDf70iYWGTSvJvFz88rFV8wp0el1q3VrxMCrLNvCWKXSF
qOTeEztaRv3ImR3izkFPx5RmvlRnGzDQQnb1FlzEtvyy0tR10STNhxiG3EotsBK40NaHHteUfIC+
LbGe+aCiZTvOFO7yVsMnb6tY8TPxEeB4A4Ymqk1/qo0PY01FFFugokqN/ioUXK6gsTAKPqyI9fY7
8r9HsKsO59YLIRGPToH6i43sCONcyvOrkMjuzINdrlkMhlM+hw6I+n2PBhRApeG5HMjnsILMxKY8
JFyt4UxrdK+eSSmuJHBcQJHb4nUxVxzC6IMh6dGdJUHP4R3QZsgZBe6/tq23gdqe8cR4OUD2UKHx
xzbV796aNC3tLaIvWolnndUUt7H1uipHQUnJ7roAMiTi9701NrTMHq2/kX3Ts39Vx/J+pxrgVGMn
juj5YCCX3EzwnBfPeZ5nu2SIEbVyR9t8qSZBaA4OjzDs2f+Ys/5eYni+c8ivTSRSRRAdubGguciR
CbLbfIYrkRXiKa+qX8OAmUsjIsRr849gIyba+VkdV55qqsX0Nbluoj01oepAqQi+DwsEhQ+nco60
v1v7fHtlD2cLlGXWpRorX1YyTwG58MJzyLMapzro/A9ukSKjYhpcOxroFwLNTCW7LaTRFsjN/RGF
wJSVnBOxHoQKMRkV4e0O+EiasQOzJousUBHawAwF1iw7i3Dneykw0FF7bfEbds9YFYDUKGnhMO2E
toJLrpchFJtbNpEzy+SMShiPYv/MOy0uo6xuekMAO2chZbgFIZ4XcdUDHstzlh2GzeUJbJlX95iM
QcyU5b0lF2DjHjhLp7QDbmgKE8VkMz1NmSugdATGSmyw4vqIrFYKFuehZUaiXAVPWbQRbTyQPp54
0SZ7NX6hn4qTi2kwktEWb0f6aNh0UdHf77QplfxPWHVD75fneHqnANNePQVgsSJnjj0n2cTYJDGP
SF2cTaMuTiVhtEtQUAG4ihcuDeYW4UxxCYCgjuusOvzNyvWGHNpn41XGthtpoP+mTtirlVD2jznC
Q5TtNp4BSOz8PArG0XFvH1kcp41ZrqyWS18ivFaO1HQoLoiT8OL7AtcjnI8TVSrVgEsEUDv0dmZ/
YlMqJjmJmXstIJ5KzLUFwu6ngWdWKnHH13sDBqjpg3lSrRPWdZ++QWueSlNhEStO/Gv7BPgfnpHV
ugjZvpWw0bMLC+9dw2x/W8s16kRMM10uj0IwPECiq/HTwuxEeWCsPcWarxX0B6/h0iIt+miyHwTo
in5nXUnNOX5zsoHi4riZ2yt3Sv43bPdJhurMPmCHT7LcdcZyn/YpoXxVpfJXOHKzla1Kce8bcqZB
yCcmUPSVuiC85wXmFvkPebcYw3FrYngVQrAsc71Q/XkmvGK9YEVQNePHo1zGDYOk9dJ+3t1U+Y1r
1E5blcG51j+P7VRhgLRs0ThHR5JyRwPbkdTsx8WyoFTz/XSN6XwkQK4SE9eFf3IogpWPegh9N4xj
fTaPO2Y9p6n8z1/r5civjRf5F9VnQ5MF5JvsucNQEP4GTnaYhNpt19QBP/Ch8dHkxzHvQ7HmV79Y
3utZ6Tof7vI7uOtRCWH85nPkcIfI8Sp/f1LkzJqEqsF2gpbX+DFPfpCqw+KMfqNA2EnP7yhEsf8j
Iwxex7xzqy6LVP/R2diAz4oBYO6+i78FQZc8odwndSRYAi7WlvbC18OAt5+t5Gm/PFBZWWshGewj
Khk950Sx7e3wf3f3bu0p7DjCNgejKMArzSUmP9FjN0Pr2pdwsTLpum8KYWiPUpj+pXKCZx/mXGmf
/3OszBvkChNFTH17TqD+quge9bP7ztc0218mnYAy+WPsOihAj8DqKcioO6aGJBSEdhagECtVLsS+
s/dJVXOYrlcP8gmidvSojdU9TEuYgPLpGAPuuO0WesZ4jzy0Ej0kZaAZpSDOwiWGeJF2gPfDlmZu
GdAtItACt3WARCGgcXmaYEVy/m2/pGZmH/XLCfza82zTMLgTDL8DLIhQq7zZf65aFdvEIuviyAS4
QiVt/rJe6ohosVDfeRM0JaKp/vzJqpEtSJWLAs+QkKCyus63pGXtnj2J2G2GHdNXpbtMQoD758XS
0d1C+j0/XF/wLCJ4iOQWjEv0d+tfRFhyjYfaaObtaPpKzphgeOR+UudebjYxIWJ4/PvmpU7XpB4y
b78xCfBhdMsW/reFiJo6JPUp988IOI6wVVhherFvIZfUVLYpVGd+gwMyMGtXl0y2fbOMjCR3PHh7
w6bUzoHJp4Gv7vlx3ZozuZrYVYtnGbT0e9WACSDGR4BYq9PTpaUj5NIGMzEfqMT5771jBMN80XQy
w8cnHJ9pujUFyWPavr92ju7ILA1pHdXhrNeUMPK81j6v8qx9v16T2HwHBp1d1Z/Q62zTMWb2LWbL
Oplgps1SfV/yMTAIXlZl0fDJl+Qh5cHyafSTQi89yUP9uYfJVuInDXYG2R4XGLJNkKwR9dVDfjxp
CEAgvhyEABxWCG04qy4eUCHZ+Rce8JvdEL74vPDQDwaoXz+hFbjq6VjurprCbyo9gpLFWsJqrQm2
tHuleC7cMOV40nsAtUEfgLfFUUa6AOMHd6zqFHECjWoIdTDy4pLTNERTb2xhCRUUFu5USY4039ny
X2/s5lDAo+F0vAq8IWPkr82jUPzhLZlW08dDQRQ5U5bnHMkuShSuj/w2ZH9VbRwgT1gS2NzUDVoo
4MsRl4YhPIlcHfNTWUZ70rrNIXBSvGYfE056V7VLKLgLdUJgIcs5dzeY1BuBY3AmZKNYaR791Cjx
KQkO7ii0jFtdIZlwsCkZn7qyajAptY1hZxXN3py8qPk9Iqsf7rcHDeb2niTynnoPUAuJcUDVhqVd
TspdhXJqgs5ktbsDS5po+DJJpR4TtnAyQAm5rQ8QHTEnaBNzahmbE/MF8zAPOgcOJOBugLclaogi
O4sJOowHzDQSPUsB7UcGjEj7NW8mjPdLYzS+J/39zvId5UKFT4i2qRgJeIeKZxiNpfQmT7TDuaKH
K5D4w8VqotL/5OGD4NQyccLMxD2EHDN5Xzn8aBWJbxHNXv4gD/c5kM7e716nrZ/0NdCzML/d1ESs
/DdzyII7bffG4WuYahGU1K2nkyktsSSEDjIujtLONGO187rMKtH14go3Oqvvp+oXGbMDAqsQP7Uk
nhO6KI9hTzkcuS9UCffICOxb08j3pEQhwSc2SXazpHi5S5oIrz20ZXzykD+qi/t78aMA1ULor0sE
RocFBIeDIujp4Sx/+yM4oD0MuBihfncyrT9lgKUiYWHxlUqKL+34rUSfspWFyT529qhOdjowMJp9
shFLzO9ggwXREHeDgd4ZZTrWgKqidtd9aZRJ10ZZbiGvFFwIGQt+StZy2nzeamD6omb0qarhIPkd
7w1qKB81li2s86YZInn1GgvpTACGx85PqHeBUv/YaV87WXQvazZAjV3IB8XnM81iDL4VY/SkiC8C
Jh9Zy5K9rWyz6PZf+0wyLVYkvXjM8uFTnimvepADLn289ea3BefPgxVJNwym6FPzUBPEvQFfoJJB
sBjqVTHGuNX4D7ZVnSLuT3SRfDsSGEuV+eaHphhl4ZGlF0TlTR7QbgHkVoOJRipZ7ou46KGWV+VM
dFmQfEQMosG7yU+43HxU7noyCZnLLu7svgmXqE1/CEXVzTAkzDdVsZvb9UXUmktPFzgaKjQJpzjB
22Up8swdIA5guMcUHW2qJ3dtyZxMgRJZgzoz4ql2lY3Jxo2/ADoIEy7TXjlwLNMBp++ZqanmtR66
oUnEs/OBK2GnLJmN/Yp/uebbsQui0wwOCH8k91GIQmj81VnwHTXvCr8XhHBJDlPmJLV7d1cBsZm6
u15YvyBotVH5Erw/GNvai1QW9e/IatH+nqfX1Mxrla9Tf1iNn3AT/IYfRdAujA8izMTZhygHxLd9
cyz8Jh6MNC4CRek2N1V+d5brEK+wfIrkO7sqLr07KerapsxboFva3P0Cwt+AUnTD9VRSXfaL+jL6
5wOzpTs84LImmCblggFNhSNXEgqYWoa83K3n5NEOKxR5KmOs/U0/yVZQ507ZQz3M15D0tMrCrjRu
kRw9+YYLGBilBlslNg+39PPJhQfnKUNdS2eEZenkX5cJPwTuVDlyXq0nnArh9dbTNDC+XtGk4r2n
oocW0+j+Blc21TcGNMGynIac5wBXRmWVhIV+73at0GKOv56jFK+P/TZHLzHtgoLLP3McYWHtLlg8
eMJnvbci7i6h//t1UuWlmQs+rbzEaXmSbvYaJjsg/KIzklwschYLIgAv3Zv3j2XIbNME5LgP90Mc
CSGYY7P0uyjhveTXV2xHwZn9XQhLaLr5DhgbZBgpd9L66NDQsF0spCOW/w51EJ+dlHLpdzC82Uel
QI87oRk368naNjaa1c6jyjpIFUNxCsDidkmXB9hUYDVAU2M6M561QTS6zu8Ohk2k+Vz0vSJ3264y
F0MW0OxhzuelgXUNucNEgylZU9Qpcu2S7Uti9X0OrABOzPkISehIFEN7/sD8ijxCQReaXNZofFXn
HV42UPlXY545lkz98E/rTnm643J1qQrn+upbd3wK50q9mOutVfi65kc4Xb23uR11DDvV3IgmTp1E
qDvgzEJzMgVVNe6IvzLJsb3KKZnU6XS92rHYG6A1QScwcHSD2kaZbEeYPN5bTq7+TWzSpi3YPCKT
pLTVc7AE7uzL7HSpCdsCgLv5I2URWks+ogkJiPX1vG1PKf46bqeijKtVdB9DJ5EW4TojoDu20iLG
VeVpGkP4OuCNOH98eeCBnqKUebWqyO9GpicPNWzb2VgHtHXQpW8rXJYwSgArxi/9eGWhoP5kYaRd
+VKcEy5Jjo4u6C8Q4B//eXFQQJu/qRzrb3S9P1mmQjeq6zKDxmKdf0SGWQ/livZEzJapYq/Yphsv
oye1ctbPX03Uy/N3NOsO9YaiaAaDUOZ+5ZJdwgFePJJLiwH+XAaoW7RbAHICYtS0JzVJ71/slYHA
unLx7DlP6s0w4lRzkYkjmfb7wo3/0jDWD6ZczKu2E83OotVJ6I4I5y19BxHLL1HVsu1Tf6O4HSLB
1vsBoDbYEkfGhtbmsPbUJqAyNuMJgbA2J1+iDhXo/XO45a1JiuNi98j23jcdYZRKRg/My6CTWYXC
vggyeCvpU+qiDUvBbjQK6iTDA/brvbrKOqBCwsl2WCe0y71FmV98H4h2KsNTFBl2d2BuLBJtodyb
uYn2db2F5WK/wsg06y0ZGYaqcY8dmx6cPh+n5pKXKDl2uL+ZeaUdKu/nuedtqI/SS0vvwjdAelJM
9tIP6z9jMQGzDWxpX0pX5pkrzs7cXSQM0L4sJLx90FCPF0XXi2LBB4bNr0dlvgYka4AKYhvlSUDn
InXRhdMe2Xb/dvAu99Ifi63084ydAS65B/DYdz5NVAvbEqWpp62pWcEE5vZO+92w8pYhQE+9/mNJ
DEoW+PHWp4899ceondsmrIpHWMaLFOnTVgIKfHhQhX6djjunWPmsSP3xZ2WoUYqafJohxpzyCggQ
B8zGE7k0aXvMyYQykHko9HiY1rNDAhXWx+6UgOQSvftiNmR3e6tc80Ub3XvHKyOB+U+jsU9bkBUw
wQavga+3JMlKL9PAYYn1Ruz+ck+jwNwrfTGli1uLXBgs1zHfpbNw6PYqNDB/X/QWQ0wtFbDVnDX5
Uj3vLX6mhfP8/LYQQRd+4xfXeCNjuRMA96LfBQIuH29NjzcuUntrWRftsBQryQcyPyi9rvrnqh3X
KVi6N2wioWF/8trhmQWbwxwQw09sfSEnEmN8nvoW2IvWsP8TWbnmE/5GeX7+BHo5k36k9XHByuVJ
3tVaXidh0JHvbqxhcoYsRKGJbNZjU9431pC7JOyGeASmmGHVqhwzBkL4awZ3J+9zbvepc+dHGpuJ
JmWVQYoMCAqoXlBbxUQH12xzlfrPprcTn/6MRJEKxN2+7Upwv64pNkjvk3sjPyMa7+5AHu7Hygv3
2gwv5HIJUPI7yeYhp1FkIQ6msseknupCZWxjGSjH4PXP7etUoTglRw4xKmqXSGZRRRY5O19j4Hl7
n3dq6/iLP5ssm966C7sUH4KG1mxcTa3s6sJ2NX5vh7+MEM7u8+dt6oQPfOPIrNGRRwFHC2hhYqUY
0kAoZJyl/MY0sh1tynNn6paApfYISUsTJfMTvVbYfM7hqP5Ex2SBQgZBddLVmMEpmHDyoa6hdQup
MyAu8ADpfEYRrr9ZGOF0/6ElyGqGD3ZcD70FRqJvkH8KEBfeKH2DxL00e9RyguWKrBtVZjjkes1x
UTs2+oJnyQnyMwHa9+Ov67yAgqWjKHepTjNM5cz1hYhoQIG+lPIbTyK+9l2NlO59EjMsklmLqKpo
9sQym7wzote69ko89WXylhwlvEx9RUJKjCtCVJOB176vhxtiwy9be1FgTfrfywj302znDfmJAOWr
oTT+TYT8Zrt5cEDp2/h6G9DLTwZSpu6RlVdsN+oEsx4JCgQDy08jxFyF8EMkYbmAI9qiECFaz2tj
H9MPvUytiP9SBxxXc/BsO0P10tWko1uyiskiW2G8j38tRkh4AxWNk2gvSb6kPi/z408o6b06r5ra
e2YYDkRdZjDnAUvrhHm7DVRoJjNZavPnG7db5UBeIUMiZZAdRDuOu4Gs+rb2SiltpmKDst94plkt
FT2h5ooiZK/BDsdKEZhFLSGRA/NnHw9GKvutQ3FoUoDGykEXf8h5L6QyLdEAYuO6XIftHl/7ltbF
6OXmLosESG9b8HmDNVMvF+nZ1LUAa0nCTWLrSilzvLQf4MRDMYdEmFhffz1utBT1GDlaE7gEDjPE
xYKJ3Ep9pwMSXtinewqbDm8sP91vYjjJjZEMvI9yyGIt0kA5/PpatT+sm5xwP64nw1QwM6olyxUp
GfVrMcb1gddieOt8rdti+k7YTJvheuBAtPA+TjPr57JfKIZF0gC/etud9ZNp8GvmNdFjxqIwlHcz
rrN6V8re4saBGIADAmb1xlBj1kuKHqfv8PJHk1JL3TjJxJ1CgLSnRqRak5lMcKmzhJ8ob0Y6BSXR
sx5ks1VD222dgHhDJdkh8DMfQglzI98BP9Fe9UiAwETgpLHewQThdluND1JPGM7VNgbIey1rfuYh
NDUfO4JkLDytbz06PiIkju4/jJ3/SMbFvhMx4mXhD2k31APgDDYfCckLduxjxMFRnGIgzSb/nKxi
eqT/4LhZtCqkAfT1eIERlp680LGMFgO/ZrtFuutnlMyZViccMK9c6FKFFP6krYZdawTJbU3BGl6V
R6ACnuGG2vvi0GUgnBALrCCDvmeDIt4oOleqbE1HYvPF3NO0EEtDwdMnsjBYagCj1DsdrurgNyCx
R6vWk/pud27WW+K9wlr3DcKn6ZwXD2YUOxHiqhHJ7fJc5VqmoOnyNT12+u1CLoZWAkAkAK8s7PhP
tM59q22TbQqEHmbkRx2QrRJgVDLK3eSVNDGgO9teBkao8VzBmzbisolZc2yqv9qmKojATJq135M8
XoKpsXskNrw4w0LSsY9rYTgWe1KlLic8/iZBx2Mc9LB1xsvNmfSB7cIyBwqBTs4EFjEUH2OpTW92
KkVFnlZb2/qKgz/qdLJg8y0MTz1Cq2DNN131kATMddNW6v0RxGaIFbAdWjW0zVViKlKPIMHHrbsH
bz4ZgKKAp3gkH/4bJHLoCSBSohnqN7ik+KgG5DYg4TVXI8yMz9froJzgXhf5PvDW9mtX/ZDySdTO
0K21N1MxodUl6ZAdvj4PBe/M0tdcZXn2P6RYjUM9fqcTFyJc8Pr+Go6N1Ztn8v/cckUAXoLCfh2d
FWmLzVGsVQK1XZG7+cDfjca55Omf/ocvd6Rz6dy4kz5tHUe8JAPQ4YC2ZTkLj1fGpOF3hJAYK4vq
5ai/85dVRFREJW+Qy7KN/3TsdS1kZa1wstAdsTbnyDvlbF4z0e7dTkUgxSu0N4bn6loZ2KEwaf+3
nCOH14nQnuvORg8ZV46VOcoL4QPDY6+CqZMREYnRI1UId+t0OOmqciAz/QmWIZ/T78iQqzagnc4Z
njnTMG2RpGqqFqyRKQytnqLY8Z7zc19j/QPGKOtGnY/v0nXyPNObgvvf/nNesoipPzsrl9O9XyD6
RaBHYlk3T9eqb2nqSWKCNb4WpDNRjtdT9BM03diTXFs24/sLllsRgnIWqSFQUOQJ9vSoYdPT6fbl
ZlGTd+QyAfpShYwT0R0VLVtARetonhRNS+uiDWuI55WyjnjqEDuNXrHFjA3sx+E8Y+eUJ4smfaMO
BFadJAV9tacU88LnzoKlxPMpBxSD1VeN1tXXOkVAchWiDu9b+wJLcZHCC0iWPMQl8Ifvf3j21lI1
4LHMzadIIyGEo2pnw9hDwhjz+gzDxRDJbkh/k8/jy+/0azAuBel0/ApLamoYvsyPp2ZcxE3x0LxC
K/MWO+QKFJzIBIRbWxmLR2HMQS0xxOuNMGdSmceqIgrDB9CPq7wPN4+i2zgmEqRbmUSANzhLt3bF
YXQOGsbe6WlRep0W9SIWgi+gGmCFMMVtF5fKEkKzdMyc6qJrTSDLQlG4EVeftLgJtNWgpxfugpTZ
pOrU5qzkuAPHgVaoHWM6eW4ya+ZWbxvvUmLHd5rx5o5WdBUfl+/W24IFvq1LMscHZtohkOr3sH96
nlvQyc1C2ceUWXNY6NyiQYaAzXv5R2zMmEQ71qrJlQwAerEFiZpYPIdkgPjg/fMEKZ2OGPd/bq/W
Y4MC+rMvoM5Zao5s+b5GhWrq8jQYT5PZ/ZDsBO7WznQGI+OND5Me1I2jcMJCqKFVUTSdAIRFnQwA
QxnHt+yuG49X60tsQOhgCq4FjRcbP5UcD724Mbk6rSFw45T/I66VnaR4kKqefgZLyrT6XA1NXDcj
eA1tetkTx9wQS9kaPGZAXkqcyA/XYVkYF4o+VuYOWFLO9ABWKC7Ud3vLnSWAKWwP5MBGpGTN1FM1
N7t6gzC5z7APVCJ1IkHL81OS17EWeNqP3KN+vGfEyqX7Iyt3MTrBahLiNbCNNgZ9PFsM3b6jfsUC
K+hrP51HuSZitfAVVKkKpup//MND5IF7xHfg30G64uDT+8E3rbLFpaQFY4N7FktUsMpBOywhlU6L
PN6WSlg4FY8bJbK6XdfV4HgiScoW+vJUaRI5CGiP4Zfu+W1TRNriQt2iptyGSiCR5UkCPgh63U3f
YcbdzzfnWNBxGrm1iVi5+xj85AJX5GgZ6pb1kfzFUmEUZuv/MR2IwKLlph/OdAXe05VQ2Slkp7Lw
I7Y2IfBhHEcvyaI+GcOsPbVElTVUM633x2SuXL/Uze1L07HXlGnHOA7CvcHRPd4PlNLxd9JEXx7K
kBplnzoAleEGl7wxO1HVR3lEYp/dPKNEDDEkJxGOaQvRe804ikuQYS+bIK047e19BEGp5rJnBDjL
g5WQ7TUUmESSBlS+pn+H4bgB22ZzvcYYyECcmHVRgo98iKlZCLmATZ7NTBHDPrm792fxEc9oyI1F
WvF8GaJxDVgtnb7yi5sYYuesg+5PhtQ2znPE+A33aV2x9FvKyhzghiSL4Aega/3oqjEgjzFJbEK9
W2hFWaRiFQURCID1s3UcwwvlLcJb1Q+ajoXrjrTzG3aXvPcPj+ULuJZrwtNUYNzDHyWxxvzx/Q63
AbeDf8yeaDzs+DTwZS9T21wR7IJ0dvnntfIZIOstrgpU3kCzVnYFgy2ckfYoW4sXkUYvOPxto99V
92woFD6ZQV6ingwKLorNoYgPKMLJ5NSou8n//A82unAXS/iTocR6YVVdfLd32OOJbtJi6HScw0po
PWdpd0RvwxbFVJnCbgZfcamdDozs05n1ky/emGqq0DwM2mqUD9o1aqlSCUuKmz+IAOA4ZisfVOuw
nWuU8xYxlZm0P8lyBmYFCIHwjwqAy4qTRfXPbB4M2TOysmqgsOiig6evVeQwfZOYsg0EaN7cbqXI
ekbD536xk2o6YffPQQnjQ02eZsP2I7FzyCOv0X2lmn75mhqF38GUexpiFP/Zon+JFfPXEjZ7wnSr
fPvE5Hduc3l1AI/7i+81Hpz3uRb06s+fwyko+tEPaT/KYz7wRO+o+O8/CfIl50gDKHVOe96XR8uJ
YMf7QwPXHkYa2ENyKoxUl6kYuYPjOzcR9qbNmhc9QLhBuysVFv2XDUo/JncIgm6MUxpoJcX1NWBR
yionD9OHkQxr7VzIGHa3T37lPMqD1IQA8okcsTgFmQFkCiyJs7UF5rVrmJO6p3sjuXrovVXIsXH+
dVvPf8jharuHy/9WHpcT2ExCduCeBRQRQcInRsSV969Ra4itY9sEF5nizPT4ZsxhIAnQo4+BBDqj
h8H1JNJgDYyhJ1NrcMBLI1Y8Qa5mhrdsEaKZAMtje3j+ZVeC4qZYlXcXA9tvsu52yVrOEThtoMxc
C/vM2j52xiAjnPEZuNBDhATt9LPM+pO0IgvyjbQ3hva/mg9Y5wf+7RP8Ldl5ya/JNQyr19ys/Tya
K29hnzcSrkec9tB2TgSoBW6NHX2BHKC1b9opehyt1w+ieFdooMB3PpA42G9rejkkjh/T3qdFJFmS
Mb8fSVq9YT2PTsD50lK/paUsk6OLAtt3ITgqIjUbEOdk9U3ki2IxnszMpncT2faL4tfwO1EN6m/z
Wt33jOI24k0794iXOnIjPh+BAW8+6tG7rjiou0eycPtXffL1q5E74HADx1IsPYye9+blipyEmeNj
vS7JOV+h8iF2uyqpil8Vl1YFGcKMbg9nomCQti1GS2E9UCR35ibIInhB/CaxHcUe6XAB6k2BFWE8
OATH4gSxOS5laz6wcvU3OfqxwG0ErVudofQ8zxfh6PtGCfnXg/3P9EXZPX/0yRknGG83xn+X3QMR
I7NrzCYZPSpT2oMyzDxgmDBzQU3I4btm6vDcCpISkhrvyhf/6SpUVETJXO4piaCGJyiQGIQ/4dy4
D8sUaO8PZxQA5JkE5uZSHuhnPTdOSaZ5LYvG5RAYLj62Ee/JzVf9Hg+Hh0vbl+ugS4Ymmd8eRVYL
P+euk4UEAzD3TYxJ6v70uA/zumFRTrl8XZc4yDSPa1XRszehzx+tdiQs9azyYz4BJ3+KFsJb9S1Q
eO0UEtStSIfHjtmcusJau0ByWuzXfZxD+UZlTJ0CjDtyPGWYNiCunvnx/oiszBx3iThHyNit9wRo
guZn2AKtF5Ivm7SklDS79NyiAnvo0E8M0rsiyR/ioDjZ9jWm6JZjDm0NqcKvFFB1KKzJDGDUcDFK
yoW3OizUdgp044BWNMSXU7yk+kJ648JZBDRKgtDegiMuZtcxs0NWFuy7E4w5FCiE4uqtb1fuP9g9
gtr3W5mG+Au4pDSW8Vdn6kExOORW7Q1OSlaCHxmtKydCvtlnCnG3OnvpzRXDXioDE145+dUBEca8
CLbVNFgcAXnU0gRDw0625C6X/yOFJLSNTjkuQbhOZKCB/1LO2Em9wwuZewdd6VJa0AosLumwsp+c
EPGS6x2ynxQpnfFSeuEMlDbDqTaBlLCUb8G3UmZiJdenvxl7NBmRlmYZ4vLEetpYfRxm5G8zDLYT
YPQlDckPPwDxeQSoDagT/iMJozPo6C3N+c9XNaLRckL+FMiujVPISGw4aphmTP95r72qMu3oPAR2
v6+rRuulKoBZX6ru6+PCq2SXstrr0ob2j+M7oUpsSdkG57e5Yal1wQ4IYCQUI2rWkts+0mjVeOll
rFerGtTB9x221xg7iP4siuoEgko/gj9PLZnpGgKSNiCS40jd+EtjAPf24aqAFPB1w3rWJsqPzIpL
wkCeygN583Q3Yb4feifrDKGXVfN6VJ3pg+Cs7yLGj0qQ7/H+XRLPOOe8uIseK9RR+TCsu6lRB6LB
pQMmJFL6nHhN9P5jS0tljiKwydlQZRsMDN3xKwVewno7r9d3TufHpnRJZo5I0du0xwig+3sBa9Uw
uPyKrwPDWEYajh0D0d4eikDIiYxEEZ6rFWpr/PVF8l4gL7vp5rPj6NEyCBBDmBdg2APnS71fgvfn
zizPxYimoJDybArZJgVAl1qAvMybjC/sEi3iNGsR1CTPxG/RAELB+V6Eo5Dy6+mlGMi6SDjEUeJv
5Wf7OvcOk0olkmm8FjIlTSc37sjlDmORYgurDo5USzcrCNYCt6ITE++MG1VyM7gGxb3ithMtscS2
D3Cj9heF+ejXv7+TqSbJcx9DRu9qrmVty/5yIZjneP3dolaeyfPRlo4DJOkLVg9985bthKv3XLRf
TANjpMqMngiGY5QbtxVna9xjpw3RJP8Ew2InUa3jxtC4NrI27Is2jRkk5V6XOUs7l7pHAHqRBUGE
K9MARZ7uW6MYGCjRilMvTugNWW5n/thL5uCR6+4mT3rkIsKPz73bNCueo38FEje+i+NRu38y3cwX
Wy/qobtxh2fkwEJ/yc/vT57KP2h3/K12lgiSsUBtDrxkinqIs32NmlI7fCY3u8HjuWKQklpUfguR
XZiEQF4RNBqXj7uCLntjKx7mZ9/ZAXRMjz0CduUY4IdGxWkWGVDw/5p50mUqbMd1Rqts6y0ibYYM
7XPZTzyejaCPqD4hUxFdZCvtY6c6dS6IfTihMXCZpzvML8VsCh5IObuo1PS0rbsOy2vQBOym5ElD
aHLl6U+f8vCUfHNWaBVnVFSVipB0j6fz79MaqjEKbU66a3jkTw2aHYHAN/JUL+BQxcFWsH9tLPVd
3EIXKt4cqdDqRTMFWZs/wxEuknzLVsuaToAg/EqdOqF0xKlwVj3K1Mkmqi/gYojnYJ0QNPFQ1C8Y
4tUHqNKJ5L1LKVOjQCm4Nl6hAMxGkLOL6C/G5g3ljHKw0heBtIlxPelnvfsW947aB/yUMSG5ghli
fAf8q+trJ991lFqNs+iJ2bYcixU/GfFkojXBK2BiD8VgTejA2idvwelnmsc417tODZUAN48E22Nc
IX8Pr49JrqssCuK14tLcivTjXM34JVyul1yopuopHtGJTHmfZGtFtJj+v5+7zsVqm+fXrNZL34s5
9GMutDRLBHxGFgak0O/0lO66k7NXhtdQdD0TM7pZqfgq4QiciAiJPmqLXyTNGRqHiqPp71hZiyga
pgVhLRGfxu9IB6awnZbl9dUp/Z/fvChFlpIKxdJRG3F9Pqy8J3swEsTnOiZ3xFz3FqrJs08gNaKt
FfhsBGfcmnUfA1LYrp4XpKIjbSzzxPj5C8peV7uMrcnWC7+oZbWGUej5tvaHOw3QFEysWKqyzrTr
EEygecS1e+aerKHx6iu3jqxJFHExO2bWI3ygF1fo30hsGOD1bEGmH/jBNC9p4idVMrYc360kNJdV
sbF1YRknWT5lW9+gRqwUqESAnoePb+6gbmRQvETrRhjtGrnW5OQM/qiWnMXPw81rI7drNyL2JyiZ
rrd5Dz16JBnQD28GZwrYbJe93GvC6Ep5or4f7j1XegBwhFPydc07KQzm48Eih7zsl1EI01A0ukET
r66xizUttmASpmCnjtSkOtMyx3Hvg3yKUJc8S/2pncSgmymIWGP/Rvm8Ds9GUAGOCeBQ876s3/Vi
VixZv72g5SgtoKznrN9h4fOJmvOWrUlZA+njFvFEIIP+Ey5iZlLLVdXa91VskcM/do+EnqDrHh0x
33Vt/LwonReUC7YcjTa+tIizN6CqGSvmGiv/VaGLtty8L1HGCyaYjH0Nc/3JuahEgwVaBRJJQrYr
6YYEdZt+qGMAUlGRzximwuRRnewgqUQXdaSTD3BGyrRKEE5DIZ4gKw7blnRqbLdCmfFcPskh28f8
tHd4F0AMiOdU4/Y0lObEtD/5EyBwRwhheVpTvqQWCalovo4RW1T6AmqdMnf/rI3oMx9Cq/ZxHz3C
efO7xSaANSgSXUKT6uwTrQxGWIi035Hq2ZxXoghRIRBP6K7pN21TDLCZI0GXjWJ7P6b5VTYDJpz0
wrjxIWzRZkLWUlEJf3tEcrYEQ0meVX92moiM02FId0GAXvqRycd52PZO8NqMrfKOEj/yL3SsTA4E
4TwFz386r19Jp7lLzfU6NAIGqI0Puyb2NJKjyyN5RPRhd2tJaVZSlCYFnKonOCdquSSqw4zWKYSD
adcmkTyCqqVWXOI8MOUjxHhCqu4Pp0B5dNO+AcpjVi4jp82Dix8kLFq5PiB3je8mPDv5Vs4mbSGx
v+/4PsZyeB6/MrmwkfJgMYCw2QTjnu8moXrpP5RpqHu8pHXB+WJnU8xd34eryxAOqxL4TCTn6sjN
JH9hMCM7qLlxidNofM5Quvf6X1Fund8/e7HEQk+yTTPd5BNxkEio0UhatjKKJd6RCSb26urqW3X7
EK9u1N9GGUkjpV3qcX2aHKuEUzGuCJrr4qHmUUsZKrlbprR3CBXXyFTG12ShNeoSdYBHysw81yXS
vjHAWSZ5lsFk4b65SiQHiBYI14JfO8qlBwuVlwvBoa8wQkQFlFVrdvWeQhb5rAST460R6IEOCNjN
WkIqmcW6TGiHPKhk0Jt9EksWkbjZM++VL6HcIPpDsPslbUr6fLTqHDI34fruBS+6XZWK62s5gyuZ
uFarmLcpofExjaJYyE4ZYQ47rMlAiqz8EEYET53BZgoTGOWZt0OVyu8XhN3lVEzGPz5ZHLp69JMO
fWPu6NJGmsanvbQiwRKTGS5zBh/BaiI4d2QRAdB3wL8AfIe2AC6ziXKSsL+A7JO947ZWpoHXKQgI
965nrbWBEnGLOpgEPqkNXnKsk4XP/jTGNv4nG983YVe0BMGLYtuMi4OB2SOE1oYaBb+mM/0CSfMN
99r9vfYmmRIoUrIJukap4G+Ap73fwe/n3oiPIsGmSt01sjheeB+Q2tEHQUiL7Y7D+N/0nIXWd6hs
Ewts8zZLU2EIDwYySJEmHFDnhPY3su3ZuTrTFih3UiV1gKuFv5XnJlQZo/6RJkt7BdbeW136r5Vd
lWqoGeJiQ7K1YCASjlT9B9wIXJBzQrLTLUb3jK7F0uGG0OWthjRJ2AAx/8Ejs/7iElOuHdkVEApw
VxwtnAUJKPutBrvxD4473oKnH3a6ufwOsJnri+SVqInqaL0dTVys+IVhMve7hCGR7kD+BoNvuFeh
+n+q0boVAMRAKYh2goD4iT60ho7K/YULRa97tcrHCZNCNGdbFp9oBUhR11/rLYlIpiBJ1MPHHOvZ
Zc61Yh0Ld33ZLM4QUJC3n4Egkuxl/nt78EIVuU86bdgp3+L7CZvPubInhih9GU6pKkvJT14/43bu
qkIb6BmUMUV6AZj9AsFD49Ebx1kSByzD67PqdNBB7kZRWV0TWEiXXmvdrfIfBQSct3EPC8RSa5ZX
/sChkBTCEXygh1HcY0sl4QiJP6NL5uDn8cc1vKCRLzS1rjbjqoOB93LlP2oY42V4ZtSetLi5+TIt
OixCuk1beOnUJmaUAVGLZ8abY7+FUNN5Rc2NDtGJ/3ExptcyaUfXfdklC8W1vn9JSqVTQayuDxnj
qew2DbKsoTtwUJME97vuig+IMCaI6t6Pv3R2hWg4CEGNUZRh+VN9MHCbqzH1iHGyFtyiOBRdqgsU
mu6CLnw0zBo9AiOpe+8pWF9xb9RM2hTzSncbbaAqik8zuMJQC7wK59/PlgMPf5KvrEzcSfFLouUe
SE24+3VmI/O063bRtGil2v+ZdN8vBuOie98YQVOB6TwNbv2+vN9A5eR3msZbBT7Uip78p5Re5sQc
69JxCTyHz/UVIyPT4MEzcT5tSe+JT+msXagjfMeiUjZPR7ffzay551zi2e7P56O0H6dnyk1lo/WJ
6t8rEif4pWPC708k9Erj1soq5YtjMLH/SnKuGw0SDbp25I+f60m8tXWbi3IpoCGvN6UDRRSss/G+
7H3h5KYwpnSjxxK56CRuE8mP3ELgywMMEQlxNtj3RFy6IVsJZ6d1PspcTp+lQzJw8+3MucxzHzZN
BCHE/yWuNPVo16s1lbmOzB3UNk6n4ninu0VB/ghrFvPoJpKr+9gqc0vyw99PAbkZBsmOgM4IuH7W
1/mH3adRjkuwJWIQD1ZaY3+/CJk37ox/GHr/087DrZ2HTz7eENrUJaXHC5hbtWCif7WiwZndqpVy
Cpdrn+zmjFS/v33PMjImlt6xvLXJ8v06XPaOlBYH388oU2PTGY0Zl7otH4FG2f8eYp3WxsrBUGP4
qprVaBRIHALRPSsxXi1bTJxpWns9eUteRnXLFKHS0c5d6M9QKU14ha3Lq/bBZzwCAY3avIyS4KaG
WGMDH04unJF1frLRnc2AX6c/c38QL9xF3UNXxfVp7H4ARIMKqgljVI8QwSxCOra4SJjgah51/whB
VyofN1H24FQpAnzYgZiUCG2F10MphGtps4EJrylSl7AU9R5DZDqNfZUMmVlHhqEdulgswk2lqrKP
iRk9DUZfkcevCvQeux7h6ImFsYJq/w8YW2Eo2NWokwuP9x0MPXYjXcZHppHWJ4pJDcoYpxaqyVxs
Dc63xjPbtG7hYJCBS9bUGGeFsWrJfMs0FwLCg9LSO0qpczFlLn67r7WUsF3t7ijXf+dMdERC+QDp
aVXIEt2XWd/ZX9Y06l1ZfdEqz4hB71SLoEPHgPLLpDOHpipZN9MuP7pKCQztMkN8OiEW7HnRTGg8
2Nu6gtOzF2liK5ODSNmwY9C2418n264t0+B52aR9q51YnvjnwNjZLTh7lzS3a0aX3k7cmDebfSd3
kyhWPzVP5RI9p0Be2i1OVxZQ7PNK9blwPmASb1WiPsu2S8N5fFPudTGuYVl4cPMQor7CIAEi5mVh
6VPUGfEd+bYzRQn2k4qEKAKQ1/k4l1WO/DeJ83hJqn40x3GnR4k+Ru1jTBwpgNSBxfWh4EDF8Gdn
nCeQfNSd4QXQ5FOlfGW4q4dbeJKZX6GHnnfCTi0ORypzV0iW4NhWu8e9eA6e3Lpw3/8HSvGFQZP8
nBTMqmQJr5UsaR2SIHSklCrFIS/4+C9syibf5xDz21FNuONbn4CtJ363YhX+W4/2sQe06g30/SnT
Ia4u9wOyPXWr8+SaszNJtLkLPcCAloDOdfBF2Ajc2R8V4mmUZw1WA6mpm/NzJq0OO0CvSkfVKNtH
GSREzGuBY/m/Rf3+JjBpZC+t+Mi7jCLitrr3H0H2+NMH6NVG+/MvSjwZfsPxkJuS4atDbfC9MpR2
HjS0gIW+XiLzaNtp+Mq40DLyY9q4c54YlwezKp6a9JS3G+RCyibgTo+K/VfMc/3lmS4PKEB9JRwN
9ibfoTaglmho4xNjhbPztUtXjrjXJKqf0sTFSTTotzKPsMBj3gHOK2twxywbKD4puqoCY8dMtjcV
IWBEMMke0KR1tSQKXwdr6iILvVPAEKi3pn6Bpvo4fTx9It/hgQFq/JW2Xh8/pe2zbfOOSKXaCaPi
RBTj8nDWbdUCm2mIqy5u8mQRMMV/7DV4twPv+LDdL1yqQtLObMl0jLxtwNxKvlSAdy2HOazRI9Fj
sxoKo1Xvw3BtlFPs4EPBVVmoZ+bylMOV4K+7ZoVig18cv0e+BOYM0ahBFcT08WX3RxFurPnWZBd6
+iL9KwYERHE9a5AU117XVml84VqrOR+nVq5tl5fhh+2dQD9sW70Fc6Y6LtxAcD8zdXmsi2K29WZ0
zBUi6diY1xX8bnxFEhsvufg8uh3MeOF7yT8/ww+oSOX6r2Boy/8e0SjrBtej8rH8AmoQuK2Kazra
EmPRIY7ymDgtWcgkAeYphIgQCx1EWP2t7vkpFC/iAtQClpAU6Ms3fMkqj2ffrEGgcwQ1zQf5CGd2
8leJ/sW8zuucssHSqIU1sOC/2azeooDb06dWiP0qeaWvneP4feL8tK9jOsSCeDqKuP/q2zPRdaNf
Y0EMwYFZWln0L+cy5ZHJvwSBFyXFbAa0Alz91clwspnxvLRfheabQKoZEHdvrHORO31zX1CFXjlt
n2RN2owkXKt07G4a0rIXHqhS50NG8k9DgtnaWpZpovjPZnbWMLSEutF1xgV3Qb+DjlAsPOlwCtKa
JRKVzheRQzPyLtmI+LHF5Fak+HWOVFxXggTRaaK/7Gopy6HaN7jqLDVyvTqnXJNU3iqFTKQZ2Yej
5aEGEYXsCUpTVOo3lJWfTeFTDG6kYiuuQinmbhEB1SFWHjbiIPd47HhKeHJCV7945UGB55y1cM/K
aXso2aD9xDoiGs5EniO+q7Xf8X+o7fio9HYswHzQj0rYvzGrE2is6/fOdbjrownEtjMDZUD2SdJM
704bW2eyvwivd/ZW0PMizIo9bQ3gXPEHpCpsti2lx5gtcTIwcKuKNgezRwEBqRb7w+TQE8HG+say
It1ky/f+ATevG/hAp2DHJa5k1ltH7VkaCOlV9oDpwirwAgrt3EkYyWwAAJIaiIHGoOK5Jgn4Sq2c
aCUpVMlJnn8+wBJMpg/wqZost1EofAZ6yMu2EpHTyTVuWGnYpN5O7KGNqgd/8/cMl+fl7X48pSSc
K2VcajMphiCYWd6IOTKnByitntBL5sigebI4L34cUqr5gwFrPtyZuqlZLIJJWkrAiRmCRrXU5JRo
TODf8p/0KHH9PJBwv9jNCU5Qq1pcTwOqO7enCmeXQ/YAC1i7WqUHscvv5uXCIaIeKdby6vZzG7hD
kQHuUHxHipkmU8XhbNIqMMZ1uYLr369s6tTOhdvwlHrv4llZY+ABdvQF88SXSuaKTdt4ynspLXCj
ljBnektNzikfUqrsdX04JBgYAJLENsGwpWq/Ph6FrT1RIOm2vHeIp540uf263nyLy1hsZ7RdWnUv
Qov4SS5qRQYSN79gQcrGvYTLFurqFQtW5tTy+HFctzMrJrtpkt0M5bpP2JxBI8rIO3h7IpCr6Fa2
v2h95aRrD+xyiiE2BmRrUbRe3URMmjNdjxVWT+VG3tgYtfuplbUA7iurhy2lpWPOY0ZSMSfzhH6F
duii4o9OQ3G5RT+yT/0H4esprmZncVDLZNul1QK8M8V/MzIw8PMyr6LVSsI8Hj0G1lIz/z5Lx1iy
DaTNUCG16y0QxmEmobQOL/T5bSvgZG4aPcZKYp++6SUPUgzj7JH8qX4fVoSjLEbRMnQmB/jJlDsk
T5j2GiXo8vWUEgXKSGItHyVN6dGImerWwIo2osHQXkQ02CK5lgDhUtseuFsACBXjfixQw8irS64x
gva6wkF8NwMiLkCYn/CDEzOJthQ/IAhz8T6W46ZLSqZTDTB8xZ21ihpwSEWCW3WC6eydrrY/rlWG
ywLM4+Gtb6JkAzE+3sgVYD2lkvkZZFYwV8IVZz//dzl0E0utwsCn6r34GTTtcTRCQ40+VVtXCGJc
BgcdYt7gM9LGifpx+Nax8Bgez2UUAS1uVzgj86IEQfFsnb2P7uRgm/h2T+6bPS9Yhbgg0tvId8YN
og41B1D2rWZCtDHEFOi2VZ2GnsL+faCjO9X6oN+iRIBEq0+mpYnLa8tAnx6FWQA343HJOM019++T
ParpvEJUv5GEn8NstJhVRpG6Ssf2C6ww3cbOtD7nn0HqyZ3Zynd4NW2GjCMKNq9YFQUk6Ju/L40k
KCHaDeI1KJ0+5jJuj0tJVacXDJqi5WYjI26c15kWwXQkFvqh0Gg7LKp6oSf2RXpCcN7+cDXnkO4B
wiFo0WvE2wQOfX+09+zeLVRYaRU9+ixkMRvjSOMC3RsiDEl6CQAQC0K6QO6Jyg8QwRJjNFh6BWdp
fbxk07m+mXErlUF4R3hRwlsE5vpB3cIUnXyeadvjIVttApyvmU8NMhsXewFmyxSsikyfKHskZE0x
2KQfOZvspEj3uSaxsZHe7ow8MKDW9EUhVy0AIt4uC42iAbvR8t64s4k/6RFfZUlqgrhJwR+wBUI9
VSMFYPDif953hivRoNBimk7eyFU9CjXNDFXPlWtjpmFx0CN5WQSL9QmPqw+hafuxmtc54tI1YBB0
FnbW4YoQE00LebK72xRCTzz4avtudqkANJShO74JIsIV7PmZarvXqSC2b9EQ/e0+o9AjkkdBmgo+
K4ip5WgqMMV0Sd/NHITwECEmBrREzIjzpDg0tdnl6tedbvOocxVTv/9oPjjnoMOxd/r6gVhJSFOC
xaRdpPMQ4SujomuCU10WFbPzIIEYf7boIW6jUlYwdZWdbmnaYEBZ+MVBzqarfmOGIZUwegML/81I
jlCSESs30CBPEkPjukASUl6x48C3TkDzwaHC0SNQaZJN2i/AdRdjsKalnwKF0Q/Do02avYW5+PE2
93+WEj+chtyjyQY5MnBsHJGYccFgL1kr+15Jo/5OW3ssk/8wBHZtfZQB07uYxdhElFiShHhXebdW
xqg0aOVHi8auGaWs2/z03Rxnd5jdjZWIhPU5sH8YADCuvql22NgdUzplf0C3TdFKhz51ZmyxI+5U
a6u5opMvAbKvjCGUzc3VG2KKpzPGG3n6RmfPXwsVr2Lu1DAKZbqbjOWqxsoa3JIFGUM0O/QjvPEk
w4lUkXmQHwL543slTPCEZqkDUaq6lyIrq28GkxoXrqOZZeDoQhzpTftdEDqlwWK6h/6eJCdfS9Mz
ZanKqgeTWX+Mme0+dRBL5kgTCcYmW3sGWbbred9AxCUg9EjdVprRL4/o+vvqXZyOkoO9mwS6QNH/
1CK5SsQtKCiw18bwDvjfCIFCoJGYFSJXZJ8pAtGLox98Mn+DHpbJXYkBitLEF8EfjS8a1RA2l6hC
6DtzwrzGZsD4AMICEIG3IpuOrgvXacRlSto/ngE6JHAR4KBvGF3AA9ERlJ7l64aMftk4mHxfs8Z3
JQvOpO1Eo4ZWmOytLCNY++NJ9sNXOQkXRm5/+EZWCCKq/mwUhCLh+2HeZGApg7ZTiAAv/J79n7f8
RR6yU4WlK3Zn5hFx4XAhdMYAwLZAm/9Q2Wz8mLyOPEqqN9fVZ+PbItm7kWDmJsz76taI9aXcaZuJ
rmTcnejtspgthncnRo4gMt/W33zwiZPnATfIMydGJ3/MunH/fH6FlERmCfWswHcIHg94XrJjcrVQ
lPKiwNmCZ3C7oOXmNAKkkLqKSNdT6qUt4xs4RZfQmywygRKkBhNpyzWH5XPOumhjq2fyWKUvfOFY
QKGfCAm5Fh1etAxZJnJO5gILjHUeOd6+InDjQwgWOysnCKCtb3OwlaLExitkrsO7H1X1RPOfpJd0
V2FyoBagS4lXtfjMWDDsZtKQXy7IS1E0RHpD+t0VdRBDK5AeztondmwFZ2z1MUMhsCBiBQz8F8QQ
aWl9zKI5ebwC4UkUrGrkoWVXYr/5mAtt1SZcewUtrhcTi7mPb3dVdt1H0YD8SAqQvoqEz8KoPh6o
/PZXYv+pWeNFTsJPI3a/KFnljeW5eQYm+CJcp23qNSmUZHua2IOm6Ed4PYPuZD2NczHAIQid8037
PmW56VXBYw3kv4yzOv+EIEXDm1BzqF0Z3UhCecHpNUqlYtZR7xqekVd6XaAibh1jXq4YocIY5ttA
6h+0A5Q0zu19Ohf/4/W7nHs9Xns3zBoMl2/DmxBcN6W8ABrpvx/EonQPTJNtTgc/+R3pADZ2+EY5
/1PmNS6Egsfp61z/Z6g5f9NOc9g1mOjKPzGpCmv5DXM9W1qPc5H+7apFNAjMwv1uQLEKwDwUAbGY
vPs2/mX+npb7O+MxzamiPB1wHADohLwVZhIy2We0WQxCdS4PcaAZyqg8p/j2wCQojzEGHaeQV7VJ
CMLReWS7+cpKHpNP+R4wD0zEIg1QAAteA/q1tv7r9SHxVhHxMl4RfKyK+P/pwIWpyBTmdn8y3PMh
O5ptmfi0s6uz0uaHQKK77+E7+v7ncH7pDtUBtfjdWFuDpFAC3oFBLcFP0TATpXRZoF6knSSZBnKb
aLZz/WovrMLB7n4a9JXIs30iTIbGcAdgzzbZ9i+D1Wext/bDZwqwrLiW85Md1FPTwhmGHyTsLvQS
Atf1kkCbiVlpxLhvUIe6H3XdBFrpv8wBNERtz6V4p2qMHeK5QvhocxEZ1tHswPeh4yPhuerKZHX7
+CYLLAzbQjYCYjuHgb5+t+Qx2UM9NC9Ew82SaakLvNHZKCrq0QSXlcIm09tU+sxK5VF3XRqB1LbS
MP8G5IrMrFIzPnVLJ1wzrm5oME+25Hj4FAKv4Sc9TfOGujYL01AWZvdbmuOc7K5u3cpOsH3SePTg
yDshSWVV8EKf0U+sNzVP+2woxJZXgc9I23cuc6i2RRI+Qoe8lvKy18gfi46elBld72dd4mTTwwWa
yu1s1h+VlzONiaaP0XKECsCpj72JLjvoLwu8JKVNcxn3nZcRy5VXIK0CZbHSARHYWwNT/RspnAhx
qgFL2PcWCclILN52ZN5NaXwcQHz6DAS8A5vgr5T7N8+Kh0KTSDeuC3PDuokkfsd1YTy9r0bmGpxs
zkjOP5qNh7Q25YdtB8pcwXmPWIPLrMkG2Lro4sZDGM8SIrXsCQrM15+GdR/XdcIU0FvIjrJ1ovGS
XZaB+FW6ms6P3KPMxN55ZULl1Ztz/WO+m8G8VWkgRP61nOBqTuamiR+MYzyBSdA8qfOl+XERuxVf
jGiu8Bh6shZ7ka0jJlQe/Akm7msOm+PXgPhwxh2DngsuM2z5OoDfMaWkjq/gwSU413rzTewdbvd2
mpE/EE1VEcrxmAC5S4SgAE1cOF3b9NPtVPHTF068NqhNPN4UycXSskLgUC+eLBFzklNp256P/abF
7uijcvNzBWUP+AAjaG9pkSKuIMiFWBR7DSiKlgeishbiMohvgnezPpovWG/qFo+FUFjZzodJxMYi
wOXTDZ9OFfREBwR8lPsBIOJEBoyUoTAqErE5/c9wELoc8tslQc10rOOe3gHudERrqPGJPxLNXrGk
6reRQWefDyJqlY9gI1n7sc7mEfnd/MNXATGGvanh0ohudGIrzz2Aed3lUWRYUgKd2n/cZOAe8sgw
qkSRApboNdt/Fz5F7Rfvjp/3/3dt2Vunt5redYUh0KWpgUq+Q5oImujCPQADpfVs5sCvQeVv/ckI
SA5qmpXrcJtXJqW6hLfQz67NKj37QdqVv8dZZ7lXAmZeOT+pyxVp6tliA60fo0Icm03421u85Oav
QlnxIx/j1AQBNgGarHTeIrZd8FIqQWedebnCnzWT7LjWdmpVyZawpzTPkYb2w5YF7ZnJ/m4GKg+x
NtvpST9q9a+iV87FfdMwjQZ3C0tOxTO0uRV8wlPwRmzW+JkbtTJST6AFdy93kPfigepiZ5a/vjaV
teT+PxIrGJE3z7SByc9TsfbAeBTSETa5dph/YLe8GCxtWKFnwzrHoKWLzwsvsDiU4mzFTseVMzwZ
AxPZZ77Kp+yUXs/4av6rlIcj/R1+1jGRp0cekR7N2Au04TkOyKi13ulmTL+9tvyrrcVKMF//EVbN
aw4DzzuKRMvJZNQtwDPfJVrgxg3J5pKWjq9pIeeqKqfFC/rdW4Wm7ykQhNUIuP+ztSLZanxXgRq2
uFVyDSNuZQVjXdKl+eqk3lba7GktSNEEqEzKtPNDuW1p1YJByNXfj59YLMVHRdfPKbdFO5tibnuk
tRyX+LSZ8nxolEJLNmx76PvKTOHHWmFVMn/fe9QpCGdY42NS6PGEmA4wz/DU40yfqyaxv9k2TKuF
S7xi99Gfe8CrF/0lLMoB1HXZwfj6WF4huebFl/RTmW5R45hgg712quOXM1kMolaBG7ws2vm1MkjO
kxpxpxTcfOJtNmHXhf6nkUwevmfFSRGiPd7XYe+/y5/hd0Tgun13R0/wWuPh7kJTscCuy+Ghm7kU
1WuDhtDK1BNQSkZX+FP0sYv7EQZn7oGk/+M1cPU8I4OWOz+RGSfi/v7J+pI1DFSyBIeys5jGpYkW
nRR/BM+HPYn6BKK4G7c4m/GSRS0WtnrJ0+9PMRu3Ntib0xofrVs7cmFPqIzfKtrd7Q/iV55LXml0
b8Gl6xxm3YfIZ9pMfjG9IH9FyOSaNCeTsRybP42RpDXIEWHwB2lGNK2iTkREGPXGIiHmBCUrgm2w
XWp5yxo+np0iUvkgcUR407fGXUITJqVLjK3IIEf4UK/eWSHkDU0fBQx3w3fi8g7uCBQj7XlVyieC
Wq3A0Gr5dTq1QrnRr7lokHES9NTCjNHg5JOYU+VaiDIFHhNVkrFoSYS7JQnBEZdsCiaTk+5c7Ejx
aGgqtU+JIxAs5h2Cx33oWoXgXoigQNfwUb0fMXNyrFbqcyt3GH2PQi1thSrlkUB3fGdCMJBRuIa1
XqEXOdK6Qu7VhGlFwk0nTnTUKlAhBzk29I0Uz5f3oOjQcjT+Rqd+BMM7f5ji/zHcESk5q9JTWBrv
NtT3iGFus3Szi+Kmn5Vsujseh/m7I9J3mGhb2zW+2uTlcX1KRd/GsMmrwjfo+gAV0S0USm23GYtg
0Pq/nUPLBNTnHk5uYIAY2fnZnpfWoNW0ps4pvps820EGPAssQDsH2l7EDJ5+ZehRWHMHz4E2O9cc
WX1OtMGb0dz+vOu/laFvJ9scm2WyyYZwxom2b+zNNfF/4I3mHDNR1PXWvWza/Khzh9Tt9pMTZkR/
aIzxrExJF6ENEeI//mNewOYiXmw/39B0jlEezRiQ7S8wYm5Tk6Y8FOnRicL+L01St4kwqibj3Ma4
SLDyeHfTOlxdGEBzjLeYMzCFdob47cf+4VmmHiNnTlMXzG6EKJspEJeiCDYss6tt/7hjYlfWs0rn
jGA0RQuocE+IUMyIW5ztA5t3BJf1YSsmoLopdKINJrhF9Ra9TAy0HNmp60nkuElfeZbQtAsp+nlr
6JVfDGrRZQ+rfMnuWnIm+13UkSYC0O3a5TIc5LVtcqnchQ3JgeAfzhGBJekD+dZS6fIqn3Hi4PPx
BRngw5aImVm8TZ/3AKQab+eQsdbQr3TNUSOUpeixRIKaXt1F0DHThDV9NKlx24mYUWR3OiiBo3Fs
VbTi4vGL3JnuSZjVgfX7EsUn8vGtEswZZg1c6LrH7Dzu6Yj3Fq+7hgOcrb6icmTHGdvRB3slXnuw
Fmb2SvZd0LIXq3pLVJ/1F0t1Bo3LZK7qyuy5ozvUTGUVrmm7qmwTu79siIakB957xjvpFbspXpOr
wDEpdT64oHI78YwqkBnIFJFmy0F9ySYrXt3xZw/w4wIcqF4JfX7rysGYJEZr32Gfmt+TR/ZqNYmc
+bsN4YcwIbfhMDxsT9BfzivyEQ1y8vgMo6tvOs1lZnEV/R/cV6lbd/qAiaBPFipNT33dAafY+v+x
HszoriYxToToyB+irVZk9TpCxjuth7m6wOA0PO2xVhLt6CE/yJz5u/cXeD8sRcieacytNwluCWL/
+ptVqdYUP3zO3pWR5ZWMsDBrpkW6vK1hmPPNPkrY4gCutrIE3AtE2q5cr3oVSl5YHBy33VaIPu6w
kEx92CzMrENoAx8xLIbcdPJojyppIhqE4g9ZQrBPRfkHZY836PcD7v5z+xJ8XT4f6bPiOiw2lQRG
ITj6TE/9nJYhe0kTksfcCBJNHCBdFJRCmbhF7uDCSFn0I04RMKK40bNR1U91Rn+IKhGA46NxkLfF
GBfIhAv4U1g4R4IuJ1JZpb8vWSqcKzMPKqHLF59PhJmZoUigTpWXKhu0++dfN3NixlfoH3YOqj+Y
OD/wQUUtEY7oDODj6Z9ZL9u7YTSy2SVYV1xwNn7+2M9BCH2FmyQwjycr+MQJxfBAK95dFXdU9Ta6
xPE8msvkCaA46yEYqpCO7wyM70KvUOKJgCf8KIxw137NbAGcLUErJnezXD0SDURxNffDuAPRfGdZ
5U4UVy3uVPr7uWk/V4bdEQW8c5tFZSowYaW++ihbe7IQBCcs72W2Hkn+yHcSKq4BkWwtBRBMEYog
DHJO/eX9HSPTawU609jYZlG4OKWP8XiWt7mjCKoZJu6lLdhnl318aStsvOJZ/KFGxl6ccpyapVlX
OjMuG7vEWr4UB4cgJ26EuKPBZbsVyp9hRV3BTryGTtoPZWVTUx1WcD/UbSqxdfescUcxB7Pm7BDD
exX/gPTMyoaHlp3VFmQ5icKXmmh5pEupmN+LKKAg0rBlxhFAGr8GtKFMLYOjButChfMatHe2Rx1h
G5UJI4GHf2GXtjcuPAT28xURsEfrDT5IvsLjiLI3SXjdbDSo3c4SXqedE9NSK06vkaI3N2NB13kx
cAh5KNDVxrjJT17iV1AaeK+PIen+lb9Gbt+DZqE7tXQeLccSM6ZTmnC3ISXzuFHPXioMW+yeQ98T
VYAx7x2y2RK7Ux7q2ykNS6uscAthenSG2XQb3fSKg62ZUnB7UOELWhZ0EYA8Zm7U0nljKALvshfD
F3KYRLGjvOOZ1KPsNT3bEk1iw8x1GIy4X/9Dmd8tjKGkWVx0+mxLUxNwkAYs2lzooQzm7gxhy+jy
So7zZNRZjIWzyvAcvZcaRnttbDJzgr4yd1r8TQmybsUxU/dAt9gUH0Si6YV1vAves917z670s8O1
lEU6F6wZz/3+q2+xZjm0qw5smz2OzQB4wHZVoG/lgDA7hAuW4t978otNWlzlV1ElqInjG+FvEmTI
pz8if+HXMXzM0tRp3cOYKxBbD5w+kkCSHoPLCcF/IUP/4zRGYBq0rdloG+XmYFKwTYJV7sPT6MVW
//2GUePplzwWYmtf9hAUwZvH+Vpef+PzxMirLsHcixJoNVKy8eWgN7nMI7t/n3Zf555fvwobyjuD
FGthRvvNEUZBOrr0CHIPnSj63giWhzmYZVRu0vWMNFJFOjEBx1YULOSb7YVtv/7XNubTEVAZv9Zb
4s9TYLw6xPXzEQR9ENbgPcTgh6u21HibbljjTcm9AaVjWTUj0Q1zC/VT0Fw/CW+8QC+e97QY9WjQ
3nz2a3ek+2fjKiqVNaKVnnlfjoOEngK4k3t+VQEqFo60BXa1lRVWe7R7KUOyA4DhmZ7RjLM/VVmB
nfS02aVnvT9wf+5cx3ca9eSi6kSSaPJK2z1m1VELAEfIjJTClFu6PIVUAWEZlEOoc+UWzhmsPoUZ
f55gfSY/5dcUrVmsY2Jj8WsrM27yX2RPn/iQxattqW7zDra5IZ7h5/dGqrACBE/5hi1qAUHCzH6+
DtkJQTPX55TlQbX+CHzSfYXtYvHfiKFX6xvkouB2jVwThm6JlwOEY4pdYEdUq2o25dH3Hc08Uj11
Vd2mS+0QPI1/m++14OnuHHaXZcxXFW3pXmPFubfrN8hytyR8rC000Sy1I2ltfAj8XsTYVlzFbCkZ
vb1vySKOKE+769FgR9KOzRlTaXsMcYbf+kmaCa/RaNQIIBwSnPbR7AIHVUr9qKHq7S47UBhZU6pW
AlxRA1GHd5dpaU5e9CPd+6xKfzXgvho1YEQ5XZ8oTFKz0g9/ELR1+1c3ZkIuxJlvbouGKtEcDRtA
q0EYIjTaIaOy6ybtrZsD6ZOcgr+kzOLlmMhA31tjYvTOpD7JXGbhw3yjO39weu4ljYrNLZOGwg+F
m3FVTMD7n7RdcLV6LjFLlC6EA2BmnGcajkTI7tM+AHyI9GdvowKCavQsOWbpZWPaP+6NhUcO7VyW
lUm73Q904zKpro9J03heZFRNwrd1eHamdVuHRwOZtGAuAuXed60qOxoKVvscCyyTE8iBb8gf/5zf
5hFxxYC1JgEzALW9qtmwKWzR9m6zWTebuW8IWXc5itovuS/DZwfnCa7mksOXkY+Fijc2dT+p4rpH
FzQRTvovV7AX6AofaSUeboNCkHJCWSopOxUXpPE0eyjt7TdYnu7qR6hdw50JTPh1JaqYXIVFfdo3
38Zinj0gzmXxOBKVdlQGOVJpaWSO9UsFZMa3FQIbowhnWqppsnlpSa27kFnDHXKhNMBAWEYReayj
rUWJdyDYtNuPaw0QDjkdCttk0pjSTp3RKGqzwUOdPEMCi6BBcM1vqhw/9Ajc7vuZLIqUcGokpSrf
HfOtY3pltqmqmbsjLUM9mEiIwqovTsuIFeQ9o6lL2Cjf/Xj3I8cRzj9+g3Cn01mMUN9YJKUH7dAk
5R2UEK6SRbAfl3xRySlb3aQhvSNcaoOykW8zNIqYuWFu2+8tmOnGx25hLTa6tBJstt/LVevByjR1
JfWoXxBdzXAOYCCVrSRgGoKQ7FDtfzBRxInHtHN5UoCqUipppYYh23dl83aJnbTLeD20w7KjEBuz
UPAPxriocAqCCdScNzEmWMjDuwmKTOGGJXeYkhHpFXaufLd1FG69ONcpIJkFstPjkuFp+o2SQ3UT
dSB7vYZChWE6cvLAJVHFSF1sunsJrui8zr4qixRfT0x0nOw93C/dvsajXWst+efkdnKrDy6Dw1VD
xKC03sgg3eLafh7York1UTl3FTwxUTC+8mTVciQ+yYJwhArA01JE8Pt5zH981bX20DJYSh7UO+qc
4GpSbMDbxcy5dqHNIHeq2r2pqf8raq5DdfBiwJtcOTrCkGile9c6OiieNWKOMr/sO/+ZiEkdP5nQ
dOQpCAeTyGshhG7MyTTi19gPce5Cy36JpUaQqm6/uXakUjsL+OPbRaH/ZAyL7ueoDslBTFiJLnQf
rGPtkYQ3NyG1dNMh+nB2Ynr10yvn7Z7KKCAa7sEeK0x/1GM+3G3FBd6b/HM4MN4DlE7tjyWV8Y5b
6mzmd/Fi80r/YtWtxedvIw118E40Zf/r1HuTntpmhjP+8KEVT9YCFmOxco+6BfbgOl7GuT0QRJkt
iauwEgvLART2mYkWlP5Pnd364SksLh7EMX1wbuQkwfueXIfQlS3ysI0woslXoTlMLfzGz5qT5PTw
y7yK41WSkgMaOZc+vASSEpx7DkAFWAPBd+Vdfn4fwXatuVr/c6PAxJd4VPNqWWgqelLyGQbjjhEc
A4sxrvxuyhszICIoHiT+kd1rncr50tggoRHns4/2Xf/lbv2B+ZJSBA7Wa+qbDZ41RllTU+swS3VQ
B5GdK+ykTaVeD3r7LZEXwl3EsjjkkXMwaAgYh2hX7GUxPT7IdFk0NKks0JxAokyemQrOyA6YR/Ql
P8pJpf7YQQKDZmV1YDEKpDFLJakfj7gAcSxIRPLrBDsWOx8hs19PKtSxX3VpeA6z+7fIeFvoE1u7
opbHbhxMBtIwzXR+cJ/906cID+IeUr5AqvwzfTSdefZiKy3n/xb1PRONvxczcLFgATHe+niEiWFD
KfC7VI8LmQwWdX2xxIuzwawC26V0r/ifWU0R+ndoSDQLDk869YhbKxVaSy01BQ94oMRbuXGrgQAP
+Mjp0L/kOrAi/NjX+Ckr9UA09u15d7PQEF7QX1+IaDETrHy2CZSyO+n3qVHsYJ1rmSScQu86yMgR
PLWnxREvtaC9+pV8746dfzTliCVjb4v87yUb0bAxg9syRIC6T8z7XRXLNe/63MGXaxHYxYmUz4bS
RmBvCq8UAYTu4hH5umUjectDn1Y/CtwyNClUB8ler5Wt9HmivP3NlgoulHy4fRevwW6Afku/FuMG
lv1Nxrtyknavo4uUXO1o6yYvSlVF4tz10Lscq/X1K+/6Y/nW8j6/LlvjxAj5mF11+Kjaa4W8vh/r
97beZxtm33X5l1DLOF+LQkzWORci2PNLPysLX1BWOvNdA5BcYx4D+IybMAMdDD2jVXN/suVET9mT
lqf7RIfCpTvU1UP8u4QGUcgSGbJyaIxpBf5XXs7q6B1PJDnuN6TN2lB68gQG8Nv/AyMu4Weq3dOe
tWY6a39Htd3HMQXKtnQubtgg1ie4Nfx9fiVXD17fKh+vUv0AnHWDZnlP0W0p00kHnrku6SKoitmp
X2AIlso0Y3uiR6gxtuvYsvsFosq6ezaKAdmCWtEaWO35Jl1Jnic+3WNqSOxzLJf1roIh3aktMr15
CIjJn1Ge05mYhL3TTVaiox1PTP0EPTQgOxcdZr8wA4sAZtrVCvT7lsm8ep53r7uPq0flEr0JNt9Z
tYRCc4sL9/csM6f1xHRpSQyvQQ+ETG5Yn7p4HNJEe4+mM7zzrRpxuEdxiK2QYRiJl65AuValz4ws
Sd59NbQlKLc9fHUKy7VV7RCxFro4okfEwketuND/s977iOmwRH3klV/r+BqRn9Wq4CSYBRUG10t1
NzRmH7+fnLn5DjJsiFwHlHbvfw78OWyLVFD00vcAfduhgBQoHEJ/HHhLZW39n2fp2dIApl+n49rq
e+lF8v0+SzSmSCuGNVdRaR++SYW5MZ2PlOJ3Zbs5UslzdnX19c0mStePyn3jW1JsEheATptRn10l
y9AJoNzEd0KH+TYGfBzI9u1CpmOwdk0pJ9zNJ18FYiBQAuAy5W8oYX/RJwyngd79wxFx15Y++eWs
/Z+diWCCzZrPHNQxEOKhwCoVe+AK6GlQeWclWZWcdqBo5PLZMUoWI2fPOFGfs8fwgM3xlT6CqJ7Y
LSpW6QE873xMZyi/W9xVwjaT9H25P81X3s4d/ugGm/l92vc5BR1yPdgCEmG563vwPGDHSmEEntWL
EwHsNwQJGheatzGYT1cFMWyq3Usbqxl0xLcvWpy+Pi6B5gfpviE3rulytkgtJdNFC+FUyjjvC03M
TCCOMSrexpFEO4G9KoJrACHfJG33l1xVrnOuIF/kVNjporW8xDoEvvUdFvKlQ9+qGlP+QyXhSFD4
j10D59ZGAbZsCXDPpGdwbc3irRvCRvpMsqzI37SlLC+dKtHawHkhtfQuyCXxDA1t3mMXw9kca1J2
8vQUIHTUwLFIyWqYVr9Q9dwfw412GgmTcgzpoyHHrsVDw0o+ohdj9Lbosh+ufN5ZczDMAbKEV6k/
yVkgrxL7rIPV3UCgns6+Zah5rxmBrYFAuHXLOys81RFud7FgyjEqlmmLfnHVLrUhEDJ0DxeXSnor
ApghCSdglTUNFZAtqROfOvx09jbA5PfpiKWCxG9ftpKNWqPDk5oBrCw69jca2IRfmGomZdUKcLeH
KdGfciOT0e8Gijf51JLBNNph1xo5W2uNdvEjlQxvO5U/5exLaTmlCTdzuVdOyYOli6lMViRHVQ/T
ehAoxPGoGOi1CITeQ8HDk6yfOw9mwM7H8jawAtR0cYFBYqNHWCsSGNYf4PNkTQ7PbpweBJeboU3F
J4wL51kmJ+KsA+1lm4kEhZSCezMoTBCP11yKHnDpAY1sWztojlgceML2h5+so1H44/yFcmUNRBI/
jK8aKeldL8SholqQS0NIOK74BuEjCjAdnCDCkq8BOO2RhkXaMGGbY1+pFUMwoq/yFgSlrRjnqN6Y
4jF5VvXMgl2QKpXEf5OABbJahs+hoA0Yt9HB7ImRiKRmCQfavnSnNigEMTUExleYyERtG7BfTWW4
aVg8v16EC0XVncN/H+L3R1pk72Ibg/ISF4uPJTM36MeCHNjBxRwbX0BDZB+WBtmXDIxmE7QgubYI
Ts0sVLhan4K0OFN9livG1xuVzArSSgL1lAntGXRq1TFjicTIxoNPGITxMNkm5qXHHaM+EJ2ALScF
1vmlTcviLPABc+Z07Qd1cbs2396pYDbyMuw/NKvXE7bF54kLQiQSqHOjXz4izRXplv1cdYFKmT/Z
75QKEV/C5MpYS3HmcNtH0FqBcNrF0iCMB365dnEEIPj9No3tI/GeQ7+lQOg1Fawl7xOmqwV4enbj
cWm9aJ1zU16zYjyXlMKJIs35dMQPvAnAdJP/Sh8LkgWGNsNa00qXZVLgboxOf1BifQhsnJQieODU
3MMdITCY/xjzGnB6d99l/dTl+Fd3I3nLk10yq4axpsdcQlx49PCTI2rmgvi27Rl1+nixtTRvCmCO
NAgnyyDyBNfhvlpZyzHewdd897Ald30MkAbKQZtYHAz5lgezZUzGZxqyOkX4p93wwNAtwWCkx9eO
Ms+8HqpHVabC3O5L80KUjcv1hYy32ffKi8obLkj9wkCQkCpR6j2YuGuoYXl1j08etvX7x8jjzQ1D
RosONacxM0tuXSIw02YE1+obHzXUw50ZxBbNBg7TsoYKe3GFMzZgmneFxVVYP6dQf3g/xCB2o2Pj
z9jgoqkmmvSQmcPfa6HaAMDILjTmU632+seyf4AWCT8BqmNMcueVkzRCvmaxpE4e7hTINgsJm79b
vAO+wcellou7HRdgolHM7loxq07ZBzIv2rPhFBt+z7472BnxKwrPdoXTePHdLu0u6MFAQxr7cOp0
b4D7o7gkW9C6vtJIbOJsu8edUNGS4Kza+DHA8Kt8hFPs9AbbtdGfiS4VQmV/FD7TzUUSkdxPFgNS
GOiFCJRo/dwVx4GdQennp/Y3bBlokDeFCr7CE43cArI+i/cDqS4h17qNSVCQw63MTvncsjVHxNI3
s6ylwjKPepMDgmMio31xUV3KzYjzIDI6ziqsfac=
`pragma protect end_protected
