// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:21:34 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
omRSI81e5FKbdN5ogWJQC21X270VfqzHsoeeCYgNnB2mqIl9eA6Tekkqf294UYlP
qxnFW+0bhszp4mc4tEIvurVMlMXBWgQXtcMS1JTRQMJ5vUQ1l0vQI97rl5fiNDfT
UfUFlLRdXEXf+bCx4E8o5r+r0++TEw1X/c8Ve14dxIw=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48368)
Xo6DjACws/6xfp7Cbw/LUmxjuG8MKq6Fwb4i7/JlU8yz+Y8A5/JBq0UZURZo6JTA
gLbTJOfguciUcXp7Uh1XGyFa66JdoVPyk6vTza/kE3fuPi4xrGWGVS2iVphTBqx/
y5loHTBznMxm30MqUSuoJ70bfDh/C+tcF/3FpXVUZIQbYSZLjvk07NvxwRaAe2s0
WYzEbIK4+bCZMn09KaUxoSmsJQ1zs3gh8E2TxjsPe7US65atHTtJOiS1i1TFpYE/
P/RF+qFO8TgprCmEExg/yCmjcY3DdrJaw2qb9pfWm9ipvFfeELhLUchpCN0HGYG0
V2xNlmz3hBJh0svHQ1Qto+eB+Oegg0w70jRftGBGxKwDGJFdr0wAbJGRK2payEg7
Xi6HX/FQoRgHkK0JSQoZpEpO55fTciuaJZR3ieY2C0cEsb9xu/Kl4qaO914Ydo1o
T8f/kZfZ3JrpXnfGElfbhnq5k14FRANEitPchj/hWlNuO0cKGh2oxhMDSHzSfotA
GSR8wJxm8pfEDbJ9/HtM+enJyqLd+YhD4VcwbmR5O9Azu8NDXtHHdMEbmqHV8Y2r
M3JW3hNRWPqLYgdlYOTO1V7GXuOFyN6qm7wRQAixFjwblYOVhDX8+w2fY3JgE27u
X6d39zAmVHraAIroId5+2RfyRAnHlkrPux4VmLQdpfyPJF0lUQDmCeqClycCEOIl
KK2NBVgS316J/qr/sLeEg3b8dHY11tztG7z8EuEoIU9k0BhZaW/k+QvgDuDj1/w7
FeRvLeEMfGQsFOLejhqp6fiMwCwpu5o/AjeTD9LbHFQe7zoZtqF5EZO4gGMJo6Xy
JMMHYM5QzAZI4FEfLQoeqq0wPp9bzetwUy2+tjHWh7CjgZoeF2ZJBUQCkRdfr8Py
0/NRMEjPtID52BEV+xKhSDiFnge4mjwpZ/uOUZWvcQn7XPQF0oGtiUqO7YIO16l0
FSf6LB/639Be6lGAvHAIqmeckPM0jmKXfpFgo9fllE9P3lFTdvvrDwg2r61JkBtG
xFElmMa5/XnJbpdGyrqeukc8gWE7q/ef+ume6zQP/xSj5tbtIrmTbbZrlk/5chMy
isR8DGHZdM00f7OqXJbEAxf7JBXzrEqPlhmXqP6VSZDlqdbjItF2SoFYW4KzEx89
mUIPaobP/brT0N+l/6zZWDywsriTPm0TZQvxI2/gRPqEHCh04jofM8xDEhfr/6te
K7oN75AkRMnE0P5PvYLTB2xuMIJ9AF9zI85+63hfGjzV3IIBqEWHRqpaSbCaUm11
8FPDo+XlxJJzakPwz+UKYfc7gZ4S0JbzpniCxdmgUHsOizXp8s3yyoCP0YrFAGn1
y9QZYI2Kkn6r0cSdxHP4l+gsBVGPtakAOnR9Z1z1mzstA3PhWVD17+6gPkRmc8iX
pbCnIHmkZzqFYWTjIT54FSE6nDWIx3F+d/F6qdwGY8Xkp5/1G9WgkRkPwrnQB5BL
JBYyWETN1fX8fAWIxlMVUf/oFNlWH5lwnEKQioNS8mdUElgN6R6dpL4RuaywPHZ9
L4yQZ+3SDDc5PIf6pj3VoaJtq2LJgYtvp330Ga5N0f9RohoA7/9Ue1hZa5XAUcEC
fbaBtEG0/8BndhfLfPU+SxsdVY1xkgzNptwAvTyXhyFwRb7SH1TrMvTc1fpvcVk3
V4bPT+ubd6yF7y7ZzIJlrXglTSgi9cNFFAmO/LVqWwXE+nuz3qo9WMNBdS0DQXlj
3OdVhVsheZvszSUArSOGXgT6yob+qpmTJ10FckIw+nw7P9TrEGDPvrSLtWwHelF2
Kkah5Qk+puR8HTnrsHbE1fFe7JVGdtgp+7xgCbeH50MAxlxZP9lGVTQGHhhA8+uA
DjJiODT1pg0R2rOQ8MC5TUCeA6PjGlTTfmjsSsulBsjJZWs/wJBOwN9kui70+RTa
xINQWOIHdigiu/2cUjezQl5mEFb0g0DXnZZ7ulsO5yp1SIceY8mYg10Ug60ptlbA
OBSIoXJubJUrlh0F3avdD1gB6QkXoNkJXxclgSGilAL3wkvFJ/kb3/ELthICThVi
6Zc9hWLJR6Ch7dAsGf1LC3ToSC0k++wy+R6Rf11zVPXXT8vgUNZltlV9DItsMHJL
NCDtUDOeIscXlh7cgRHve0yXpAqLprylJCuWfdQYKHiMtde8gTuvpPFkiNPH3gyp
VI7WSKk3TNguMt+twWrUKIB2PRqfGbVQxWMWKbfRK0ITSmH0kySj9RkLgn5zPdtI
n/cU69PunIMLOTzKjcw2QPKOf7XtoEu4SuPzcWfsifHVKYN1anZvzYna3NUgqBg+
mr4HmpkxV2b9pOL5egtZgshyju8dAgG/6KSFWOeo9hbXRH+3N1JbCz6RKJPOlsHh
tWrm/3tNO9puztmzJm5sXf3s2rLwsm3gU6EJBBoHdj0YCFeEr693+6gbz/gifieE
qo+bXSNWogj7RxPF3f/Av+9Qye3va4VCAhM2jG8mJFNF0OBbiTodLASJUKra7OpP
VE/0XWHQfCXBWkV+3W4DQY1YcwMUI3NPDVnNpuwHYKZe3RIRXh05qBKvWzMRrQ6d
UidIrpSsHo8U4UgR96whd8L/cocIq/Nor6SxJobXsTq9LeCA9IiQTLYdotwwoCBf
3AGfADCLln3NIjg1HkRa12nSr30ZZrBR/vBf5ugkzZ+C5+ncJkx1pBH6T24WEyzu
K9vQRdfsNwZBvpqVc2A0m470QemvZ/2HgVbCBEbORFc2IcUpDUFShRckwVBssHr3
ic/oBWfnR8aHOAqIshUKOO+gaX8USDM/Y+r/EHLonBeFsy9YIXK6DMyYeVHnOebF
iDJXfYwxotjGGLXl4b7cTCzRBC33aDxpcWVl7xwY0hEkL3kilEv4kk2uN+e2f9tz
SM22/Nr6BL1uq7YN63naVQokxVqsOURsWVjm3jNLwFPXLLKsrd7Bk34GC6qE0ETW
7C89Y91M3vBIR2vhd/HW5ODsRkgWoNwWgml7n3ZU3EvUlONX8DWSCvod7mKGtGi3
KkSpHsWpG24etvsVC5o5PR5qiEwQDNBNAbSk+tbgw9AcIHVb9djj6vAF1CIxp6R3
PlyhnPoNIEUjfPc7r08RL3P5rO9XWyws0eyJCxU1hGmtwU97k99XEZpfanLZXyhw
Hb7WZqiVdSrTsL0kunNr3k+ZaRXpvq3ENnS0hcGaJrYnhks/prR4uNIJuoYO78vC
yT9vhLyTNY8mf2zdy+OE1CFFJy+F2faNY+wx3VmpH3XGt4hHlpUPq3ozZt9kjSCv
/fhnug9EobHfIwAxtyA97KQxA1D/ccTVZwjj3nBcmzmKawZpScVr7zOqme965nFD
7is/W/sdVYdtzfi3oF/FAKWcZ03mglz2Lt9VWJd6ujgwl0C8bQrkEn37b6op/Twn
qnfSuKOmdHsEz++rdjtMj41mKSVwd5ddWb7BBqLA7oICZ/c0UWFek4pTi6EMKkZ6
6gyMvT+XfYQmmK5XLr1EIYSQNEjdZfI2G2NG52bXqJA/pA5kQ+JVIDSQy4IO6ewW
FT98gvd84VOfEYUKQtCprZjR4N/lcMeJST96zvo22C97AXv7uISueiYvQdbyCj58
yBfR7VZS4CSAmFssY5GVdm6Tfv96uj4NsZ2v01TJmcNKPiu7CvWcglDjxUWdE4JH
csIo/Ad9PuigLCP8N/RDIpv7Vlb2nBqwz8wtUoy2ZPZUza/JX2SNnSljkbdww4CL
L/UYNDap3galOu7ckyuOcqj01aLqsdeJW8aCV49lUoMlzb+uVGOE1xX4Y2yLr9Fa
Yh8goKaCRCsJBhMa6LZrtchU00Dbric4N88tA9ovhvAgHWrFlUix1I490NOOPTzy
e78MZk+5Yj3E65YZ9+tu823OSqM/OZPp6/nrmbzsAiElsF0VaWs6gALA5mSkacUz
45quXJY3gtGmu8xRqYVjhzSLIb6Yo8RB66CfFQ/hCIR4VoqSSIA350bVJljMe6ct
rY+wEx2OCVP+wMqAq2etBv/Yz2kn6GubGvykrS+lyeBhew4APNUbIfqVL4Ji9/gj
m9x0PrxnnO/sCd/VPLfNX/ljvkOBc0wxqQOcffanTGCo3q46T4VARREHtzzkkFQm
vR9nZlzT2MVTSPVrcnb2aPqs2WGJ3CkmL6X/zXuE00FwXRO4gHw0Ev9wiaPGRKtw
+w0WBnfg2zV4yy64LRkoIOXEdEAsmbSt2/pVnH0tkjckms6/oxHBU0tvy/Dvg/4R
TNrvV+IoIqSJub7X/VI8jEi+wZRrGUl7uznRMlrYMtEhAxEr+nCDkWlQYuoJVd98
OaMYxBcvd/3nWWUFW7zJkDUKS/Qef5lhwzGB7PFveVtEzabRYvaL/aWN3G6QlZ2o
dL12gwpmTk7+pChAIKDG/W3E6cczFwsakD7z6a/z2ESBvMmFDcYEnEsCOlct0pHn
O2Ss8fydUTX+bxEECjh+e4unNb6hFLGnBdYr33MG+CSYt/oULl574uNQjqB5kXFd
3I6nY3JorawUaBamuIo5fZ6nkRIojPurXxyc18QZd3u2ovRYl2Xgqm6rbC/PwvUi
ZQUUvLqrYXQiOZB+UleNsiy6k+4wJY2Iro3cHBpv6yz6P9A6UjlKV8DWrdQqQcDQ
v3UZ7zw5XGuId1tx2vBATPthksK8zZL3H84yFMdwunx3TMN2Qgy5J2+y4/mYYxlZ
5A+5ufVaFYKj7dprPJhu4KPNJpULc064DWCySYbfpDn7b2Zxwkc3aZJvEtSDdF49
PgfCNkb/WGWnlF9MEnFsObCzSopk4LBP3zbzojRut1kUWMrKdSWaBjVw7sPsq4Jx
4CG9rUpXJ4jw7cau47TQlS56kAbqasrS9wFioNF6MI6tD93RcjT5lIhsx67rlqSz
qvXQQ2yaovjUk8OH3I9WiTlrxcXPBCxZHXgXpe8cODUOZnu+0lwYWqgfUMOR8cTG
kUtMNLu+LBBuesRpJD2jQf1XzBMzkWmRe73OGeeRfhD2kh4f+0cXQJ6kHc11WLr8
8WfSsJGPO5Ts0hCFS0PE1YAIUgiKi/27qS44QhWI47FBB70fwe5ctxOk6eSCF/KR
I8nJxM4ZztF2daQDHVYwvSoR/V0dyzjUBhL7q479657daRJovwiJvK8tJnO2De4X
jWdVwueadEZ61dBFx/3G8WF28fCUqzHJs+FV50nGVD8cqtKQ+zxH7TSY9MLeDxHo
AofsdXKMWksgrQU7TsixMad5mLfOZTFqL583BLu8r3diHjBJR2O77ryM/kgEgiPL
73qABekKZiNfyXTC2cfTJDaSNzoZDJdY1Ach067u52J2uSy0AiqMvx1Rzj204zRR
PdKhkAwIGxHHErDep/P7r41FSV4N3ZCdSyvE1uNbNL1SbcDuj2nQdF7PpXWK/qDc
lMXMA2Z1WyvOdjiZzATitmcVx2ojDU3z+lTjvV+6rVMCnoemONc1vJJKkG5Mouqw
PSO53zHOSWYIosW72I5+D8fUmCXmerKJVR5lGMs7FllKnqu272bqKGdfNRiebF/U
BGr++1PQP92rp9SkbBkGiZC++wTMkFi3BnSS8uRLUWyKw+bi2TlF1eyDNMm2+2dl
xxjPlY3jXBw896MjlaB/HPa9OqjQzRJ1dlcJZ4mogDm8dYAQ+qMgpwAuyqmClRtM
KzS0Ylg9svOk0D0QZ0gDJBu2vOIT1OhPkvLckw912iWdS/ehiJ2JgYCXSfqhwzUy
olif7qcijKtoJNS1EVBMRlJoF7uPCpjn6N+DKgoXcBBtOrE4ZhILGmClxBcqMFsP
SpKHe7gNTyEuMofTpIoII2f0r8aoBO0h2yf8PkHnaniGCXRYx6op3buyRy9LZAnM
uiIWH5g9u6lAXn1yfhSZlFeJWGpnlDxSuRhxPcaeRID0pomVciYrq01XcEFZVHdg
nhnfiVyadRf0p1di35EyzL8jQfNdJsirhYfE8EpU+SfS7rEG+rsNPIO6pXwoBt2f
nMOet9xEOlOqusaR3h79nynKOUV1FPa4lRO5edosn7eAoJubHElZIoZEfxkDQYhb
ZQ/GkRTpCnEyk79iA8mVcIGIl4g6/5SjN7rwD9v34ogA6iMlYBfEpjfizG4cOvfN
7v6Y6N+ip7NSod2R3ENbsccrZCsgTh18zKrgGmVEn9DPKgB/zQMaSQJwcq6WyhcB
vxRcEYhmLLZow5k3iDEA9U80+bJldUKUm9k78J/jBeyv6itfk/rsdAiMnqAdN4a5
s/S1y8THd+yFHJlH4U6Haw4qmiaxoxC9OMqz2YKHnLGAeU+qd8MFKjEh5yeHsEgp
EnxOPWFJv6CyeG2fJY8JDiDMRmhc8+3WX8J5NsE/5KokguPaqM6BbyfeQBpppbL4
A9g6864ksYkThY3v3qLkpMDVCBIsGVkHnZ86ib84cFM/TGITHBlqn0SGLdqhtPXP
XTyirR0gKjQf8+BPtPGJ+pXhQpJU1gQkgXxY2U5m+wTAmQV1PbRrXcL/5dlZwlL+
PdgsL49CfUTEvrNtkU5G4GUrlNXxOdI77qMuFBugpXYBh9pzShNS6J92dxb0fL5n
9WpvSaXu5U3jjJSVGn6ZkpMdNuk1Q3aRQp5gYBVgPj/gtOTUM0oocM9m06LaCw59
2bHhDIOTFK981pgZPrekAZsfFx1zeTxZBYknUnmx6EkRtfGkJ/Pa0DinPvN2RZm0
Q1gvC+lw7umhV7b9SwuvS/xB41hEUt0Ym4ytu/dwWLfGNPWeB35psiAsneEAWl8D
s6yyxjxmhHUAT2kqojSV4Tdm9Yu3lZsvlidAiRRQsJp2p8MnwOYbN+Jm5vtmFO6B
yNIQrMV+728QGRkA2mIYgnoz+J0yDFmjBwS1SHpA27Sit4/lp6YjAsa4roY2RhPS
binIXY6w016gBq+IRC36LUz1yiKqdZ00HNDPKFTVROBrjpYstahwtjhcv0Zoz3ky
/fr/0XZ4I8YK0C1os5dsN+ly6D5IovKPBoj49uwHXDp5zsSFplTX/fjc1WcVufsB
QdFQdO8T8mgPtECcN8fxeYmrHx2pO7FsKetMzbni3TUBd7xDPNW0ikXXEiELXbqT
ouYg4Zg1azVeNU+jCDQJXJPpfwtlMqaDTNt+RtOOOIog/ytIWygkCp+4wWXOox6I
irX66DGjfHXq5kCVDx6fHAUh4TztsY37C9xFpN/ZroUvBPir2pCJOWPo8VA5fOfJ
pzrt80r8AZzhzaJBAFYz9x8PM8NHimoHuexxfFI3VFslL5ruA7HbIPme3sTsxwJe
ko5XNeJxDwqglcmIiOR7B4camLmR4u0YlLLklvWlxXTWTWms2EK3flU3QXhFRSu8
ddXukZ15KoCEC+3VaXZMnh5iH7RKbOLX3Esu06j2AgN601dzmPm3g2JvbPS6mkuX
TOdfXTFSU7FhaOjRcoHG/e76OGTvahEsDvCEpSom00Ks0GSLGro00rvKkyfFOlJW
/UFZ9gpyRLF7nQA/iYtviUrcIF56p+or6reQzxWRYC8FaJJxzVNZ2odDtE07YOOy
8zzK/8wrDeZ1xwhqZNiBGPXQa4mXrfLyIA2PsKOU0xQJQt1LmZZNWwr4g3N6mo+D
mg6McgAnduM91Bhe0vTg+NJazF76r5i0KzfgbmOdhZfZfb0uqFc3DdMpF/YlYzxa
MGCeh0dMmQCSfkaes6Fni//CndibIrLuJszfKQZzzvcFG+wjcvu3zt6jnF3w7G31
VCJzJw7jOWY5hh6YeN5xW18kP9YArLH365zKGdBsYgZW08EZexQHOQ7Aj2x/dHSf
J9b1BeHEUgQ3d/OR6ONfO4NcdzJCvUVgjbqR2j0g+wR97Mtxbx3AroNXf3OgPrZd
ZiXj+MRPbIV05tEDBoO/PcaCCAnRs8ZiQZy1E+RL2V0US6hOoYtaOst4aEXJEpuK
w1U3j7O2rjGzlpt0N+tQg3AGf2Z/XcVPCmPYJTdcT4gn0TwVNgSH66S+pMDYAwaO
enaYlsjU0efgTThF+OHYVLlv9QpOzMaacUJnLWTtsx3bG1KlsO3hCBppLH7JTDkj
TDYBsb5vCaQ16p/TUUSPNDatTVRQkWW7pWok/SzUfU/LS198mwhan8m2RTDWy+zK
nbK+z2blwUY1VV2Jb5ATd7zXrpvW10AJvGtvukkUNpihvYdWdVJs4lvJdYbru3gr
DpzHYZmdfKDkle5QiLTBMe5rTCkpVhZJwfBvL4WqOoGAHGLfFascdbl1wnAdwN8U
qyNciXcvHyALPh1/n3QMUNEjNNknxxWs6FbZXIAdOCJ0KeQxiP8FLfqO1/y+S4fC
kG5CXhn2A3YIQHke2zz/m/DkaATPlj2IpakTZxb9u2qbX3i49RkLjqJyVUEbdE+Y
kqceLgrxEPp40mC/GwXOCtk2bllSveQ6Aj5E1kXKpK3J4jfmm7TrKHl17pgRc5nS
g4SuL9pAMPAbW8f6w+zvBdV1WBHSlO5zhTBceD98Kevlw/IsODU81ZK1jT988tn5
CtqePDY7Lm8KB9cslUhrlWwYokFaula75t3Z9ZOPCBBldciHquSUKQZ4TqRuFvGI
m9OK6gMBiyEBCMR0UWj8dTR89sdCsNrqomyMlplCHmhTbFLQ45hqhEEKrhDm/Km5
OWFGXq55ohK3T/d5LCFFU6x3Ajamfkbh/lFy9/YxhKMZrejtvIIIjn19yG79RWqg
GFdsDGIbRFUXCzk7zdJLJXVP/Udfz2n5II9GqjQmx0AQ9AH2q/jSGKByKp+PgJEj
/7FwW5Lus2nVGomco87MrNxi3pcqbP2UlASrvvf6A9bKDKoB+eB85S9iwnKTloQc
nq22IlJJXBUlrYuPNyrUnSd186oVY+19LzNzY8op5RUyFz+WXMm9Y9WSepD3QbRm
QSPb/UhH8SJlzYVZN4AVqEEoO4m8jp+RfHxgXoDl5/SvHexXKvq3y/xAiHEb71qg
hLFPkfxqLOlfy77ih/aV4Up3jgxgJq59Pcvj2kata+Jg7mU/0A53iaieswOKww/3
XYgBMDYbNdywoEiRv3aKceJtr1xAc18UHC8nqh1rPcK1LfBeN5ikzhYZS54+PxBi
wcaU1HnaVjHfKUVTvfZInS2UYS6HlpzKfPSRHrRAYWVWCx/UpHt8POiI/8ScJsH7
0isE9atgKtykmdGN6yZebes+H6H4veG5eOimsttthZ1QTWvvLja2fngATXAFDD0f
dJwEMBEE/I8tsczxLzxAuFrRbqyx1AQsREi2jARCvLjDPVKQ7xaoAftioq1/odHy
HwwLvb4gCfmwHVK0m4znqxG4Gs36sIJiKhFDwZV5a92UoQ4KaUWG5IvUyqZh3YqQ
SrV5b9YC4hck82UuGe9+HJJ/u4POvbDhXo6OLamXXLyyyF2aRM2GRnmg45oPazgB
VfH+CWbUmw5DM6vsK4eYyuK4WPw++IEfHvz1PeT9O73iJWAgyqGsFfPcJH2/Ghet
Or3C5iPENe4jFtagH/aLoO7xDJoqr3lV1EAnLJPn0y57yD63hvi4kmpPseZfw2+e
VIW96A9wUOdTYuCWt2R4A4xvKtbLJxeg0+3V8hYnHQLxG+n9glFMgTTG2x7a6t9y
IAIe6GXX8ELz82P0bNcg+EhX9G5t3U/WjntVP+HENQSxysc72G3Qr4rZq1ilqOP9
KK7aw7wATyzV2bLqpAlUCGNmrOV62vxFI9EA5ijv0KmSe8ZT6KwF/oMz0op/tAk+
m42dMOhePM9zAp3SDYhPs94v96qZ4LdD+IyuiGt9SoMUzRi2YRfFpaax5XM/FQWt
ZithDj8G6LLHFi8ii/T0JSt0dOh2PgnvUe1/er6nCQHMplqRuJVc2A+MW82n4xb1
Egnyw97EhbVsCj4CrSLro+hZvpbhTVyJUmTzdKfYNkJ4qy5eoaPmEmnce9+echl6
tAXnhqyuwqqfLtbs99AUejH8KG09Jjbtu7rU6T173UUgcnZRR/Vent2kkP80nVk7
uX3fLomeV45ieYakHIafjCTRc5U0YwmZhDeW3wb9/+Dl6D1BlQsRx5G3CPQW+LaX
/kMIVFJmhb1cPN4IatyT5BoKsH0SJGaRIyjOvva7ZYMN+2n3VT06GkcdlbOu6WVR
b7g9aPOO016iho++I7aRoufcweoQYqMdFVbOy7nuKCF+JNoCBpcAnfV5FwmauTM7
NrFAnZm69GHMPlFzydePTOSgjDFU05gfv18tBkccqhSTv0C1MJMCVVTAymnvsQEs
5QuNmEnQYTGwFPJoJqDJX1DQufs2IMHxCayzxWZTfriuJeILNTbHgZ0xQwg7e5bN
MRCXi9tdqN6Xikp0SBKtrUEMSEh01d5BptNfces5uouGVum1P455LYERgdYDaaUq
K/dw/H9oQeEhtAMGV/RERceKn9vGiANv/02+XnMf1E3eMIpF/b3dR0lIN8aS1Fpm
jS86lkBKud1/N/gBKNFvyKoz/OunrVjYAx8ce+7+0gUEXvTAdVk0ISvMdN2mLgJg
wTr/FA0S+AYzZVkAglUroM3yXogQhInqVlvH4ryeJBpVSTp/7yNk9oX/t1nfDa5y
8JFJfu/AURMXKOsku/oIte9/dXLuy9HHB8QCbb08pnVJ+NJbPMmxfI7x/MfoH+qu
kvEpq26t7ev87zBI9A5FmM4+yyzXmTc+IK/r/9w9rhF/xIHVWLuUjdRzUXBTS3lm
EeF+k8JkHQZ1lqLMq+HnpE6xpmzznc6nALxOghs7hCidz8JhlHBLF/8+xRXydHod
OUwTdNUZc5Ha1B7EO1N6FIBlmUG0nnnepLkSfqVVdRk1hj/LBJbcqnwlyCYDJ1FY
drKozlUAUe7YEMKXEBxjJD+icIrUl3pNnUMeLewatrzYBBwzKXJblZz8B5Se8jXN
oh3pnFoL4YCYiFnZCrEEvt2YPb7l2v5Irr42RZsGdcQf0Y+wBEiZLcg1Tpnh40Kj
AOGpmUw8wNBXJSP5glfCIsPKGytdhtp78zS2jfLt2KQ7kb1C6MnjYBlyxF+RxLrm
2ndpmg3UvNMfmqizeOx1orwG7UmPKY6bQy4rMWat0gVEniQ1lITiJNMNepjXqjbl
DV8HD7zYykuhQFJLr0sBhEcaQNBH/kIoL7XGuegv6lCishb/xmrzB/dQg6C4r9yn
m2h0KAvE/qT8NOMuHh/GaiB3ftjR4hudoGcdj2yM4fwALxG1hpid/6OF3muzID6s
oYYVBnsJ9B5urrRoQ332O1fPBoQ5FAvL5i3c1/z/fvQLOLtp3TlRRgoUu2xEsLx5
s4QpiJNfzSmLoxuyRqneQyJ89yXXrH+EFIDozV8zNidG4RqtdpKuRxOOyqBWLF7X
dLQP5XXc8rlh5PiJYFbWEYuNt3rlU30Xw3f2IES70Rtu2Jr6mYy2wRsegvv0PCIO
BWGE3YsMxXq8juHr+4K91ewlvyRYlhfSHBllGii8K0dEVArKeIyC+Hfd8M4LmrFb
Td9z+qFnBOdylgdhJubCyib0qGT287FfZEK80iSR2ZajfZm3lwa7xjWveQLaCfiv
aMpI/vWg28OKzJBSGSVcP5XaPE5l+YjSlwYi90k8524dX9dMCN8+IWoC+E4+LriV
QV7ZH8O4QDBaE2aIdMsOD9Y8MYRSLXYUh4J9zayySa95Xz+zpq1kDpIGNTpG5J3l
gqtuS7nIIs5CwVHaT9e8L4WBSXfuiYE5LWaPB3WejI5XfYCvrKtRrktuo8U5RIGT
xATsJhjTzvPx+DTVgLs73QCP5yKQ9BuKbSCvd3uDmHCCbjFHIevGnpM74yHODBtc
dGb0L3L1w+mVc+/Q0sf6Jc5bOsxDGrCPLdsmMjAhlwEmBUTLwHhklWn6wH3J8RhD
Ch//rQR2Pf0iFBtQF7hBSKBwiiBw8ywG1JXqKwfZCeMVd4FpFooHJ6VSvYGGVm3e
sGa9GnJ4tHYuc9eSexeq4f5RVZmZTZ7isJoQumLYV6a1b5i/9aIVIDv4lJmt2Na9
EN33DPaRfdGm/p6hpBwxCp6jsQaGkPBI3e6YmJ/8JTcjqu/c2b38IYNpvd2MIkFh
nrh2ePppijgfDHLQtB1fd/xlcQB+IwhCH2vTH+g1zheXh7lQpl8+tD036I4jP8b2
gWP3/BeUJSW/bEecrHB1jCFAKT77jILPHpE/nnwRLOS3fH0ZCKUhG21iYVmtd/ot
S1TDgg5IIpaiY9e9M/V4qn2n8UBOrXDwiJNRA/AUdLIBVAx5Amah3XcWvkVdzC9Q
9CX2g2aZJ/uDo26W3m+qD7NBxMJ1mpYAuMeDU1r4KfZrc7Sd9S4UYcnQxWzHX1T7
ubg9cUPV0e8GJ4iHOQ9sBc8R0j3aLLZqvTxkmFanT/CsjMBb4x7ksYTHENHQ4MUg
J+ujPa7/v11qgnp55U2GY9rCMuUrEAhBzbT5SIcbK8oGQBvrePfg5jfLCKF9I1WZ
wvzJQUDKlilcn8Fi+wHpH5T2bjokzDOHWSfh66q+G9jvUchGz6K2DPpJooT1qdso
TKElWi5i8N08YieSacby6fwmyV2x+W44zZqlnlnXc84po2pDO0X+AmSKMX0iJN5m
RgD+hJUUQdg/6pQ+/Pt0Lh17AZUrLWrS37Iene8tjBAJReV3Zdsy4H7I2Q3muD9n
XbMyNAN47ry2U9QyGoHqYFv4qKX/oeW3iIFq0k16XmjEzHEQw+silP/QEHu/7HqF
x6RzNMETVX/j3qGm6fqP+cD8h9N7Af2dvtg2td9BptUKyijoIEzFSvnOJeC1XPRE
Z59lc79B3FQA2+Lq+sjBD/sUhnsAFSQ06xPXgBiutI7x7HIX0nvkeHj2xNO7RN3s
WYDa4cjw0vWzSO4kFKt/QPEPLhY6O7wycJDhKHeULGE+0JcLwpa+rhnJetMv5I7g
DVuY8ELt4L5AWz6OvAhIvEYx6kKu54iifntapy7EanNXjl1RciAUm1X+E7Zkv+H0
R7OJP82c8NqqFoPi8bStxDVyqkbiYE6Mbsh65CSucZiaqK8f9v3Q+gtqhYVbDTWv
Jvqag1d6c5KhpGFBJ1ZnxFy8NlzPncAiZCM94fLJO9+Yrp6K10hsVB5nH9kViQBG
bvrPPznMIFkoSDNKbtVEVaQzCAW/7MZspHYpE0cQDJCPUHrse+m6wpuK5iryx6yJ
BfSHfX0bqTww5iasoqRwQGEuhXvR1KO+Q39AkRiJUNvKAMtrF5PQ2FHULTw+HCZj
cj5rH8LPAxFKz0Itp55DAm39bFWNCwf8NL7ZfND/Q6ihbtu8ugFKQfv6TfsWPoCp
5vF6GYYvg5FVBZW7sxagvCNdk0sVqWkjM4bBrGAubxD70tFwRLHQzJOy+hd6Itqj
L/jH07CiHxRiOazl12XsSYx9yJV+eCyOxiHT71/hGdS7N15uCGC50NDSvRtqomYQ
w7C1U507OljUMj3OziHMKApcECxX8bS68mrT3K7Qua2bkxYk4BZqVk/UbRSxGta7
ql54bC5GCtcNKdfqZJID6bbNr84qD/+UQz7KSc8Hx8BXfToSJO/u+Wv1ydwW22Z4
YALq1EvK350ba1hGhcv+MpJ2We1pdu05r8k+DQx4EWrDVVvfpOTPFUMj8NpTb9CK
xwq267lJCJds/EzDZhsvys38lvXwtNoo+hyGwJbFFuM163gVpdcC09K0c6c9LbxX
paZhx0Y0+bP8RqIkJdYq0n9PucUAntJXnubMelSYGyNqR1p7aBOf8CmSA1cFmaVE
HHWm/bUkxR6aqdFZObJ5jPLR6IFJ7RkXEFtvvLIq3F5ktimgRz2x7sFDBwmKE71a
5Sx+gCzbhUVSdqyJpKPPdhZANjdMEye8+2eUud/OysrNEopfVZLlr7nfJgMNfUVo
zcnM7r27JIq3BN/+FFnnc1wY5oRgt+kad2N4/k3H7TUIuC6NWCudS7Dnm0Pgq6m+
vTbjV9nFlUVJ3L0NwhiCAD3Sf1mQzxs2xI+jaCOzJ3/g3T8KRoJeLkB+YUo4dvyF
v7yH6hr0XFNllzv7PgVVaSQpqOWMiQAEeg2x8404MqRI4zbsrk1iuz5CTrhNNSo/
nlEKFP3xvhR9zReU0IhExf+ecgVYi+ZVeg0ClBvyW7TGevLBCsjfKXbfThgnpO8J
XP50D9vmET5VCt/McTYrLjdLj+koLivvcNcpN7cfsgAK0d/khq9GYKGVnTBzTX5Q
HnENkLnooZpZpM2R59yosCi2e8ZMJp3EfiGy3CKrP3bv3MyOFbwh4DKzPnJ6EIeh
lpyYt1eGV/zL7bXEbjkhod86UkaT+P7dGWK/cXRquxxdw3m8gdUB5bDvr+6zU2+x
yVZ6tInEe+gnhDoECtZ2ct+Wt/0/RGd5+FRKSyyUvesc7BMiFyJT79h/pz1DEmma
P/NqO8Rg5bp+DotSaf8xmDBa8B7RWPncbJ6fws9vp452WMNkrASX7vAL5vRDDW9O
LV5rm2MtrPnD9Kdo+fxx37m8w2bsvHUN8tlX83JfEr2mzWIYLYnBigP4BxcJu7Qm
xTAuawCl28cPwTtIlDkQE3Gv/HUgVfynXq+dLiBH2M4z3rBDvmOjgHH35Fi3gBqM
1XlKZnqKGkw5mBtGLjquN1OvbAT0Jef8RmZiKF86ezdmW+pM/ZS4zJTwv5f6HRfT
EKVfipBYITA4bRfGFXgpouVBQgCz2B5h/qocKeRAQh4uYC0g7Lted6zDGq6r7/ML
+8dEmWgB4l7tW+4j4O3QvG8oBTiJfV823HyZBpGcwTaWy7gH6dnxxaTx77ucgdgC
oz3szZ6LRm7PBBGIWUvRvaA0cAej+VyD3CaAIwyESxo4WcEeQXN7kQBD2Fwtwtmr
xy7t3O4g0ABUKkOJKYcSWbdRWeeqQc0QyHKRTscC6aL4+pgbg3mtZ1n5LrW7Yh84
dHTVBu07yWIWQGjfqG6nX6ZKsGlK6ZmvqtSfEKbzXkEOLQ1G1DnbKa1ARcl5k3Pm
XpKeCk9VQP6Bz5eXnycXyXqM1Y6i4yY3olzKcosbO/YcOP1Zi+pj0g+FXX7GJ/7c
UwdwUaHCw18Mq2IgIkafnpFn6TXi+QnC9JjiJpFeAIslEIng26zHzbYuLqIhypvZ
OOiOaFZVgXSCIv5AG0JyKzq29S5/Km7Pd7fcWzvs0ue2zX1ccZGAVi2TDTQGD1zd
StV3gKBmGXbLlaGRk0jHLMOeOoPK3hY2r/ZbZnKu8wcS6sSBC8ZZSLT5dCqWaU4r
vgQm2UF03g4EG42Is7a9O7cAr9stBbS8QhmdAK2SZig1VXhprH61GOPZCYKHCDX2
EpIOFkzXVo6WfWP7u1fSY86Q5yfZfACwaBhlecPxtGKvYCUCMOSjfNqiPfndLm0Z
zZ/M/glMARO3F0JcZv+NZaAfVDdCr2LwroTG+vB4gE+ZynWL5jKQZiQNfEToaPrZ
qDa36kdtZxjCsv2F5R8l4VKVj7KGWnojYgIFPOfwBrdlwGNcLcn36RItaSP8bdhl
VPtAK+rO3t3dQGxlwGtscBMtYU673y1tWeEkbIHRrJfxTn67SrumgYmRiWVERiux
FHrRagu1wZaYcFdJKKh1VRjKpQYp7rJsgdFM73zQd09vi13YBNw5nQ4RON0IlcDT
vT+hTi1oZhPeVCEYwadiPoAQ8dItydHuMBBhpTKio2S6JF0/OdT4Q/kV+bcnTOrj
oXIfsRW7hW4t1PnKrfH2wnYmFPVrjKI7YdM7pPGwrNSHb2Kvxgzi4SjNgg+Vp3C3
fPGAL38tPfx92smgrnBt10+OprrrVCGciB44juDOrKUuk6G0ShseGdN+bnaHsGDm
yL1RkeKEO2suLJfhNYXVo1dbPpu4OOjPBpC+SFiAxrQBIgx2UNXkE1AmxARnCswY
ParcOWkyW/a4PLbI6PiJJzCNMxHWV2m+NkK3feUI4TT8x7qETSrqVzsTuumixvjB
UsZqbipgGbz4dRh8QMu6MnepWEv3RZJoG7jCJFet090vFJbuXDtBhj2QyXgozPQa
iMAUWYPrIlcsFkyPdQYpmEmlPRKwGJi9VdRq+uBu2ltplRgCqpdwdrlSg9cEJ0Ki
Sw7j0RbgwTjQYPk5fWZwUEuPn13rqXr6Cv0Rm6QpOlsTxpOZwK+vzkr3fO4bjWBC
ow58LtaQRyzfm/TwgxEex+3+fvwqARTTngcdeEvrKBUJ9FnhzLxhT3tVFwokwKxX
eRyYVMQ6SNlNcIdU3CqaQzF0XAeiYc51cWEQFaIhbrJD+7oHodPVPMODc8UM12Sv
misz+y1g89xRO5R+6NF/KL+ViynJDtyTsMyuEKOOL0n5mr94nGNUcQ+6zqv+rM/E
7kBUXjRRAftfgDj1jhTUzNlanW5V7h5Cbb+mtubXOISze9Aw8kQ4jESLn/+PGMEV
rEdzJ/c9eFzyHS1o1a7Q3RUL2anCZgnOHA4g865WkE8ahQ1lMeY82yD3rzhOloig
IK/BwDyHHWwRPCfwNPKK1ZC/iV2ofY9Nrg7S5FbQntGHyddNjdmaCFX3El7rcLEy
CdUhkycWB92EPp0D/X3nTjzJqmFlvZXWaJh4OZtA2UWCpk5I+Yoh222yUfjuRUM/
qEc88U82nsHkwenxpXYkbsv2tLN0zzJU8iMhq4NJlrcg/gihYFFk90LK7FR+kdW7
m9zzxGqcpjK1G4vt5yzYOg7GYf+xe0zaxZLVnnzkFTF7NZfaT9e2RNqugRaaGHim
pYBWo673ZdNbCF0AHuOSih1MnFOvWw3i+fLSoRulBkkJrXmnhODtY0c35lF0dm6b
5DEMxg5fyd7lqXYw2L4RSf13ds1Yeqsejr+D+YSetdge8d14Da1sBiOQaURp49Wv
T/pLOSaXW9gP2BOQ2bvcnZ0akZ2G8rBYoLHOwPqeg+QZj4PU+VttKp5Jc1/Q9yLF
H8WFjRca54Fc240j6pC99MyGaW9gaEUxtWbaJee/T/UvKvtJWjF+sjF2Ghhfs5VF
yZoelF6cfEhvCiBmGxaK5a1kOgHV0CxXlWfhn9N+kWBUSF1v5u3i184jf+aOIs6S
6T2RVkjwO0hUTyliszuEgEZSXnFzxLrvItBcBc0j3AvFhBTQ7ds4uU1L3rxEI+dB
bdinGZViM5pu4hAM6HtDqClBGdOvEg/UIEc/Owyeeq9YBOBQqgemWB9TvnS7OAVd
V0bMFkw0KHiqh0V4hzgnp6CEfJIGfP5mY4tabuM/inBwPJdf9X+vqBotcWXEfDgu
j71HoTdV2wEfXU8ZFWyFooRf9aPUnqSNr9jc+gsfslzlsaiaI+9PQSBMCpFlArsD
XuBj7gAl9iBAVIh4VeqoRUiqIxVFTNiKsiQ1PdBn04Xq2JDOf7PKMoJlZfo2HxJa
fTk/scbTcfPgJXd7v/Zt50l5rYuNia+4fteayEOheGHUgFmvvn4nC2ybjLFetWJF
zWZpRh7bp1he/PiIlPVtoJLticiZjyEW4VZGePn6av36dsr/b8N4VAnNVv+YEB1T
lrrppFZ94zwc3KLHymKqW6Z/y26ySy/xUFQBgNPmr0vXIX6wrPEZRxETD+eDA3Jp
kRjv51WZa61yqWpu1kvgkbBaE67N5IIfCUQg6v47cLevDsa3Gk+OfegC2fkTcPmG
IuyNU9kZQspTsLsbRg/D297vvlMaEkI3DCa2GHFGITq/6cJ49r44Hx7BtEzQtnch
aSOKo+49Kkbj68b8II79igSYUpKA9WMiCNNqhDoFMuAEAL6ML0MYuQnXZfqSWSAV
uCep8Sgzkfy/B8KpSfd0qztRn/k/fXAYab4gMzC2Sivqbrm5yuwaN7Sd1elGyhas
g8+C5uUvMLH3MjwUYq21w+tJWgI1sFV4xZg9CIxxEmWMS0NmqojdykZ78aOZzOVn
O0EA7WglzlBNs8x5m0/Ow82v7XgBYKbfsG56qTeUN5BllT05UnoFAC7nZDe0tsO5
KWcEVgPWpnvQpbA4ccgin3h1MDvurWG6nIvGd95Fj7olpbh4Ct+13KqBTopMBoML
HaISugPqhooQZZ+d/60MHWIxGB3W7HMtWZHpgDH0yiRvoYfaO4XkjaasCeNirIT8
mKAEmumytI1eRpS6i/VenWmPXbbW9C6stfzUk9C87TYfuSuKgGA8eiJ7LqBrbx4M
tfKj0xIGD4IZjctuPlbJFVYY8aIzwSqusPWrfnkGxpZaDjg+TimEiv9wBeGtqvN2
JPVqnIlqFX3edBWrG5GwzFswU0cJqopeA7rCwEwIdDyPdmqkSxOKGWq/SFxXMZr/
sFxW4mwkrY9Pp0KZoqRxYzvAWqpB3r3IbK009OkvPAeuXYRHhTl/gPfM7YQrv4vI
ePOdTLVUS/0YuiVwM8D6YiJh/7ADl3n3Vb36M9B7uADf3h9Da2rPlf8rbRgwOGEs
wvPRpRYIbB0MmSv55B/fSZNjiDxAWF1mG+F6tLqYwaNewyZZmzYBXR3/b5HJMaj+
86Y1k69gmgLAogfkeb5isttmbxHI4PP02GAG7JxAxak9rTHnrlLQkPEfGb9uFnVP
kI0CBXwo/F750eMWFnGTP1x0qHoFpPG37kZ2Vjk6HDIwQtZsug9pi8UTNM9Jp031
zTYB+h6vRSmR0iTodvadQlhZkIH0NrqObC1EccPxMb223E9qcybfln7PAPPyhGcp
i9hvoJRl9q7fZ6SazCDaeTl0cfeggbpkxLWsNywril/lLr3rwaifzMw8joGu99Us
tKTwyc/y0EkLx9ry3qGIJJ7WO5x6JU4eNF6Yv/PmmwXAfvWKGa3OAIGkrUkiGPnV
Ei3yLRgu9/x7YIL9caUg0P2yfu0pvgyyXOyjBJWhL+JIZVIcTP2V6a9R0ifNJacP
IoXVpSMDL+COtBVqXr0Ar0kKTVYn5jiTxb5qPc6ITS9luaI5lS9J79lP56qDXnt2
pAs5AKJhVKLAuY2v5cegd2Is5EFjWh1h3pRutgP62eMH5m8baXARx558yYbBfg0d
r+v+N0YTlhFg0Ct2briKOpeTjBKNSmEmEafKL0WTlt1tsk6C9Ljr/3zajLerOJV9
13K4fAuarUEWkrt0xAdx9EUpaUba7Hsa96dlXmomnFcW4rebq3q1AZIgsxPvIB2r
00pJ/+zvQdRvQI0pOj79yiHXuvt43SnqrJHlc6vmIlSzgEUvKC3HYVYtDg8KL0jZ
D6NOA/P1L7qE7nqBZ5lLQnBL8qKAo1J/OeCnMg2Y8YCvzbq6PxilwVR0x3PoTqEv
/2IDOCnEUgGn4Gs8U5IIm7hoeAeMZICrW7QKUPPcZzMd99ilXtOTGxHuf4+I7PSy
aP4OlqjVy3ByP6LXrcc+QQ2vcxtIEPb997BQ3VyruzSBSxKqCW73LWERMIjtuZP3
XF8V0Fu+v1Vi4u7JdDKu2F3KN9/yNgxPk5Gjs0wjiy+Gd4Uv2CYhR1XJ718STaV3
cw4yAAOVP/F+irCgG4A/7IKJ/CsE99qFFDQeMTi40p3DLxXYFCVtlisfG8BnFjXP
ZVlPlxP1yiCR4pqUxVT5sle8cBW3PMi1TQSXj8gGCYTGlF1c05mi9QdvQ5B80WzP
hGhOY6+J/RGprke0VJrHyo75+oDVN5bMVLNxPsn6LnFCOuSGE9hIavnMlhsc/Pei
hZkb/dVkgI3rnwCbsFKl+V55kyTf6cZa51hPCKleGZ2p7Nf7D9NcIILoeaoAliB0
MNPVJBa4Ce3t1Zp4ayGe6X3Js0k+nALOgVGEllpI7l9hUCGOENddGWXg4aguQ6HU
dYtrvEVD7V7QWsBbSSyQOoGNXRzbwa/aS9R03/4W8GCp7zM2+g86LH0RJcGvaMqF
99dhkGZvnmL6J9iLzpP/HEUm+OyI63Ik1LKZikOwN566G1JdE9+idF+gcgDZA+YJ
IX1Llo/5CsTHTaab02E85oxCWC+JjP4DE8MVOpFt7m55CaNKSQ0RXbBujT9hMyUr
mhtLJ3We1pO8BTUs9cA5ywppxoQElJ4lZr2M/CQaDSV7sN2IYiHcfCdaP54ya8fg
PbwLHX9Is+ECFLus6B9YeGV8xfVwtrchWe0L1rScJgrzJC2S2UTbT2dG+L5GWB65
1J+EkUqhWkVwU2XdPu8nK7I9x5NvNjCedtQwRYbiODPFtHXoLFi9GsfPoddbxI5T
zkZggZ+13nzP8uKj6HdAWjS3WmImSQ+23EiHAa/ytM4MytSsGFvpe+XcABf7GEEH
LeUJuYRUf5DOuOzII521JBX+d6egb6gqCKZsgWgVkWcVf+YevPXWKulsmJniBNQD
YCRCbQgwqbg6Z4zucEawyrvTsGcXkT43e2BNU0pl0bdSW9LqfKNmuOCRqLaPra2P
KjPywWt2hJjsgysB57khL9KYaSINI35SjF07zrMU2nwvRH7qTZJ9aI1JUWhc6gBJ
Qb5qH2UKGo9vXjDp9Y3Ul4Ps/6KL6+I0vDl3RkvglfjIvnTmvTdOG0Rx3Fm3j/Rr
fXy6T6YuYpMlKHzAQxMKVQdXj9T4tiyWTJdrJFEmfzL+Z5wv0YEaDIhXEqHfdmfx
fETXBhBuG/BraohilWd8svqZiBbKb+Z41mMBCOlpqCg3//jw6PS2dnJdZ+lRJha9
WuXcVTIFvMjpSv34F531N1GvjBgjqcqHfh/hz6dm6pHJJd+Lid5dR9LfOvdN6tvf
+oO/kV3mKCys4qhbQd7uWFaD4Trg8HQCsGIsDiugRfR0e8U7Cy/ejNnyY1nTHLgK
AM9TrSp6tXGEWD6OFR6NA+yjpL+VTcZTWX0sRqGTRrrJ65NvFVBcS+QHSU1faveA
ZjFeI1WRuOoBya7f2qp+Fi0956gXy79nRPbReoG4fZT6Pu+8lQD79hHK8bmnnzGq
Caph9mV7UkmEsoZIe7p9giy91R29LpXqqufMYLeXdMA9w/nMv6kMOkT4Psmo31NZ
PETIKEA53dAtguQJ3FpjdMNS5WG/wLOSceErnyg1UmUbZZ/mKm5ia4zeCoYzoZJM
884NKkP+T/jJYZ980rFH8MJ8SpHcR8B7+eEXf1Uh+ng7K1N+8cpfMoLKfoCUsxDD
1Mfb6E8gh9vShrypvRQivwc8Tr1WAek8MChMfrs8OZDUtguHYsIVMJtjc/XVizHT
Oh1Se7BRrcQhnugXtRlJQ+bqqmjEr+aq2R2KcAEgZf0SuK8leo68DUfmxySd04Ou
H1PGk2QVJWwT8jQp1Vi6xq8Alggwi9EeNm74EW1wGhUPdJqmBgzF3M5FkKVz4/zQ
+jbxmUnlbvWld9FIqbfbFCeXIx0MR0+QMGDr+pMMzYLSxP75X5KhTHVEo6DCWTni
p5CPF3DiqADS+E1Db6WzkHs/7fKgCgbcb/sad0cVc+sgUBKGFAHktVrYQ0KlIUBk
vc+5Ex7sLdpv31w7Sgcw/2c2Ec7Bx14jvjQ909O2+WV4cDGLEyaWJJopE05pyBG4
wrREC4/A1hrD5JhmqYBWJvcwp3VWkqC1Hi5Z5ZW2LaIr97pMH2UVSyTWUbW2zTOw
izTS2YPMYcorge10aMb7k03DjMjPaeCmsoxTifje7AT8UMtPkeCSgnYYJ0XImIoT
HqO/5SSQEIp8UQfLvs52oH5oT/bF0v2AEKEsEStzjipaSy01RxlRQCXtFPtapSKo
F8Y2p+lRHp9gLyZT9YfzqnBvPGaN11eMrMU9gy6vIwwcqizlTy6zaUbZVdiPBjWn
J7mOw0zrSPHgL+D+wVnWOOkq67T6SX8Y34oiI6nrtP9iwiFul/eERKqgfmO/LsGI
rl6bPHrP0bJc6bJ/w5o7TZsBaZhSYGUfLELPsqNYWoqtrihfphU1gGNOHPt9ON2y
JVciC1E7XWPbcVtw1XB+EGOS20+wtgBB4wuYYKJfbeo4LaWoHyV3i9EGlmVORmLY
0N63qp9j7Hij9IMLFx4POij6TqE3xZ28QKds/oZxMbV6k46z0G7P1i44EIGoG8FV
Tuhn+umRRr7GxmjTwDSnUhsuyrvY9RVQkGYRl4gpe486Z5mqQziQM9mZEtdIVK4K
KnC8tYAdAMCNMI5XCi0hnr5qORkx7XWv15jsYNFZxXssZvw9vBfIsdCfaK/IiCs8
p9zNb5rLDPCT4g2+uGnGeRSJMGdNKkg1HT3oeGWsf4zZ/dLZHK67TyNGjBhuM8z+
ZXY1JaSx8eUGz74KaXdhs7+okEobU8ETR5Vmutl2pBO3cehks9nJLSrmJ/UCIUbB
I3xiG0PmeOExkeOlWAXhzuoR8BCl2QqWrbIE5QMyv12J7dQpSF1lAY2+Wa0jQQ0A
mhtbueolqv+tkYICwCUWeohd1stzM2a+mlxAs7S9KB7hpoxsrsGXDwJWBZD04Z4I
vFIkFeOJPOIyIG/n0YCnhZ3PwOIIIubQlEQMl8Wotp59r3wxgpxn/3gHRYTEFLto
NcI/c5BMBsGrcDWE4HjE2qj2dwahBM1B4tGvnCSnEsECpOaHFx9B7lURPWfn9Jid
PT9iwPcDBm63Y7ux+0D98bdJy3a71BZ1rdkOeYC5EdjvLYLs7z4muQ+EWBuO/0/r
7P8hloSHbRBSUnP85Jx1vlVqzgb254CFOIzRHNwt/iHvKRW4k/616gMWzGwIOzOI
UcAtZ+jsspkybej780tNkH+0J9hCXjeGPMGscf2sDZxNSKURU+LqkJcu+8MjdOIg
OabgbbAFb4DUlk7Iu1AIG4LrLDOzaXJarsJECS9dWX21m0DDqeVz/VmyBjpNEcjH
DWzPL8n98GAzEwQJJOsnu0rLUzbb8RolTs3f9X24+16imA9IAr9aYvXHqLDGQhGh
6CMpKic38hF7n2v6GtnG/wkpvDtPUq2sb9yhEgd1QHkfPiWF0RfHCrXXOTc/9XD3
1JVCyFmOXaEe8CKgwalvkFV6hzy5wAxeARqQN8gQzUgiPLAdARyMFHb/12IpLhCo
HmZRfwmNtLOt5MoJvRhDl+mhfOLOPm2Vp/F8jUt1UFa3pogxkpYEfdd8euSjdO3w
I6cS/t5sXet2AIadnHSPDc9vBGHZEazzoQ68Yhu8DVxUsZe3mZTfBg15VsXaxwLj
hUSHXDyFJM2Xa6lkrUmFo+XgoeYpfTEI9ViqEeH2TAVSjXaFcPXhJDIuPm1YgPzM
C1Cx0CsnuS3RPLAazflnmWOakhen8cifxsLe8zWeWK1tLp0hwBVZ/0+U+E4/xO/a
qK5KbSOCnfi0l7g09GRpXZRPkkbdFo9eF0+tqPPRmRPz9/6Ed+xuFaDzJrvQrDEx
t0P+EEEOMQ/DgfDwclUXZ1EkwBVp+UK+xOLRL2wSfFO0ZNPtyMjEJZWZ1CzpTrIo
Jo3KI2rEBaREKQIAPkF9f8a7AX67ZAUk0jFHHfLScuKgaaetUexn9vPAXr/gUZ1s
6Wm12rVl7gIScJWZQW5HBueZgzT/lsvUZayqENpNjM2lgtSAoyvQ2ZdOI/CqKa3t
kFrU9JKAlXUdCXx6RmD4IWvynfiFN79kG4xt7x6qLMTik1lkxNWgKceE4Td281ba
GRGimMW5q+NegCTXFH6T8WilRe2voOg6lOtluRLleFlPT2Z1M8pXMWMHiuje5qe7
MynMO/lIhMNuPiSX5oqEkUjfonMV8T2OI6GZlJ9tZI3k1lwJIHGA9F1puc9XV2mi
mn+0vL4yjNuI9lXQ+vIr4U1PyjRORDna1ykEpu+sRzXiCil6bBEAby3XlKM3qsym
nvriIzB+LB/az4vQEBKX3okN01i5pgs5ICMgRFgXVDREhSOnC67HajtRTuVdEJyL
ryaVF3Dvetvl3Aa/M16zndxeGmQZNNpbCEHxFhK/OzklTtv1IcRA9O9UF7cKFk2s
WR6wHIHxKd6ptD9nPvJTqMXXrbljms3MUFmecCLQmKlPclLxjx3g9LjfTO0Qzp2Q
QAVoPf3ii34HpLormSyUGN5teNuVRvi8IuLrza7X34XHqkFmvUqspEscZ0xAf6aw
I63/0KprAssqbw/uBcLqECEHIoKiMEfJf0+qI5HAjdS1FNdSHs3u6/vSBxHtlWHm
afurz+MfJmkjwE8gSulAVxFQYuLyaSiVc/9MnHb1TzAXE3/ltHIQi6jVChuN8Mk4
TKmJdFV+6dkFnr19hiqYqsPgIQyWFNvJQTf9M6SxMqbj3iUC3Z8IuMe1ne2DNE+3
/q551tglwJi0mmsqPdoY4jPwNegLaNgoFMKzt/gHjV2Kqn6lLJKCTUqdhtzvV+W2
lB8l5JzOZNV5cLImtzD7sJcvtayfWAB7m7s/OWJprmo0ZUADyKtLkLVVo/4djFsX
DlB+8D2Ley6UPRRZFYt/dm9OT+28qThc/W05pXHMI47s7EqPBg9K2P8mOjm4wnZ4
ku+earEYVxnQVM9bmNwEGk/YDP2bqM7IvI8WZ3Cukj8PbUv+nvuFAntstPiMpRy+
ad1Jz487iT9Nz+caWr+oKbsWpESQAhHTkWYIePEd7sywGjaCunCAzU6qObnnJ3Dz
eLZd/1cdv9l2a0W88Vv6y0WXBTcHeWmLcxE1DqU8cHQltPGPE/OX5jQJcbOMUYma
pgsLPCY2rkN/HwgtpKORHWBrHEpBvKuBz+oGZHgR4um60/ZJ0Vwz429f9cwaLPrY
vIEmPALur9iiZT5eAc7EWbq10Q3p3ee8dJgg2LI77WHG3/oQ3GLTeQ10NI6YzZSb
VjfgDYFOmh+5UpTPgMc5roqK77iWzAfYIgmIiBFJv0T4+ZFL7aIVyXMrkfRTRbLr
w4jHglgK/0etD28067g3L7rDTiJMTE1x/H3wDiLkklv3bK6i8vtZDH8JVZpU/njr
sUXPmRpMeuXUU7+/RjoW3TccNKZkCdOs9oROfAVo+KmzfTyuj0eUjvmEjMeDZfZh
7VS+GNC487y+w19LvUPG2XLPNeE9wuJ4zRPUsM0cb3Nu3HWBr57ugecnKO6LZfgm
nUwfu+tRz3d+CFHKRBEMQ/FaAEIa0i8+f49dW6vFg3o8FyDk1X5SGFYb07wTSzwK
RTsxoNxZImlHods2LKxnePgiJc2rZUwLPx0XfhEvpDJ6/TIkMULlFG6kTJKfZBjH
TX47hUCgXljvny81aqrl6+Fp0VhT7aRVm7bywREy/pbg+LXPHcx7xZzWzUCuVeQv
qMsyVWqy0KUMAjlJsIxMt/zrwmh/zFaMGqmahxum3fHBHToniNvShASewRFW04Sm
VWVB2qwwUDLso7973hm7ITdroz07PDVVoMjGD0sllDygxaHSNoYT0FmiwyZCheeF
k3k/iqJZ/yzeT4VebrFyXr+D5NQzqk320fnSFEbzZwtRkeuUkTRA9jkUYAqvJLms
WGnA/oD6GrL67OVfC0JazgZT754mJfOP62j5sOGwXIzyNRobpK8bgHOo7GCUNGz2
kjPceQj0plRxWdmfzYBgsKNjv5c/0nAgfahA/1/Q5s0KwkH+0gVbMqWXYVYO9xci
l2qUMqljHgRO+3ZEjdzaoJVwG64TpqkPr4dek42GagARA99SC5MCR9kv3R+ZmbqZ
JfzG+GG9YlXjd7IQ1NdbWNQIPtDx8Erd5gID4uK5wcpD6hv1I1vG5rdI4bjhSki+
NkFoaqhZ9mOtNOJ0TQcDYihDNyP96CxfHro92RlFD9xxDUafbkFoaXWPwVGeviLo
1w74PMLAcn8Xbj73bjv6D7FVRomod1A8ZetxLCm7yw2nwrSsIIRby18S37um5mEm
AVKWvR8S8vT9Wr/CINi70wus6FoI9NvGSWX9dx4JPiM3EACVw6YMk+3/DzbHNAuU
yMnC1IY7Coqy9UkYrS/2r05JhMaVLkakMmzL2G+rYdTivFMOVqkVBuTpEU6EOm0e
izqOvbBbBoqAlvyk7d6rcfin59hx2NnfWAQnb05uHELj03xDEEHjSumHGCAGXtgN
Pvvu/jzqm9cTnvUVf77fLOFqvw/Tf+x8i1NAslgPslKRmiYWNAq4Um0M6XK56wbW
yy/I31eF9tPHMz2yjgRL6F8FJLTtiS9YI5uIbh6bdtZvb0O22qhFvq4aor3wOgO0
VpbDZtFyU3AKI+Vyzm5Nhla4p+KtX28HMeLDsPEUuHBvyB3RGSFHelnRAE0wrGZM
D2a3Jr01F4m1qUG5lpYwNGwDMx6w2XckyhiE9KqDx+XsLzU+Gh0AXJaZMv7md0r/
QuuBLLCTYphNywfu8cv9K5ixJ78uC0XXfmd6vH8v+IsMsD23csR/YrBQOZOLrn77
cN6AlNBf+IEBYTiwrKjafjYzwcfV5U4F3ukoFtaQp0J7J36x06miRmua4AVd8iyU
l2CoTgByeptn2iXLelLaZEAH60b8jex0LiqACpXW3YQjrQisyqQBcIYsV47w05Rx
DPpBnao3W2beBq4pcwzqz9mgCAUmdDUcIagOlVlemoCbNO11thPDu1G7722uEUnP
IUtgUW2DSQ43BERSiSQ+koAQ3pVYI5Ol3Aa/5RB1PWtjeS8lga8v7hM/qWDCZy/f
BBOh2MjgLACHBXbSfzLypg2s22IC835SP6lQJYrxZZ2gUHapBOK/9Y5z3vuryfcF
3iRRhi+Bdbs//FQYyeS+YapsuqAgQeLjOtwnj53Raw0Np83Aji10MBuyO6LkRLGV
s/aPCkycz0k+VgBehvMltMkQ0qImRlXoxuYMTcIGqMzMagnQaEDDaxMA4VDQgSas
XI0LWMhNavms+yiwkfOCOZTZ9Ap/Uw1QLbqFRrWQhSzMUJMHQr6o04jxPsv4QpLV
L+yIfURroQH4kFFN2UIfgjKh11kIrVAdx/vqNaIv7AyicEzS+uNcV/QE/RWgB6fC
oQIsuc/qFFufdOgPocprJRpZZ6R9lXlgNMGrcmQFBCV+3QWaJfj0wEn5myA9PJEz
srJB8xxZmTa7mclpx4yTPq8M0YzF7iXoG6TZNSj7XG5eWBgwOpnFSvM/OHpTZjTG
nKoM17ZYLAGjxTxNLqCU0tibzKQjn3WhsGCmRmL0whwd7gx6M+QMXDl2gJ74Qqa2
viJnkF2wp93R801G3ZaTCDUWbuRPCRu/JkjSdTwj2MCflgI40aUaQ8aWYAK9EGHU
W1K4JV2EN47hHWsffQ3t3KLm1Lh3t1cC/AIL2F+vJ72QIZMA7Sz4WmYbQphfp//+
gG4WVuclHWHuWAjGIQ6xl/CHtbp8HU9nb6y5S5ztfzpkkTzYSCvC+IUed3yqCtQY
rO+hVqvlZoAdP4SwcZycv1H/7Wo/q6ii0kWApJA3Acn4itcl2ZNoT0wYQwdu6EV9
I/pPcI2llVAzpcQpzo3f36Cy140EXyBiZd1gekixKy2HFQd2hx3yGkSuu3oI/m39
KymoJkbaKmtH2lJ8Ix3W28Iya1mck/jPNExAa4sve1Xq7PbORmA63E/oLbfqmfJf
Vx4OgZfMLzUeiInSV31ujcdlbpgPS8Z4CRpHfBC+xafIC4+6VQbR3bxWDKblnHFY
OANc/MmMFjlLUTCtTIl6vIBAAfnMkl5MpMCTv5qgsEhnobQ9obBWL046IKWHtrOW
KpES8Tcb5zSamE5wBBb/xuPRp8pRHofod7oRPBPaleOhJ38ZIgI2g46Q+CjFM31B
fThcdzHaVzp3ezeGjEQRBRsVujwHWQN3yDxGtQ+OaFy9z6rmL4Stce1+0Vl2myLM
nDF3iIZ7zyWwzdNM8e/93bkHDJWVqbf80zmueufBbUflnHk5aOkNqanSSAACUdr3
E+/qXAZDV9b15Ib06Dh0TT55gQOkAcHHaAXP3YPEqGQvYGENObw3LmWm+8YLSCMl
HzrfBYb2yIeLjx1XedaJBio+FGbqestdmwYy+z1+XCl4VbjA+OZeow04DJ83pzrT
BMFRCRYV2//cccqfhs/bIP2/byntO3dof2Xd4He1QZvKsSwtwgiRUqLQkWn61Pfh
kQoQbOy9F0egHf4XcgvyaGIne0B+jgbvL2hconqd9Pn1yHSnBT0yzuU/7577BccL
Q8wKCujBB7RIu9gDgscljtiPU2Z3U99YIW4XzgnUMPjVEuX1bnkWiVa9fnd6CR9L
1MsgMLPTmZ3DF1zVnJ3B7MTLg0JZLthf1HtNoOzUnPnaOU8xVRITeoruwHFNkA+L
kKtJdkh9iABhmg82/iu7f5Vz8axCBMM4UDa973AFWe8Fg0ZuhXEiMmudp7hCxp/H
ARkwvuQUb0MR3kd63E4ErKP+NAmOH2vkT6vNwTo1QibWUjWlukiPbFLWPeddzU1B
uMQOJZlUWPBXPAEGdaRNajEowry6QqGjIl/E0hDpi0LvQB7mqZXWx2FiVMypZjx6
KRK4l/cx8VPb3uzVOwBtO9fAxPnqdsdmZrukvv5aUZO1RepJ+CAzUeM9X3XDWC11
N8r0lUkVSfWSP6gIKWuRP/PfCSEeiwKXZz4J1Zln0MtcsJXU61E2d6bkmFkY2c82
QbMc7l/I1oVvu275IH8mt5KJ/YTqgW6hslkvQ5C6zZLlQOpbzdd7759T49wgmAkH
yESv1OsItbTmyA6801phltRtP9Xu5WHe8pM+P4QCPWOYxQEcNR4fuZDBzmYbK7IK
iu0uNKHQcxkhmGKpZg7tW+3Dr50XQcmO0rSznTSlKiJfzxrMkGW5Pi6oNF+8rv+e
cmoSsIvujN5pjBS7SBCxzMJ20DnRErGVM7xiVhA4TqtGJjjD6ppEzwMpWe9Z7vXx
viRnFBr2ogyBs2K4IJmrzpCNYIRhCmtyjxLP80x17a6d6C1MjDr9Ikrjiw0iTd5D
Z5yh28AnsRNyaT1HIxM6Qfywgh5VIfer8PSNZa6DmMiC023NMrwqZmk364CJ/oGc
k+Vh8abhukofJvpnR41LbVx90aMy+M9wiVx5TqOetYSJnDDS5PA+CUX7cK38dgwp
DTxg1zGoOxv7XizmNp9a/B/kmj32NS5OFbqYyS5EzOXnC+3yY3emIz/i1PlWPUA+
W0xPmu5Evxjj0b/f6aLvyF4T7j7FtzEbtrxLnDjbVuUSoeTMtzewdn6Zfi8pZrX/
nCrLRyfTZ4PkqpZPfj1aNEOpof5JQEDwtQW6fEm7uD83INdj0Wo8k/uWP+PvzRWy
3X2g6p5//FEj9oysu7c20V2ROxNXW7okVMJRRIK55gLwp5699hHLslSYxXocTski
Be/banUHwC/0bew1rU3XoXa/EVp01sQjw/AbDj1fmJAJQXEOhJ6Z1WcqT6ETb/b3
shN/sNogbF/2lfS/HomQ8ZLJYA+bFNQn0ojc493i65YW2b80e1dkfca/KPiKZGpk
H3jMEqSy7l9h2Nn36N+KHxJLLRYXauDb46DLYwqi4zwp8+z27xZOwkJhbYig0dVp
AdHjTT0/9HIU+ZBt1DtSrH8GtBAc7d5Iga9YyLM4CBSWPv2zWipfVYFGPoW8sIIF
out9I9KOIa0uNn8xXjQU+c/TQq+XKO4AlHSpqizrNszNV5Dlw9ojxRsr/Ca9I//C
wTwhbyOt6eI+EvgVtfN4DZbFTmSO6jvhJxSAqCDk/jfH+JS/qPvfCzqt5EoHibAn
S7ZCKZrf143Z2ICw9vFcsYt6bXzDcpPb9PCVfvFb8MvfXwPRpBpWvx+cdUjGuX79
NAcPANmPO6YKaXVaBc1KkC5rPRsGi+5kLB4ejywUIInvj5z8BFPH7oXrC1KaW/Kc
h6tzUlN+Zz5zGbAJRZwqwOk40ViC4GvR4X4mZin6GCvKoMwz5II7kpqZKTrXaE06
TMBKSHdQJbFr+aGo1GQ9MZ9xw4ZpOjYgW86+eCwyCjAwhB6728/eeYNEq98acPVP
T7K5aADgvFJTTv4GFgzdQ71uD7UrGFDoNU4Kw84OsfHR0VCUTu19gsWxt/SUvAbH
SyXcSt3qh4xX3nFdDihFcy4j0tcTrZX2M1BObnLPHhEsJNNIKLIpTNx2nHE1G6rf
UK/WYy/Kij9VCUVO+LBPfuxGJ/EL0mbXwJO9F8V9axlYXwAXYc93nsHjh/HsygVK
S3rQtk7Q6iqvLPrCKyPXZtfv4/pr7Ty626ZNrbje9/ZJ8yMhHtcjHryuIxF3rDNJ
5xuktwpqkFqJFxlZrx0gJYqYioDc2ovi+glIbxIzAmVVvknVAg2SNFPJEH9tLeYP
OLaDi2B7W0kknVWPntLACz+KOtRFE4hjJWBQFiLx3ENGLeym5UNHBzvpoQDvi6n8
4l2fEmFFh6z3QeAEZMRQHVekDbhkA3/3pG+1og+0ivkWUZJUCbqmhhF3tZ5PIaMY
pD1CUCJNFAaZcYexitIHbv2cRqAbIY0isUoONEO4tBl2ut634ELAy+HMq6gLV5gT
8ickB6r7MRx2GsBrQk4oTsI5PUr0/3AZq4QYcQCEWZ8Tsonhh6RVt4cwPeMKpgha
7wgAJ/gPg76HUyICWa9WTdG1pOIqkyUdYhl0TsE9ns24TjUkZPaYOck3Dus1cyUk
lKEOJujkSbkQSi8BmJizrff3LF08ucOTSKygtH34z77sXtEb5So5Fg3FZVN3N0JQ
7ciSnLHYd/UEJhZu5I2jNjpBR72o8AkdESX5kQfP8l92iTXPaRCvhNL+G1G+JJsS
huPVht5sLPl5NFKJsbT1SwNmJXUr2Az6NUbyyGCRjhCJpP3D1R6K5aLuIdMikzI2
102tJ4rvKBnksb9R8NUfhPaS7NR7QGL/d/kPCBv5smWgT2k8iZj9dzRfueftrE97
ry9JhKxkHBv1OIlXV9qEEz7xJ7gtTQPZxq65r/Qto4gKweEvEACo4iWKnQTVETaS
tNmwogYrs5EtmVF+zqHTjZR/C5stLJxpbOl6ivZWpHIzdEV/SvASOLPu3kPd3YFN
TE3kARpW3kjb9TX54ZKzrCv0j6ei+EZ84+N9Y+5ma4vL/dutltgfXjIl7eCQkUsY
dP288fr/Uk78lJnvkfyHK1f771xgMJQkSQacUVogBLiw8nWHvhvQwCv4rdRicPHw
XIFmEbz1ZbhlmIBwvMgyMrCzcDVIvY15QDTfB5q266SrLpc6XE9pD/4jv3cK5UqJ
+VgbfO6EBRUPJNT+Uo/cAHveNYOojMaEUXjp3VzQeYSAoNsBKY7e8xStu8yTJfl+
avq+E0QXOcjaIsgvSHzouSfdQyG44a7fQIQkHbsg6x76GmvELU2WYSHRhtev+1al
kizFU/5at0A+rQUdtEiM1sYgXZ+go7t+hjctwB2poFiO6FcIO1XKiuSDfbkKUwXL
nWQfgqHwKtnlnQ7q8W5fJyl+v4GqaJj1YP7X0pip9byg50ecT3ABuCvw1Ft+6cnj
qDwNQEqnnil0/ySmmWljflnE7m3eeL2RTGznOfjQ3/C7X01Fz9VyPckLKXzd4ixf
cxFdsDlser5bxvVD0vo751/1rYUk4AwZo7d9TNaF4/Rtbz5RqbOlMqf+mFfN/piG
t+DC36eU6pZkq0m1TWeBx78UMCI5hTfR9uWnpVLOeR6JpFTBrgvw6ZVLYj78gl61
mgB0M8QB/62qD6wDKTrpjio3QuU/Ko3g7tafeEmXVsbY8dnqw2B+6P7vRajkhUjy
d+j4bAJTGRrtcUwlukoYFuY+gqAmezqeANzy0wg233+wLK2rPed5eADeE3+XwNYw
+L5UBoU9mAh7V9ZPKmYBDr5YOzHj0q4leMsRutr2I1YMqOxq6pRfiOkzhg3+/L0L
2tdQW9iEtu+XvgX4sIVZ5Gv5cBMX3RCfqIXnKYE/kGta3RZHsdX+8HXs3quhN2CF
MHO4LQlAKWUGyTT8Irc+4wc2ZPjDCdLRXB/d8PrABEVjkUc8MXf5GeeSTegSmOKc
93wwUK8tAgGWmFzv4XuzHI/vKAJkPDU/aVNelffUbeTib68SccEu9HG/C3kMXqTF
/yXAhaAT4FRufb8mErLkIMT9dJi2UYLub5+XLNd36jovyGWDqzmdY+bb/YNb/EAU
m0xjAp3be8fnbyw2mtBkrUzOWupC9Ki0Q2YH6n547UDCGPczOHeEJgqQNhUGpvn1
GA2+vbZTOwUjbvaczwEaktLREX/8AwEDa7ND3B2QFoCrJxUoOBPHlTTkA/ny8qh+
9fLL0OQeNRg4sJ/+v1CRnT0Js04c4tzQGvVE4ATRCfvFZUkK5BVC5kwCwNnXNgXY
b6k7eBpqkqvBLJEe5iAqASCAlmfbGaJ7frYGpLuj8StJmFzEqrHwK03z70bg6JyD
eTJD3ILjqShWuoqMkS7Id8r0zgwG8a4Co8W1XZjVeG3lPSGQSles7W1q++TKQ3VR
lMgHy9M7MuT1gsauMvWdJ/7iPy4lmd/8dlYaqQOiobsbyf/9muaa8KLMS0lEOpvG
vozpdbPF1DGR3SUtYkdikdR1lx9ninStlqKH8TYPgujhmkiTqUgAEK1hYHHdkLVt
HU2TEm01ffmrkaUpUIjK3DpeQQPNT1x6xpnko3kc+lnQ+5eCbXXBFyvmKulzDl1f
CR2HalOWlh3KqOYCllNPu5HH2mNEBQzMDE1Dn6Zil5PM/np68R667aSfixIC3Tuq
PE2hGcczEmBD+x+PE2nkDPK+srObAbr/+VOtAxLbisHb9+RIH7LD7XtIR8Sz5pB6
63Cozc+lhG3DUnVlWJ4E2WS1ZWh3BIBxA16DCWJvip2v/Ka4QuioxTIizPs73/4c
xHoyVQh0Pv5Vpd6A/wVk9wIB0P8KvDh+dseW6G8lZrmXGot8aZG+/L7NdyjatGYu
cSJ1bKldHbnZyv47S0/QMWVrWIOOPQ7Jb51BmoLdoWs8SnfFM6rm75DKvAQ6gqVZ
CDSe8GrgDWTLGPPrry+ABeBdu1OrASBx/ze89wAG/sNxGxgTWLfFGBJFfv/MRrhi
BHxu1bkVNW/ArcRg3SLbzn2bsStsaJzTHO6Aw8MPgKNQbNSfcH7bZ/ObfnJ0wXpJ
3p98tbC+aw6nEXQcAlEnsWNUku0LyfNiBTecN5CxGCDNLm1Hzod2D8H6Y47ZIiy2
8wiyaL4l0JxMT7tc2qvfBbIll0jVBYoovXe8U0BptFvu8pt2WgIX8WWnOZkfxV0X
Ng++BfeTX2axKFbcJpl94JD/qVSR4+vSXQHIeZTg5se201bTm6WWo1NN+lIHrZaz
WDFIqFZ1ifeXcw5Nm1DkupG2t5SR3Yr1HhMPvb7T2UyaPD55mxlgMsbyycDeGk7l
/ldYm1zVmjpOZP8+WaKsqxTDKT7uGfEHJrSr2qJgDR4ISnSTbzhkc4CRSVJHm9+M
HG+fE6n/UyMvdz3CIxDBjy/mPqI0SeAP+k9qyl3hq4mnX9nC64TX19PPqy0p8yTW
hv8v3fKusJTt0pLEGkHrSABBRuxZ8yjG9+i0jpg75ac+HaMI+hJa9vUvdHBp1DZB
RfK7DOwrnUePJ907Of4kisXLdJ+/Lgq4barhZndIlQNr6rtK/Q81haKmSuRmEbl/
ozStzwmTyFM4D0wwmm8pNAsf28yFvOcdiWvORJX4L5X56FblDUGlKF4dFhbJA+pl
B3MRoDCyB4NAN+HUFwDhk0ECjnVaGS3kEfXk6zWPhvW4D6qZFkH6H7LFCGlyMGoj
KJUPmfQlqUauPOwI1qEGBwLpviRFENFNFhCHL8fTjCay+yCwNJIW0H2ARnkSYl99
lQkgqwyDAq5Js4CBA8uKtRbiaFK4shNKNkpLdZggbsOJIOoQXawKZ8OqUHx66rPc
OHz/waoU4VoZOK3cr+2pVwVpboewzfzTFP4wB5H+SCT/mxdqFm8iXgfsnDdFuPHr
Nk1QsK68J3nchr84V1ZjXOihy1+V3GV8mhX+hG03JnsA+L2hWlDWuL+8reyJzTmx
ct9pn1lSKg63rw6+6/faIMnts/JG8xBUbJ/fH/d1olGFe0nCDfzyf7UIZaK0hoow
ZbXeooYM4rtKINDwdiZR6Clx94g7nTbP+P33gRYmZb52fW0/d67p7VEouS0z+Wsj
r852RpHEaUQGS/StKC59oLqDnFDSEf98gPHVF+oUA7souVaryNeAYj17DlBBZXt1
Xkj+RYmwxKSEDV3stbyfHRGKqO9+CaL+gpdErzxy08AUKxv1o8xWqn71CShu/1QE
/NSLRgXvOwvBoUenC4Zf9IZnum8qcr2UZ9PEXn8W4X9qIAdo6eHLlVGQmZ+6x36z
0XpOpX0Qf0mKr0NgXy/D2zxMYKjPwQ+4p5lr3SCswIqxpXJ6p9MwmmMBzuh3Y8g9
hG+m4XJJ3oQEsKwq8OjcmUSBpSADX9Ntgm/hErUP8oH/gMpOLKrO+zoELvhpW6Vw
A/NqQH6YedHSo0RiPJ75ooUGIyTZcXbVzHq5VRe64/MsyH5615Kyru9SMkuVt0Zd
43ACSFh4U1PKhWtgqHj66yhIz8EaBtaQyBZhoffPr8mjCrV8q8/ygjEOR+k1zXLC
oe8NVd41gFFyIj1mHmSoRkjOyunxwheS5oa/sI4KlWvIlwnHY20sIv/tY7AKGwmS
uu0ORH46A7yx1gZ05WjGZhOyPZ2CWGvbiJqMFibS5GIZt8ZNQCvDURRqXoMpPSx2
hEXJPYfvfQ+y/EO3BOSDo5SoFgp8ZlaxXnitioCkl60yzokzSAo71RH4RWuCKavq
Mm5zcrKHERKgp7BhMWz+HOeLDhihsjRUiEImpk/IdIyQUbgTc3WXWY85gtB6yHI1
CJkLCHq+RVA900T8jvv6zVJsl7nnSnJEB7Xf2jSSe0BWCPGybbTVahkLOWVhtyvu
j7bgsFbBqUYlgBvzxUm4EeAa482LOHFVtdJLAIGbPZfV4+7CyMPMTof6twxbhfJg
Cw2ss4b2MII8E7z5Av0Me+odx3zNe1pzRH+q6Bq6GxIfeclIa0Ike68ab0WJKqS6
TbXYUdX9BgMryrxi3I/H+z30xblPYjJnKRoJGzgSPgXjPJvxSeZG1dsjdandOvkh
YHeUBhBMMr5muwGqj26drHEg/UO//ietWPephD5IIlU34UWfxBozr/0yA+iHQ+zn
+SwcO3gr4EN9CXCaTfMDMGhtcafQWlE5UDHIrZcGUfteqKTgO3xImUtfYZSsxCik
GoF1woUcFW/t1AUZhBbCX4aOZtahyWbi9xr+H1FpvEMqRPqINs+7KGiqC+RFy7oh
hcQEaD/7qdP7+jmROTQbUv3QoZ213zR/sFssUEVnvBE0CrJoj5hPJxq5qKGf58+1
WUy5K5hijyXd1EkAzaDuHWekmlDeAy6uTROBzjdecXHtXwzpzfbWd83UUESIObAC
88Rl4b/OtXDiKQbxe7WREpLPtCmzgRI7xpOhAHvkWUWBzpbFxdmWVBmJ+3HDh7Ug
u0npOXS1SwpkkJS+rs5yWO0XCfzw+VJzNN3UdwO4+aSU7o6BOl6/pdy9eNMd3j0+
1LHDSTYkvvwtD7sUYA82maF7F2YQi0FFwESn0vD5dI/mXWkuaDuO/MvCNp+mo7yT
sTnZDN0EH7C/+B5I8W0ZvoZy0Q5Ui5KMegBfcHwemO5r5IYUyw5DrFUr8hz8e6sr
6LY2kvCGcygwDISIbIR/AU9LonVqbTTOkbYWjNg44PnA8UIGcN9dLVuDkoSOj7kN
vgIQIqxa9NmfzB6OiDyiytIl3MCVNQDKPm9QYs5XL/aPWbdA5gBhyjoERYZVCgD/
rwvjA31RKVPa4Q7iHjbbnzhteD9azsGsrlEZiBNifr76rQkb11SWvaKzQxcZS5xz
OkeZ136ii4oFjReNPaoVNTQs7nyCEbxRKgi+Ql6yBStdBoQ13GqsEUU+UXl5Dt/O
62IiRV9fTxBNhWHUxp84nlK1leZzhiowlWvsnarQ9Fa0/t2wW8CBB0NDwMQqBAht
th0RtSJpZiiEQwBC9VErXGhPIHkhKHPNgvXL3MkMvZwzTz1xdOMmVBZxjVSHSKE0
ToppK3VRWXu69lCfCa5AC84y0K0fVMAqHdh8jS83NM5jSwLvk2sZsF0kdGr1zJm9
YtcZAWu0gHSbIMuJzK8u06hxVbdzdhoIbSWJOWl7F0urMNcYuDxDKztqc1V7rEps
LNBda+nCaQ+aBmradrwVHqhMtFcJPFPE5GfK6TB58dIFWVDiu+QxdP/ks2d0nXwD
1cYDVZIrJAwLQR9DVkbAdiL6YPacdqYl8PGxisn8QzHLiZ6S+0bMt14G5/cKI+UW
pcRrRlmQTJ9vhSV8skhT/G10LBtsgY0JHN7u/eIt/i8LeJ7DOxWk09l5qkn8CubW
jQfBWE9rJNKdUyiOXxcmKFBWTQ2/k8XJhoPveDmAvVlRiKqi++Qz7ZUQsxc2jWPj
n2qn2HSuxsPBzBjxXui1dUSdSlJQv1lzeyxyzCGxdOmLlxJG/dL24X41NLOvsqqQ
YUQEc9DWOFy54YQPjKg9dqSZX7aZe0JKVkkGszT00kb8UOJMYBc/Gcas+4sMe49F
onIEmjXs7U7Yf9tGqxhzD2TRcD6lskYGLx7sXFk4I95DJtn6svt2dXsH5tW6/iI3
pR9974ccQKrv+QwSF0zv02X88VJADQEZe5LEuSTBuTVFaZAyRULDA+QwdxQ2rRYB
JCY3xci96/xii+Qmgf6UUlHpgrd2iKcWkubcZlJnDxNuU5mhZTISx543mOaOAnPo
fcNI/42ku8FbqYvYGHeZS/1csVdMZbt5VPbN4clMQR4SmE3RRRNac2tfwv++XgwL
pC9F5XuKUdveWEhN4sw0/gf+Uf6Akr39sJvvdvzF0HrDk/NUS1vZLplU7YW7IeJ2
N9rAN8z2y9+bFxELT/iaGBXcCkPGvAzn1eIpYUssv0bHuzZkWsheI6CH0fN7rsqo
JxxpExHtxz6/qhpf/gr0SYVP2ftcJvI4m6InOcIZ6vnX6CN5v2OVZkiCTwu8AlIz
hb213tevkcjZV04sCQxO+sDS0hF2xCKgWY1SOEuXOZVbjMyZyWqKLAG3QjwkPXRl
MroOvazWLXwF/aBBp2mCu8SKgd0TemPnSmV3yVAx8qI8ebRv6ZumWaqbKtCx+EIy
BtYc4f4llIgHplMULuAlCwaxI5aSH2qq5XPDSYpGiDke8OwuUTW7zGDgTzFMI+DK
AgiMfxytYLbXloVDffe2487B70XK3WaoYOtN9ej51XHZnrl6lQs/FINlz56MSgh/
zF0WPQ0HsGFyh+86TwG003aJ8Xn3gUMFVBwYtwxuDAZ+ILyzwgj84pI4fEBZJINH
s1GkHUIflb637WFs9sl8Ft6TiShUM9BDi+jAIUrgzxi95ZUkog3DdS13fq/B4/FH
EIomrZJdJDV8tALHmQlkftFT1JeLjPyfkmRQw2aFh9vZ4nYx0B1RZ23JlpfaE2nB
ztHJFgAuxUuZAVn4SuYJ/H8a5iDhuPrnlEaEC/ljYWcl3GCwtGZ6qg7/Wcc5xiX0
gqg9T7BHXMTAciyzvqkG6zHq+P8qqu34DM2YqSXIftVhXJzPJMhlQ29m+XI5J+jE
HQAxYaPNcAMP9V6IcN01IzC9ymKSCa31fGPv2+9++T+DSONI8MruwpVwM9kPremW
n3M8GSSuzcNbdNZNO2C+70G6arSkd2XmNZXI6vfmei6193mM3KY+VWL/yAjm9P3g
i2lW0a08P2Gaqvu8zdzZR+IuDvU156icQwsgPkuxhlPMHJ3R+XU3npm5tFfDO3dq
KhNps+WKh0GFhqgBKNXXphyWo4Lo19VgKTZZnkTnJ02BSwkyxooC79FN33u1QEPy
CKZD59PdIsHgAzjrybdVYDQIiiNY7mxa89YLivzNtVxk55LDwV8q3XM29/iho84L
PYbBmd5MGSL/cc6rwq3k+eM5Hnmun/H+5CQD6ON2r8f5Mp/U3Y6FMZPafAwZtXtO
JT2Y26ZdnpghEekr+i0bvxNjKV7zce3D6znPn+15oX4IxkaNK/vEt8hXcJUIdkio
Ah6uda3DryNopAgZo8++SBnH8gUH+TyEtWoPr8ut1pefKyEdTI3blIvxF+CMqKnn
NvnNmHWOOIw7hsetBWzm35STFAtCXHbvenW2uFUOFAmymXDX3vJibSGEQw6B0qVJ
uUMmKCxz1RLs08JVPBAg783Yg1GCfNRAmDVkzNKq27vtJ0a54H6qbjElFgEvEqpW
xUt9Nsf0ze0dQkRjnHcpzCpuzTkgQXE6nCJWvn5vU52zniZfPRkTcKk+5bak3oE6
WX+1TUB5kbJhYPFFECr20nMCR91u63IIlg3/ce1ARqe1foTw5WbaRXZuttk+2X+5
mTJiJE52kfoUdjtybUxKbk9rDlZufTdLfE4Od4pkDfSbBUBU5nhlnKtccbLURf6N
kN++8VvjlealUrhfmg2VNTDgRBCjgHYmQq2wp5hChu6HZJXdHvpCO8vGCjR6FHSu
aBmRc3frXdZfBjeVvIA+OPeiL6IcJNc38B3aj3GB9k5NoSWPwkWZSWDejHN7NUPV
gekVGaN1qn9Q0PQkmZhZR/wBobCgRx/iwhzfhTherwGmkIcdvgfny8lJ6G/whDPA
HsbXJipKuThhIWyADY26UIHdiMpvxYYXbIZpzhQ+8XNuFB+GSVEBD8sNejIJQntY
iL/xs4XT6zUwucKcK4VGy5LMS72uknB+1SV5dA5unpVjjUVMSmO9bPD2VcdiMigP
engvvPQdBSKYzSZ61bmwX4WouIZcI8JHu7O0MA3OF3ZsAeE7YWF2uXpIhagkvlpl
Lb1El1nWruCzum1WHvFBciu517q6JaWVGKSiUS2vt6b0gxcwQ/2rduAdCL/d8N2U
ms6qOaviJuU4uT8EXKyAbdpQk1fMwVPPXjS3k/Cskkv54e7peV3NfPNQqMfJfvLy
1xRi06RRSW63X0D/1Dv6+LnBXPYJWhzpDczT/8LdepWK/sBwuGRJ3FQBabBPwars
a41XwWOWSb9k6Jvm6IdUocudTLILcaqV9DPSl2mFkvo9yQNsCtLDXsjjqVRs8Yde
Ms1GarJSbVsrYYD13+wSRc9rcnFSfVr5l8e/OPyJ9iAin0smo2ErmdmzQQVZ0aMQ
a2Oh/pX0CMfILuVrD9R6bYIXIZAQ/Uti9dr1OXUcO5v45vZt8vCxC6BvWN1+KSAo
klqW0WThXwPC0mhpGZZWs3N14d0ILM+NdBqO/ZfubupZh5RPNlpfahd3zvapWpV3
sef1IczVbqkBWN9pk6dDxa269coa4sognyI6F7Btsjc8Cbt0ZZ6fG1us96CKD4Kl
IvqDwXY76PiJa4qeiG1n0+d7JY9EXlZqEQTfp/meEryettERuCWs7NGEOPEq6gUP
DfrqKMp6mVeQ9WduSpVsMvApSXdwPH6xBfXrPrsyj2r7smHJqI1ebPx9LsxXzw3x
b53meJzO+On8h19yKYEa3ajBF5zFu0st0kWyH/9GHo9WooV1C0LI68w/hQ98EVff
Mq7pNda29i/YtZRKRg2oGcadld03umhgc76OgK1LsXwLBdFW9m/AFPnRi5BPDxYx
s5Zgy8yHyifurowAy6//CLYR9Ys2zD10adweZYOHcHkB6OKCwa6eLdZiAugCLgre
XpL430toDxqpFiOLNaNig9dfP6IiXg6YbmCSXMR5WxwWfkVjqWjVQmd/sQmY4r6M
m4tS/rQ5QslOa61vjci55o+cbbOW5tsTp5dZjbzvMtjzWcGN7ZLi+Vb9nU/wNZY9
Nd2YQ4Joe+q/97aomhRbH0WKXbl6C5GPCUWNqE8pMHSenN/YEM444FCfTWYpUQmu
wkTjicuz5aKVnnfCEKOnimB/FgnypoWcEzt1h9Esg3ZYdc4LKPRCrNra29VXFdlh
W/+KZbz6n2XOQM7/AbsDwAhQxD97iJ1AYIkK7wP1kgjh6404NCULWVY1wsUxGPQa
x+s+nIulp7b0L8MwJ9O6SiBB2cHialoQ/rVQE6EWZTiUSKDntAXYHtgrnuUF7cJ4
cuw1OHRM3ZcXIH81eRYm1yi26saBHVjb25EFkPfmc72mC5Avye1XJsk+LClhRoUi
fUshZm6b6YGSsxgQ26lTCL3hv3js+GXxmR1AkPBKE5VCRWCN1G6LtlF4ppkMWe94
+C390oBOzjSypCDLTuSoMROpqcceTuKjk/Kj1+7gphb/QvA4vNtg+/K3BGvb4rWX
OeOZ1pE5yqoUujw0gf3dyoIaI83CDb4oVkGHQ515Vw+jhlGA4LNxwavUdHmchER4
9zC5dHSE5zVG2IiEHM0Zt6hy+42rEI3mXVn8/vnW+DeYBX+N7F1N4AHU/lwGOvYV
8/oU9Z94K2y8HBGVmh1OQ12D590aKkEgmDCX9IH4jpBfOVrgKKE75LMlXlOYMIYF
rC1L/b8W2DNBcUY8lWgnKIUq4qmjqLCk2g27L8gufXPVzPg8TqQrjhLqkm4gXGGJ
tDSGZq9PLq+x/QJcpNOnJqPWjSUWeiZLdS027+eNIyndo+ExAZLFjiAotTho9fX9
UrSVlGfukrkYrDBkxKU5rHXqo/neQofcQTLDK1ehUk81bfnMHIbrJm0YV+MH2C+M
3P6ukLKwn2AzQsUaSN4zD9U4lVx4CAkbnRhbeUiY7B1byga/d1Rr8maAx1fC41Wz
+hzYLJl4su78TiiHzmzfz8C5KPP0V5/EqCS9XoiCmTOokIlIOHo7CcMX2KLBTapJ
1MsUFB3ClexxWF5XCos7A0rNOEpfnFexukJc8uu8xaSByEIg/s0XgnBPSvXcyEE5
HK1B42IIUVlotHeozVnlroboHIvLDjTDcAelsRoK+2OcvltyzmZuNSbVzV2tME4e
cH9Q9NZPEm+4nF3DpJBvAfjwCb6OE8YjK8CvbeDO5bHhIOUOSjaiLQMqluGVS2sw
ZcoW8b5NUEVaY0H6DYNrgA2I02m/E0yjxQWeQjOp3TsYfYvaRu+X/biU3HI/er1B
8ibzWq9GOxlHijG95ZNzBIzlNRIHRXGuJVL2q8zxlT4GcuPb5Sas7Mb+BGfUKCOU
51LdBOpIZtWIPA51yS8nGVkN4b6GxHOgpPrdvLxHR+yQERHQpwh66Be6s+sNlCPD
fLt4FcHemNK8w4/WGXotRM8WpiwKOa/a8Y/LdzhiWLmkQDEH0dy31owoDFUPDm8L
oLw+zLbzUQfPIUb51Fvu1VslQqy09GLU1I4OkGWOOGxxH/oFzwZ0c2n/Nb2tgySB
2nFx+gk/tdIYYT6l0lcL2ZulCNc3eROOXe/Tw9h4e1wR8OxMLPBDCBqlzRMg4syH
lMo6TOiDxoak4oYgjWS7mDt73QMSGfSLRQCXThqhB5YbhV6B+M4qMuQNs6JAvS2z
3NZ1+lHqRIPWZhyHGniJKWh5XstIgjUg5K2bXjsicSO9V0LPFnA5z+N6+2qDJLue
fFuGIw7mW0Y+JFyZgWMK3yIpKXmD+LAQnWJlOLEhofCglVD1Lft3nxwnouHrLGl+
k1AzBQuOFrmNjnCtOoex5Reh12K+8ChWyD6ASBdLPYva5IHTPQbJi/wMrtrXE7jT
AW7ka6sEMSr2dkmYcQK6Rx1gW2hMigEtr3B7RZWyaod0hVVk18nC5yaXBZHF5IGw
HlXLL9HG7q4jTyPm/UFrEOutReoamvdQaOJOQCbOZdqHMs1G5iuPGyjBeiNvm086
ra/otkvheZETaQx4lMnl8aSq1t267Sn3E0doxIBNkcM0eHgnLNyQKQ6U2vLcjAFW
41cY6/xewFS5UCM4FTJEuT+TQS1DbMNttiBh9vKmOaWKA5f6DffBqEmHhKddmvOl
oeGwHgG6gW7D0fdBd1hkGR9VpLzDTu+fgXg1R4HUNsdO8AMA6iZ/hszb37NMiQDf
qvlwEbnq534VGAkN/LIbP+nNpVlTa/LWIcyTpEXtvfsMoDebVG0h6wLFJbcP4DS2
O96R9t1YII/QeKCJ1Xy5tz+djYEec3mU/kS/PdCupHK+mnVNtKqDYkU70CHFXHEQ
amJ7M4Pxpvf0pNQbSQkjJLsfuIid5mPvrU0ksHXgOgo56x0q8tQAsSrLomJs74SH
tCKQLohNR+fI5WfNUDBfSwVLSBV4ZEUIOdUwhTN+QXEs9ZXmmsyg13tmVvim2IrT
zGDAP/XeskIKk6wd28OwnnhdiJS0DH6ZNuY7bjolehX+p7GgrY0mHL6KEMSUWRBH
qEGEM5SANju19mSQ7seE4OOVXoHoAmKAXdNTv4Pf7K4ezAxoecPZZzoYoZ8XTInh
z2KSPuOVMY7Lxj4Zyi0mOy4SlfBr1x7vLQitGMM9TR0uHoXbexmhOpDs5eZeL2hX
r+cOkkvEYddYKau0hT+lX75iyJwrJXAg7OQEqQiTsBWUtVzh4BdWI0X8lkntSVjD
toZejfa9uTRJXFiu6zvo5hvqaopGYY+OMixijhkwDJ5Mbl93dz2vXERNl6WqObHK
ccPxRfmMarYA/BP+4Q05MZqBu2jTRNj8KOf0bJxJQVi7pzu4rHB+x/x1PanVMGjF
FqQ6VC8YY9SEJh7kMury2Wfs63cd8fCAt9f8R7Kh9EDEV1r6nf6UzIjJP2yFuBSN
T91MOGB2xlXRt115WYr5z8AZmuTeYoDMXxgliNFyt6wD022WnLXHxO7cXznCwL6x
cI+TplXF2JpkQnJbKosgmBOuC3mlfuBRGC+AVwLICmtxIkvRYbTzTj6eoDOoefwh
8rPxZx6qfcW+HsPUDQVfzZl9UwsETd5dP0u2mOrtiUEm7hu2WCLXO2z2ZVBZ3X8S
BOHaUr6QPcOgDl9KSQtsTXQqkgsggcTEkIqHzwaqOpYQTBN9d4Fn+c8S7IcmnwVD
O4HuApit4g3XVLrHVYA5exj+pVf1vx2C+k6bK7M/9Q2DgXIv8QEIa4xDmcZj34KI
/IlcW0eR8Qujv3UmxWwdoZAjrAXD3GTsRNfRmHdiJAkRX+l/iBS3IFTSeNLiiIKz
jsO4wwKkzJiqjETpHC3aVqS0UFMNFuXc0kfci4XovX+uEfL5KrC2XaK05P04Ibu0
W0/Z1eX0xslk7cLWHIZOkXPldNExmQH7O4TfQyVkaOvq/lEsI2QAkHNp9+CqUi0J
iRPqpkXLwNCnTe1pSRT1AV28/uXEFNIURVsHzW6Cdn7pzk23BJzjnMvPfkN/OncC
DzoXVpFsHNbvdL3lOEQlddDRyIf3M+K8CE/iMYl1iacgjBkM5rZuGZcXlFl52U6M
OXfD4bTIZt0SCPGG6jWjjpunpkLc84bgL7TeEcI3lc+X4LQEFwqZZ+0HagbbRSYH
gpYkHWBsVZ2Gi8XEX45RyK8mnypruOQccDRjlQTW1zl9hLTY567IJOGUPxQhnE5V
1UWqApdIGb8sQYZJbtW3GHjW8500mUf3CITxVr6fHuP7TNCTfYjuun+ms5vcHfs1
INz4WP4tGL7XxHzu0QixjwIJtn8C9X5DiGYVPmD1SQX92ca1QIP19Q68RKOdbm9k
a70yQy+BFNDZnETOH4jjJhS8X1+SQGwYrCREbSce+9cCYNzTYJX6z9hseg3ZNhrL
Z7/WrkKUgLAdEDxftvMkVA7fMPiW1/swOHEiX/Fnn2k0auSpY8/Snq/mUb49/Pex
5GfFLB8WtUu0zvTDDMoheGVb67ZvLhyRYLAhcadTTu5nCvPlKf7czkdWLFKxYVLu
WPqnqeT2pI2Gx5NrKlmaU7IsHI+OTpRvyI8It63GvVQD5BFtvlVRpLnKGx9czgLK
34IfPYkVOnDB13FT3VAYuEaq6CcaQNP5G/q/D15pcbPR+ikTCNScRBOga5I/swQF
ipiBhfZDGflm6sepY9uI6rlIAqkvcv0oe75TWum8UQ/lxFXS5rFScHagoyx67U32
d5CCJQImHljbnhzPLRaGZ/OajFHhDXnBfq4iYRwA3qaPD/p94Gcm4or1zaoPm36z
haKbZm/NvrFo6OhLiKqF9Bc9WQSxdR0d7UNYrcBUOxeUxU7ppjG60M+H/SD2Z1BY
517S9RtFUSuuAGitz47ygyQdrUEdASc5OvBVLTeLD2dm1KWRgVEFzKAPceND4bh1
qREMi1be3PrduNjXEjk31v3/AMTjml1tqIz/QKtM5wKE5M9uicQj6eQiR8cbcSSg
lKuVc9ZGB2f2omaTrgm0TgzuaG6zG9kXeZr+Dt66iGakVSJ8RPb7ldnsGPtJ92JN
kLP1f87QlJamuSTqSKIklnuqXvqej3luRXgDEQw6ZliKz/CuRYNECWdvsuzyecfa
5nuHd75gNGYA3FbI+y17LxPN7K41ITnhvatYSueTdvou87YIsg2hOy6h5VSqQrKT
pxPawcVWxOjRIsGhdmGRQjHosYN7T8LhLZ6boBPqqf2F0uqh4MYDOAYYtip+UTaA
4n8jUky7T0O5te51p/pFm4V15llCOz5bBArCw53pzDYjeMkobd4z0ZNRY8FPn593
z5mglrvrrreFvYGy/3CIP7nJZyUKjWucC9vH4iPe8jqsGtMuUu3qcWS6mTeIVLIO
95JiTZcDSRUZQISgEXG2LyDWG/TgFbPJ2u1p/PIKfeLqWjkNmQPU0YlcIet8NIlD
HzQ5ES9fSp1Ps0apo4GHvd4FZLg6r5WiiYSAlp7HqJ8vsxJ3pJtOJj1AbxIRA6VM
Xd3VlaFj2Mn8fKBwOZrj4HD/VD8l0ZLT2uSi8DuIZiUQueCDc1SJxlrSN/W3p8hm
zqs5Ej/ceQ0wjUJK9KaldbtmD2I1o57D+qbJutexwO/bGovdaVjTcvPysiFsJzVL
Gnn/oA99iXOxDRtE7WZhCLhv9ewEWSUcXhHGJQq+j2WKGhOHXuiIetGtjlZiXQer
u0fTFzj1yzC5PdHarluXlvWB4gx9z9zHMDErEvhXSjp7nyHblyfAt28iiIvPRdIx
el3CA55A6xDBRJePtV38qLfCi6wgYtsRRuZDMB2UD+oq5hc2pSIXzIaHhuWvOb+t
LEppihGT1t4GzNiqLUm5QCajqsEKQskkOcuyzduyHd2Mc6Rq3hrwgt5K6B8m9+2U
n0jmLeeEDGrvl1LrBufLezU5va3q8N8TUTE4UX/O4CLkKRvzH7fa45SO5Dj4T4bo
YMWH4kR77+S/4Gwdk8tAp/8zzq41OJ+1DxgQUfb+wqtfyTv9hSB9stuxLIfml2nq
6t1SGLLfD3CCN5pjZz0dI8YUcg5QXgzFM51l0Pr9TY4mHr2bZ30+BODDX1Qag7lj
6ndPtZqfMAPaGMIyK7ZMFKa5QXwJx66Aw7q0fUEP3MB7XE1IJTPdftXPxeFuABcK
n14NFP+QV2sYDSab52wiM+EoQzuwykATxFVghOuaPylQfvfQP6V7uGpm4KX9yWV6
FEU5UKMmnaoSBFMhfnR54LOA4u2agFYFB+iJPzRvWmtJ2bxXR3unxv1K8GeL4+CX
vLoIlfgnnQmVA3FhW0a8lWERSDO0lluIxqjK8yaSQfBdgwQH9DVMMzewYHXQ6M9e
jg/tmN+t+sGiXIXHBSzJJPmlR+gHZKChy+qTM3WWxahOFJEHA+g2PvNEjFQ6O3Qo
ETPxDMcpwr5V+5FpwEJW5J8Fv69q5rVTvSq5HGZBB9eUGj9Xz2aynUADhe+AQRl/
c6OrZGnZwBc4TSriERe5dhATLoj0GTgmP5Ad0BbM2RQQarTOuv4KAacjeVBGoAFp
BNfoixM1aV43WMn8UbO4LWjuAiQbWHrnWJ8yo4yh8sanRlPSKuQugpFTNjJzmmcU
EaXWzs6YzatYtjQPUKsrsHnqA+175YMAHOK5YnCkc73BCjGCP6XuUIdQYPRtmHiN
EOSVnjiRlaAK85FHuRAF8aN0TIhoSlLwE3NMA9q26nM/TEnU6AAUp+7IT5dulnl6
4UEX7FMOPyPZuTodLM29FFykWzAySDEzkFtw0sDarGOaZ0tNBMbvkiaiwvmUq8uW
tkzPoXmKoaEL1XYA4z4Fy0pigeopvF4nHh4mRPJ+EbO30OWIkZBJD7wSPAtzPhPG
WhiRy3UIZbvXwD477UDaSyJg0pnk08oliaZXajuSaHyDiCooVT6H7nIRYvSn4s05
r4FopaNPlNIeA5Lsj3bL6lDWxN8fluTEfPEpsWq5CD7kSfUK7pUn1rY7Fq2vQqze
t04kHVNzJumuihiykSfbg3OrZha31yH2Bygz/INxrT4s2fw0BpcM5rG0pcs1ZNhq
087S/RWe+TYLvE0LGn5qqyO1PAGlWDqbkHJkDq8ABcNnYgDn65k8bkHVqiqBsDwc
Q1ymkezMX2LZ1G/WdO+YP8nNFaNSs5ZWcZlegB3RIMJXbWXh/cbjcos0sEbA1r7/
9Nws2PJyQXF3pzd2eQ848vGzoDVt4Rwkx/60hq5xyQ54HVfMupIttQJ43aoy5T5m
d9Gkxb0uNSd24LFfBJqRDzNOk+ENVQMyIK2GtbEmtbG00vunARUsMEVHtkaA4fsD
FLR2PbO7KIi8m45XVPaIw0xBv3HPVmP3baobEvsVI+1lnJZi/2MD6lu+PwxL6/fi
g5cYJ+6G8z1T7fPc95uT4QJJUuUsVZ4PfVuaWHszPV0q0v5NQ5zmUg4M59q0XbXD
SooiWuKz2YimnQaiFAXO/5tD0H0G6BNC6dvVVzbylv5xEZYCz240MeZZUsswuMRf
xpb+Szy1n5c3kWlC9DRfxtWDA0FW1DB74eLYIZLDdBKjMHVsAcuTu6Yqv4Wq4fK+
Gz9Lb2fH/WHrs6LNEpfPxM584KJjhYXQ9dhe+IdmUzfHo30YkQ4EvdEuibNOih1x
/cbHSZffhLlgRUKO/GYm3jw5Y5qygmfdi0akINhsKS47HqU0WSQO4Ghgf+8YQ4IU
S9l4T0pUDkb9NP4ub3fu0BvFyaacoe7ihQI+EW/W3VYovW+oaIG7e0hwUjXlG3pE
iNL9lvfvz6ktosxwpLGuJfYPOc+Lk5qe7hPuaSwrsct+9unHYtzeccognB0Z2f30
MAoh23cOXYZJip1ZRBXp3mZbeo7WTXMmzuRYDNpkyoOmQlnWR/UuYSZKOdgrvM2r
BEa+DNChSSGWMizrTseKCfH+w3YFFiC0fvh0Wr5VBbfiKBBbyDzwP7Smaw1S+QY3
QL5CdNpZ8W+AncMWT2I3lldHHaebQT+Ix4aLoVrcWufX2v/bxL2oUD8hFHG68AmX
oejLNOx0ofq9vp7NGALuTDfNqaV+pfIvkTrnhZXkhDSbt/9aqGPU4YcOZGVgBL8d
AV3KlXGEWyWuXQFl6PSzGHvJvaphNu0MeU2KUgG6KLTI0/2YhKmlnxM911A6nTvx
yg1XtJfi8KN3fdeTqoJ/9fsJKspuBo9UfBjmOYHqsrqiJisDScqjw9ADCq+Let4B
d4cM435gR0ZHj/cXlGKPP4BqUu1rQ6HywxM++FUtrcGmvSMwVIQsxkDIrvAPi+Gu
QdeVavdWx2Prw0lHjjZHkjI+LozIe5kuENJUUWnF3Mhqhcczjx28wjSu5d9HLDUD
2p1pJMAhrQtEUe0Hml6F+mfJW03trUaRL2svIFQy+yO4UVxhYAW45GsDe6D2WGOQ
yd5oyCDUUMXVAEkv824IG2LCgUPjY0vJFilJlXtVlj3zbntlfh1x+n3YvSWC8sM7
+UXbbm3irCWiXLCA2CZhMeu9Ukz2GiYyq4jYblL4ZVQZbwHPaqKfMTcWa2TS8vJW
rL9bn/yEKsTWQUXQjdhZ1Wz9MSHSFPj54FZGJ/75ozxfu2A8eOT6RRZRH8yAC5aa
OU15wqZYxd1vCJbcaoUjD8u72j41BXI4t4Mq2kyDkHcUFrxcB45jW9fviyvVEiSa
Ut5NqRVcQGAJdTjvZHYqq2Fn45VbbM7WAaLhzuvgnMUuK+fqmphc7FV/lktL0Gmj
KJhl6Wct5xH5lxS0mKuZu8FZ0xu6hF8WPN6ADX5Zb4JYyMDBbs7LH1Hy0jr6PxnF
wPDGS4Kybhbm5wtJADzmf2gNAJMiZCyrmO0CUPHPAcrYENkm+k9QNd2/2owFjTav
A4lff67dyiA0676e5c4F4tF/u1hEZjiGd38KzKPgcdyx2Ba+xvR3cP5IDkYwvwD6
Iv+GjmkJ8AVT5+A/nUIqacNtcuaEM2yShI9MO23DBLvcBgi+uMzQh16KuU/LD7IO
+WAINYnDu5bN91CRPvRqG/4Opqdl/k0wHw0qu6ppLMyBK4WaLF4LElrMfAoOSVG/
m1t4xmT6MSIMHXEyJM8wMVf+ICTZRnCQKIkYtOSv/T80AKiQwa/pz50d1itgZqoB
tZzaou4fdC+9v+QBMCgG179LyNPGdG8pgMwXP4+Se60kl1izq9CYDmOpr8NCXurg
EupIW+Hn4WMbP1LrDdp5Shb+3j7uxzg1HzvzUe1D1YiIG3dxPw1Ra7syyejX0HAE
OB1jDfQSqIlXHSJ+GFklQ1uVsrSZACPc2CNo+R7LSGliXfM1NRNQ0lZEZh8HBmli
bmCmDj3+unOllF1xsiMiDiRr01HgIyDWPID37oHRp0KVPvT0fa3TCiTpO+Wjk08v
bkH+pH6mHT0DNNZZkcVEnhvOyvTr3nc85LwEhnFO8vpda6EQT+sqnpe79caIGe6W
HhRt1tOxsmoXRNfZMoJssIaT3k42zwTd4lDTP1JiLoX3ohiKACcjAfb6cGLToymJ
GvRV5d6llHb1N1oB8o0a4ov+MUqlQas+Clda4ic9c9Ii7mpNPM/j0q5LJToiJYrg
XVpsEpiOABMG9fvnPCJrV9qnw95rOm5I3/EJDuFPWTvH+tcKwtvmxrO+P4s53Nrq
FVVq6Vvzdq/4geXMdsuNnA58+RIB1AHz6S0RMp3HeAkdjM2MAL0xkVBlA9QynS5m
foGdl1mpmLqL4S4KZIIKpj/ZfnklcGD8am7Y73/Ol0/qqMhxfIyll38VIbAUsu25
g5XX2OzlnWKcIZ67hlLv5CW46daA8ISdkosqemuSZ0BLhJ4LBZtcTdW5RgxWtDEm
MiGnAofsSgBa/Q3XWS/pL4tp/05pi+0yT8S8KI6polYuyGxNzMgNPxDFPwHCMRR+
HZ7sJjcXiV3ejJeVnupFc2AXpCNIwoY+rAZPE9arFHPMvwHOKQVAUSjTWNETLna5
agJI7SJo/1sBTgwGRaJyi9IBTITToQhkU/AE+oJkw5/XObk7nopLeindK++DgRDc
QxqT/172i8xOdm+R9qHM6gGUc1oO+Iroi6rqFggvndGC/lLCWGYrAyCr9TvcuojW
YoqzaZN/YJfmduHNHay7lRyKGA/32MKnydlybktLB/98OzqkXNt5Fq1wbSJBpRaT
8jjmRw8c6S9LO4xaqY06mFIAIUTlSLajL/yyE0rkyyp27xfeYTElRLb9vx0oucEN
jV/P5N5PfpZwROsXKSfaxblZQPXTx5bcdWufGkg/mPawWarv5xvc6+C5zZfnzqgc
+xKQ5xpbwsUNK11B/0RCmb5uVhXup0931JI/ubAG0GhmCO8GNmHw39vstUIU61Ev
PQk7v0seubnt7mgYqE68HaWPWYpJD6IUU8A9Yqc8PiUJftqzftoI/bAisgnGiVfS
SuHV4pGx5Ij2vlp/v/8cRMEgunQdRbob92gUIjnqBmM0aG94oWfvhY5SobSOzQmd
LpcyOwfgtcUgoNEFgEmDfIV7zK5azAC3arTDfE8JJBRa77Z2DDVm5dQpT41I02O7
HXAaYzjVuKlxtcehgT4zTJrnFKlhjbFiDZuDfyy3yn6qeanqCx7sTimimssB3mj5
yYKLfXY8aWu8aWrqDHnE715NgUnwZQsruVa1PqEoxelRQRtZoUehRGqdurKLVutL
8EG+4uHjlNtVgKjuc2UZSoM6jIGEFtkeTCRCZf+GL/JAnI8vRlXmPXgBep34x7NA
f7e9UXaHYOADsk7lu7AaI9i2muU/SxDNDvQCDeJX6x3/XuATyzd6AaERe/7j3kLW
hGqs/3kVmA/Pnwdbv2UANBoP+9eQmEZwtpuAjFzMyBfIx2z7yCaRl3xh/prdxV9+
WgSHeOXj1gw6Hg89Q9s0Dn0vsn4NgIbmMsS9mmlwEL6Tn8OefOnYuuq6tExG7vTi
BIMmBVGIG4efqKc0Wtdwi0x23dRtIg/0XMKUTD9fHn+0z3xiOxxsqyFPVEg6T+MV
cVhpPtxNoWpAjLhNj4ngF+nAHn+Vs8109J2dWj6JwxwwIYa132D4OrHcMCR2ix/1
327XKVpmwbfFy0/3cvw54rit8MmO7FCmrPARPGxuI59C9CZAUhuJAgk8cF+xRE10
uh5pyo2u/8lZEvgkAb4EudotqAS04kFEp4W25awob7nXRRxVqR17UOaVCbuwqkpg
eXQ3GTjAU2lh8lrePtnF+oy87vB0sbYHmWQXVpw8xL+KCvv+xld45FwNNYg2BEfA
g8hkl270st3nGTE9vOyfJ6nD8kdLnQpzCHYTyrZS5Y3HQWIN6iyoK6NCnbpJ0XTd
38n30T3G05oFN/FPkha9jpIpJoM8lu4Wl45/0ekFoBJv9nZXW0vP7exQZ5tk87uJ
btOnvImVnFCUlH8RIZeWgH0a4ys2tDJAAEdkAiW7Y8rTJLoODNPfwZXPcFSH+Zdt
+JjZt/4IR3VeaxxSI3IQx0fiqAq1RaEt+rxYGp4qugi0yJTKMgEQPTr62g6Ehz4N
xJf23moDcJxjFEL38LhoKfMe65Umlor2EekP0StxR8+H5MVIPgl99HHbnwGhv+Mk
4m5qxeKskDeRZ/qMCvmgXmVbmWhtekJYiF2BOFzoto19X2J4no5+y2hlw6GxTQyo
1+b2U82SbHfAnCMEJBVkOcptvsgzY6a212JT46psvIfkUDQwut4dsJ87RorxTaNn
ZY3geWIo1ee70FnjY7EmYsu6f81ZAOn46W7P2ge2DYT66woh4bHc1lmnQHHJmoQj
55T82oA/PEJOGaTEUPE26fbvER0k5db7vGbt2ZT4qkxMa5WkjWoQA4hRRCU7gLBm
oO6L5+kt9UGHD2GeM9WFF4uiKq4YMJVLFf7PcI8NAJqtsfeidpedjnizr7JxTQrL
4HzaOf8CesvWIyH9CEPe3Pw+PLgW0U5ulD4idn4BGkMN6gJOHr7pRoYqDRD+snDF
7M2qXxHpTXFkJuLCq0sttaKchkiygYJ639aLZXdqXKB+a/871FbA2emVvWs3N5sj
3PsIYjWkMQ0wHlksZ5B3qgJ60Y7kZ13myTjqS2P3TiF1dKSF95QvHVWYPotKa7e2
6zVSFwcfbA5PZF5hpNIcyderXIY/qW6WqKooyj9nWi3Krje9JeUXZwOCv8M9M8PN
EDvJp4zYvsQ9XeG2dcFIFPrU1kkWkl76w86IJrtQC4OYQ7eE7SMPbOL86csSVnzZ
dMDZXvvDlqSm0OdywQuq7oOqbxOFrcfcJ+Y8FwoKL3eGllqJHj3Hzjs/AFE4vsEp
rN9kZQ14l89sFI6H85yRnLBCJJ1wrERIiXHx9ZFECjPxso1Fdz8as5i0BQT6IJZV
+ki5qr9tAdxQ6aEBu2xs4O+nL7rhDZzCNR1CZ/24OOgzl3GHz5ObMO1Bjv0g1rfk
5u/lYQ48YqfylY9c7BYK1DW2eV5N4lMup0KeSkmtfNSt5oiijR4K8YDnkh54Xhk4
xzPh15m0oSsO4+zupE3RHm2FjhWDZ/Ss4EYhAdUwpL9vMFmmfvShkvus9B7L/Bfp
s7WF1e9rj2UHtqCCLkFTnqqkHCZacAk7b/N9YpPuU8UHITFbfTIk76rtEVNJdjj8
chZEPTsdsWRZi43UmVSalCcZAxGTQGr+t/RPtyjOAGkM/hniAhm3k428SYKg41G8
DzFbNzbiDjOvpvklFppOwvNdFjmEGZGJdQyYcZAJQbfo9Ju4bFvQ/rxNtrpu879d
iPsIoEvQjDBsv3I3C9OPvtKbsoj4XIDPM+yOqhXVA0HeBCWeqRUSC7JWkRPvmvQd
/FUd6Q01RjF7Vc1OTRsH2R2UjZzmo3UA3yrouh+j94+ce8/DOZHydo3bMAYz0EP5
ROdoQtH1Eoy+WGQNh9OzrQpZDHnKD4xbknEj0aDRN7PwQa9U7s+1aBhd0fOGPqxH
5sioUikJt0QinTNU0+1EaPmG/kGhHoJrKiaZQFhOSZOhy/ZMAO/UAyXiqacxKm59
QFUzct3EqshxWOojCnKpWtWwxa08KDG7U5Ehh8mUuYql+FqU9i/mtx0VJ4Ncg1Eu
QFqb5r+QDlxr5begRgtchIDVB+MV0oKTfsxKQw3XFRumpBz271KnxWpU9p8wedyC
MnvkFVuz5pPnJIJtaJdyOFQmctgYLexuM8CcKWGLGBg81J5oKBJD4RtoFTIiU5Vd
Hbh7n5HNCI1AxY1S5GZxjqDtsb5TainlJ1OV6PjJBrMrEwcLtpG3XIqu18QmYFAw
FbHzHIPu1I4Dm7luMm+GRBsevf03scQt/5dS8I6P8hcBnbEyCL4z+Eja1QuBec7H
Sjg5iQ3mdl9e6GfIEQ1ccaxea8YGsgsWo/vILlfLUG4C2uxp0eg31s8vJH6uYI0y
War3qf0bS07VjbyRk/Mmm+fnv33pNoRnrHu+0aHtLKSq5rJIJn9ZQNiFgaN5AeL4
VhZhWI6QEGB98b5behISUk6wDXdZuRyLi2dByaEBJkR4N3yMkFa1LjcPYXt/20rb
ykTvobaxgh16gsRIz0BFMfQhethOb3hudKTEqemdEW8xz79UI9MtLMFlgctf3iJE
BwFtzArl+jxOW4ZZxnFqld9dYbzAkodJEt+pEmb4Uqect/Ya4qCkKN3LbhfN4bsV
4J6I+u0eMQWKSAv6tEadvkkl63jowYWQ90iTvYVjy1CQVbdD92iLsv1PgxW7oj2l
7bhP8JjSGUjwmNLvvf1Tk2TxqOqHvaKESrPUNvHIvhQlItgqR2004ChK2KvNdIbl
ZbVIOo+kMTP0vt2adOoY/jJ3AKt2XAsLAnxiMqVIptjfYz4o9D29eAfeKxQgiWc2
nHJACmU0dJ1U4OgJ3MDZPob+TIuK2ZqIRER3gnz2M5E0n4aDZiJ17LhP6wuz5jlx
OC8nfjApLg2OupTH+Hk1i1GI0cd7Q6yOLeh1Vgchnc5AR2i9vB11zospuVTHLc93
sU/3gMgCVumTzLnEtDSg3pW30r8lWkUu7XEVb5FpCwnN2p0J9xoe3iDy17YPJRLx
0ilbIUCobiKkgdDHg0wN03Gu1lJwovjDpu8Q8qNFIJg9SeiP/qSGfCo6PN/miUA5
qyk8QuC8sf0rbMtpq5xhjOjPCvZZPVaxal1JZ0ty5B3VscWbOgRjYN8IEbQEwmMQ
Ww+L1kymooivrMEN4uA4XokzAV9972obvZmK6kS2dDrRJqdlqfBANMio59jeDYkn
qkIQ7cqwZHY4G04GkoxPbfNqqkHYN/wQm8ay0cQuJrEV0vSxh+4urCXjjorAPGcy
upLbRTi+62BwGLfOmt+uEe4kx6VsmxCvQfvjvac9wsYdqA0Z3kJ+3PNPhtj0jSnt
SQp0IBto/corGHTpTEHx6ajG1jijSBIbQsFDXA5j+r0FBYylZJmFHuPIu8mqWLtC
Ht0ONgBaHM7tN+7BstquV/QWcORp+3TtuH0xnFWBK+UM5tnvo7vLYYANd2sjZj8E
kedtkIcBVYPqBD4t57Ojm6fbXOUS1F8Ssv2E5SE8YBfApisT2TaZXCh63MpI1srN
6wlqRy8KgT3eLBSk6RFBEA5mvwgEtVXujSLqaUzf6Flt3tB1DwOQ0UxNeDVJZlhM
YArUzwE8g3GX8JaABGVZp99ZWhucSG600QBbLmSVkU+3ThVvxCG5u1mM/XAAfiUg
0UooWzqv31cinJQBCPn0YPmZ87Qqkk4YucYjKE3PzP/ltG8rQHI09QRuYkyXprXp
0YrIiLeOdg4TBD5fdeDWwjHPU3B60AzNqW9nO88MebgWPyZLTX9LnNUnBcdXjSv9
6Zqzbf4V3T4CnokpxKkN6HVcynQRCakECRjCSxw43pxroslA/7kk/QtplalSRnjv
v1TnWO2+inALllwUVmzBeC2Rls9LRrZwt3WTSBJxMqszdWYw0g/SKxDf3GOw7vM8
e2EKW2Ie/Jl/kyxwmX4sm3FV8Gx4mlCZzgr0EpDjNmPgCgxYowqwt85pnwKAR4a9
2BLXbSPaxeS1AdpWwXveFCtdyO/oOSnUNnZaxjE1RXYO936u8+UhACRcAhcASZk1
iNTZEhpLl8FQrJ2jcV9KeqQvlQFIsAAt3RNLK1sX14MsbwEp9AyM1IE0KzJc+qfu
Ky7K1taHsVDvK6Rt7ZIMjtMtv6mjCwThjG/klnq4g14EYOWHn27eYf0BY9smCRW5
pVNFVKilBvsdX6Hp6PDiPMk7reH1bB06LMXXgXllXTQ4JIVJnEiVGaU7stnk08ET
Z3QT0vfuoSDjls2/RfQXlqCKdytmVnJkRlBDD5wnwPdK+9m1HgetP1BPpArjaMU6
rB3XIDC4am9L98v947FEDaPdrLySyZGplBSt1nkzvFX2ll1f04Oam567cj+MGtYe
ywMGJEXUy66F9wR1Hx/8TcbacmijhkVKpdLIxko3m+JLjmj1eESRkruJKXuv4SQv
HRWjnDlEerqdBCyc/J9hH85W6VL6ePFNhmXmoBz46jfk/R3h629PY73DxhSwXIzs
FUpXFAwP3wGVekbLoioOugmDjY3DVWMRscvV0pESPN0t6MFkyHu0FQB9PoQkQZdV
f0zNxnhRho2FCoQn8GdPc8HScHPZIkinaUDd/doAx8HKcZ8t4zOtHYDMif5B9Sby
3CZZ/mDn2Pehs+wlISDCxQPQsasuPAwO3RhFxyhJ2ZY7oosA5ZN2EwlivRvEAr+D
ksE3zwjULQiKbmCOCvFK62RoiD7ox7tNTase2QlIYHTB8Fkf1KVKp7Pz0AhNSC8a
ZDJCmZtkCoH8SldkRyoJAN3JYj0PQ0N3jE0QeeA8giBqE1WTqiHftG/t7dMC1kFp
vf7xjkqSP6/fxCY8wpNWf9PEaAkfhXFmuO3W776OpwfRTFJDrnxRyFIppTXIYl1R
0rvzbF7mTWr8JjEqbKi+SHRws7nT7hy8JCxbuKW6g9cb6xOocgKZ0wd7/zuvofUZ
dFanTUDSoYZcQv3Xn3Qbj2vev1vK/vZR+p8jTeRFk/ei0qkDIwjmGhyLxoCx2MZ8
uC1C2LJ4hZz4trMlyYUFFkISwgYm9XTEWg3okSc5lxPMF15yRMN7gxiKiJzQWzhp
4amFO8opME01FBb6kP6UGUBErVyXEdEIup/s/VEIjmE9KOVj1O5sbIMA/AEYhwzE
hx3Sp6kDDWvkE0veSaNT83mwi6exA4H5tOlST/1a6v9z8h1QYrKkZUQpf2SK5fLr
gfmiuWJBoeB4ktBAS2QByHdidwbFH8IKxy6I6OCy3s9GzNAcDOfC0+F0kzh5RUlK
HLAguCe/WtKmXuv3OfX7utH8WXMH4EQParbb2SRWXU+qH3I8lVlj2CYtxTquy4IX
kbCcZl6HRd2yJtiouqaG9NE38OQ4YqkiXG6B4LUF1leAi+uOQmKbV4aT3ncFCuYy
4DQg33lMqrj54/UXofynCu8k2NO4sfmUj7SD3Ly8gs+7c6AyGny/IbxsIk82LjIh
le9CaacFpyU7MQ9JUcnrpEgMJ8hLb5ucYUuCGQOcLdfbdSnUfE4aUHtx/HG+H19T
IoYgvMtsUfMc/JKRkwDH0XGohTjteH8PhjWJBYoIyfLDgZPY7chDe8DFSFXcasNJ
dUsRfycU8N7bT4Y+mOcLsTN06amGNP3mhOvWZD1TlRb0/xK31fTTLvOV+543KI+4
SMtV09IDgzDjeUmoBz+7Ombsk7Lxri261Z45pA2TphavEfHmWpOD8UAFBADD5IFu
xHTi3XxPcPsfUjwaPaOI47V5azyeKtLsOkeEi1+TqYstjCNmlfQat2CUTmtsCYS4
66BqDt6r0cBKVlklGPJIU5ktX44ls5JQYa9HgnmxpXhcjmV8b4Y2QSH5kGao+Mea
m6WMm29/zGZ/JaEZtfbAcAxwQMtwMBzou3xgdHTxFvC1kMBUhebUKYw55uuGDuUH
lrJUjYsqldrCDkVPWY7UO6oLb/P3LUlmqSuS2TV6hCL0Iy+79+UMcNAh2pHNHzEK
0/55dS14SBt7vIw0LbrND/tfeVZSsYssdfjTLt+0GwNRyMq2NIp7vTtPOnv/rimh
s6a+tXl4kHnYINeIDSExRv4HvG+re2IqAI4hTzgjIGgpvqf+EdZIJw/0avjC9J9/
2C+m5MofxZdCBVYXxpW9C4ErRCT9YLylaaBRhRNpO8iWlDETJd86AoBzuyVkU+3C
nXnuNiodAdXPEdG1H2LneO0KJxuBinn2+KGo2GuPwb6Vd3tfkDKXg+qfrUx/dCKE
FPf1JRfiNGUeP2bCGSAr+nTNCDSZcXuznPQjYW+LIeU/mdastD/jr9y1yjiqZnXR
zZPP8GbCVhrkSEkT3ttorIpzDUekwUTchMDBWbITvB6xzXDhdUr2fRMbPM6EjfB5
sZ1nUAr2Qdroo9WUxZZuBjXgZqKU/+AZQBZmbOpgjZ2JAeNCIB4E5hEOwle7e8WD
XMKUuwmVIYV8UcaSGa6Dd5nPCjryzVxGcXCmljHpnxFaILnnV7zJ8pwBPMDLk2Rj
4cA9GK2t/ByrPZuq/fdZDUIymf1tHBchYD24Ntuzvi6kz7+J/HIIQ5ym4eiCYIq3
skExXWOYZpNlCGNP0yicCh7k2mrax2aLbc07krsW0G0fVpj42iRSlQ6l42C+tWsu
j+oakkjQKpQcvDS/d7CWFPcdjyg9BSv4NC43qcvZKFdzXSE18Zu1+DIYBVuEUHNf
ngm1rHArgpvW4EJ2/5/ywKMHg/pFocPvwDZIm496zAJpVFruc3/fNjSPvbjJ5NNF
LicDApvXhnHwa4oy7dfB+Rq2+M2WZrzF09hhIfWKHUhRwZRGRHgqd3ZgAVq0VGLc
FvR1hjBcNH2Hk7raiHIYbSATVcNESBSn5ma7j1rkhGEzRpi81Mw4GgyjI6+wLmJP
Jhu/RZAfuK6fqGk2NJqMkZB2M0bro4aBgjw/bv5/sqH4vdB9SQTAcLgqwZnybAJe
03a+8bXdtlaOHxIZmvTYYbS+I62Nllz3fqJdXRImMpBKAUmkDd2aB4FCoq39sjTK
nLsW1y3AyYPqs3GmGjqC6xg95WJ6ZgDLhq6t1PapLKWkzhl2DKHQGS/IBZoRHgWS
ZvwWxK9hlUg1+C2E7XzrUc8mq61L/IZS3f9MuAcZjfx2RCVq4JcW9dIWWAXDfAp8
f5ZsT9yPBMip1q/Dv7yQAuPjcGwlfLGevq0+gItzhrfOPGG+f4MEdyZq1J2mCEut
gJgywHIqy/fY2FgixHbOsiYNyPuDJq6tdHcx8Q4r6Bd9RW7UakBPq7NVyqUvU8nT
qz+cORW/xqIKCU8EmmazAQgaxjrWFhdKak8YvKNptQeKjT4pZbtW7BFmFo4FYQ2s
77b0gcD7q80b78KzWo0ictfs7+ShL0m5m+285uc+eAsjq+xdeYWBi5ghchePWyZ1
OLFjc/QUVAcNdfCJF0lQgyh9x1vNeTvzMI37eR6cbWbHqS1UrXDJhv7JhNVwamM+
vBCwJ8/Kbc5azWfq1glEU7B+lPjUje1GzpoP3uIr8arHVxqN2hnVPm/W1OsTXqTQ
ELHT2gPADuB/FzjbMoIwZSZTD0SW8ADxoXfRDKNDpC1EmnWXSaeQdUwP3YEDvGhs
ZPaOzBE0hTNfGVUB4uGVSWnnh/mJDIWPikagv0XncYkqlV22B4Hd/gu0xp34eoQz
QbRHWlAKVVjAI9IiHUhJPtcFkT23ILvSc8Jt26/3obMnKpMuCBisU6amTMbEARLG
0PBwwRZzpPgSZw80lpZSQSicCn3d84ppzlcOzFbbwDcK//6h2H5rk4Ao45LtUxZ9
+8uqNmwwEw4ZcsgS+Kfwkdp8zk2e4xmY+YDF/pJHfgxjLmwzR/LeejYj7hXAFPEQ
qIVjrv+qAAL3Rf+IApoeWDweZCWVdnBXgHkM6OpqgN6m2ilxHiO9yA7XWjHdeQOY
xrvfcqk1yqTTCBJ5OD076JFmvhxVe330axRchSo7NNbWg2V2y03TK76/hBmHII7j
jJUKWSNO92hGxsjDgYg0ntBe08YpQmj0oG77TQcHym7UWZixaaIN545bc0UEp73V
TP0NB/eAyeGN+ZOOqOlg+ucEA65pz3Zci6cUL/nnj4K15zruHGVLSSff6kcnCMU3
6n6ZfC7Q/EnZobDSIznlJOxsK4v3IeCP9gtKoo0bhfWsowRpirxHh6/oD1Uj+OSp
j04Suglc4fMsJY0AnHuj5fElPYefyVLE8mEhv184YesSDlfZS5OWbysEZq6+FjOJ
rnX4/nlxJaefJtcBgFsMEbSDEtp0b9aIlFdEnLo3UL6JKE85r8NxBO0SWwX/Nhwf
B8X9PJ1Dm/HWwOG+iPIEZCPlOGJOiktLcYDiiHZZFSZPLvuaLCK9W2vCMqDP19ko
aR3kEahtQEHS8Oa9xFWBJ7b5ilK7dPTeO+qwnjMz5nIx7skkdqfBaI97IVfmlsl5
Gp0H0CqxEBR9kyWOLHpevH3A/4Z10WWx+jvZX9yli+bCYNnys7uhrGITf942f1nQ
8xfO1eKfMFN4Z1VuBj9ji5FNDuu+Ed7Fl/fKcKEQE7QU7/JuvV1fqibLIH7cpKmJ
pi7vZVELl4BYNvIY+92N47vteFJbQtCAtr+SCxOB7k8oqPMPugy9El6m0qEkBrcl
qTbcSFCpwC1nf42PasyWUQxkTzuWpX9zm/P1m/wJZbQBLCroofDNje2CgkNCUVGy
mqwTd4RIO4cLDYZo/lndkAKn7YeLaQTSXR5DjEvYL9mecDnBE92mMKG69jGrDG1/
RTSyFMs/hNyn7KSEk1AF3qOfcWOQMv/QMTc5jKMm9gE2+VQvmUf56YbbqlR/O2K7
dLVaxkDLNgnPobv76b570MPLZrRgvfXQmB4ZV1md6D+vc8V1Wap2z1bJ9Unw8aJP
f5YC8MO176hrGnwP91hFl1tf98j9fLSMXlgCTWhWIIxl5Y/yngXXPG/GwyubOl7Y
8255+PvFxHNVARQwgQwFCLN8L03KL6yMFMCC4ZN5oq2zgEYDbYoKbdWQEuLFN6yU
tcVbAOtVcSKAyc5WPtuGpGRgr8nizw0JoDF149ZTEiUxQtXB3mdtNxz4VDMDzOH3
cRSH7603Adz8JndT5AuY1du9aX3B8f/Tja1Qcu61qyKn4v02rwCRkTh87z4EdBI0
8+yKPHVxJ1MA3TpieRd+C788UqJvsQt1TEo1qlFKDXrw5Wzcrz+YPlDlspEMxgQr
dQEtKfwrU0G5+SDsoHTKvlb8RBUZnkkY3llI5+fSQdTOcqEGCRb4wjQFDjVXsj+E
LF/lg8LqW5OPDpM9Lb3cCHov0DhMrwBAJDnu0ffHgYEjI7h0VqNT3uQvqRO3YOiO
Hd9Bj50Xt8jPzB59PSvvRzANg40SqkqanS5opEKjQ/dtWdNMjW7cMW2KqsW0HDrS
t65m4bu1GgpXVEcOYFzFF7QxO+KaPAe0jctAKYtH1fw8VRpEXavGlF2JuYvw2NHH
N5A+Qu2QcWdlzVJlFsShN19E1NrFQhE9HLAczGIdULV8Wgc80Zzf8o4hMfl/3kMq
jFwEZpA0AWtHTjcM1cBwOO3NomnQSC0HAh2HWhfM6312rBJV+ARS60WnWoC3DT0h
jK3ZzzJkl1dLiBemB21l6u/GisYpnlqtxnqDXEwTI0jQqoE7yo7IAnOhQwgPJLZW
X+2VSnfyjHUXno2Hzl5MELrgzWjc8t+EXc4V67yhqjLqAQpdhH/YBzHfuKSZDdBL
hUz5aYZez5qcR+aTIfttWNsOl4HeIq4euNPa7q662uof6a+nTVwp/uPtrb1/8ifS
QE3OOFmdWBcqO9hV6JQ/L+yTqPCxv0o9e/8mCb6boIpdZKTYW7pwzKBIzr1v8EI+
MGWMmFo2Mqi6jpjBtaj26ohxn3jq/U6pACvVH26ny87FJc92gpyTDEN3N7KgeCgS
JTrEZUIoDNIYHKkr09HhqX+qyQx97+AaOkNK7fKdqEubdSzWD5b+hWkovuWzL109
DnhUYcUeW4B0En2HfURSwteQrwYBQg/RuxcOHEXRupjuGMqn1S33jhBYJe1LcGga
E9kLJAOEqznSyl58ILk0xsubJWWIAHEq+M1fqN8VxzErb6pwXCA3ItYL8QtQQa6b
h1LHQeII+2P3D81+aYxSbShwHc+vaShho2LfuPGsknAgiazfot3LlnMZyZDhf70b
3w16wKUeuIheXg1SQ5FL8MeC5Q800oExMWmHTTKn+fQCcY4ZOI2R8unDRv5/0+zi
jiN0+N9P04bXiNquS3LLbTk1rauEbczCKk+2481VISwPDbRIaYbjtxck62pES+ry
GeZd1+aHzAxXCz/ZHofmmB5D0RJFj2CYDLldDkSHhkGOl8rRz1S9ZJIx8a7jgLQ1
X7/Lvb8vT/XzU5I4mw6IAS84f/JbroEbTE28IflOKb4oxcY7N8pnd0L9FGWvZq57
Tm6NGrsRnd7z2qgtykAp+wJ2m7XBfoBBeqarxQ4tQJ9lKs5Q82k83hFJNkBq154K
UKsNN0u/+kSaDe1cHrn6/F4y2dmy3syLhARlLSa7XCSPrrnk6ENqGy0ttsyb0hyG
mo0ENuVM4j6Cbb4mBNPCXjVwkE8Hb8ycYUG3E+DvkZKgQ2igB+betK87qfhjwqbI
U2WpwPUnvWBVMNh1on+Jh2G0gsFnOxguXtzTT+reyjUkLBbfKHmJVlS2q3L8wVdj
U5j6qJ14P9urn9Hn3+F0dR3e4chvKd/FXzD6aN6dWRFVvf4TM+VZcIy2oHZ+8TlY
p/IFsiDbhc3bYcK+RZgBcAsY41JoN+dvKk/EnRM+qbSvufqPpwh9hvfd0AfYXMKm
81cPXjNBR90ixMxZpTvlwyBzGFoUY9+SSeCS2kMax/N/zckYB2z7nxbRZuqHGlQ2
Ae8f7fxPWoP5GQTz81ZEIxYkreKevREKE+QrKorBuLxqpnQsE7CNN6pcSKCuzaEF
eNBPI5Bsysb83FUyrMfKDFj0ub+yyT7JFkfrKHnnmwQI1iMmdck9zTkWQwm8wPzx
RsJz0bbG2gTY0Dypg/NdyDqKFFZKUowCqzXEGSZQ9yFQZL4TMBF6vYNems32aoBN
FT3KDvKDuuoWVcA6Q4WMwUsIJPk2XLzdsAUlc+G5T6A0qPzEFOt839RtgCHngMdT
5NmKlPgY0evtTskqT03+vTLY9cOuo7hikMcSBVvlUSN4S0PtXNZZahkfkQeBB7BG
9J0Bee1nQ9lwFMVOdydNYQV4VqPiLzBMDQ1qcORuORBcF0hf5VDW/730NlUF+Yhe
N3J/ZDykkgvE1gih/9GL5twFWbAHrZ3lBkLiRfqx3i19odCdtAKyRFV8LAMFr3xO
9WKF6q2t0uLQcPIOVst4xx1lddTL5nJ7NpnKGjmN9Gqd8hAGRrK0m212/lYZaU9t
ShvG/uXnq7KAhC+pJO6MD1EsGloFb6OdEqM3jVW4O4vziJQdPBBvMNmcJ/V4Z1GF
jALCbcbfI4mB8IQCYfafTDeiICh1HbzFzvVjC+sOyERfNOd/iNY/FRQ220AILuYY
sqYjHGiYk7pyMa7G7UmWrfVUmW6vbMZBBsie6pumzm0FbwJdaNHBKIrIgb0aKkrW
fKEVk1Ge+h+wxpbeCm+jhZRMmtGBWEcpJuiUGXFznCmsmR/g4G8qx+rbKB6aKE1v
KaRTLKxeXo9DRlILEPGRhQxLaJRqjMVT050lK5Jo54uXXfxcg9oH7UU5Www5JqPg
hTIOlubAsk2cwS/pej8R2+s2Hw2K4xQgYCRAFDoME0TaQzcG1ZtcxkzSTvTQVKP1
hDDpw0Fm8CsqUO7aYaRVkykc59PMt9OBkXedPh17RveQVbKe2qN0GLmnpboQ/VZR
PcPgUWUXYS2UIRLALClZ+zss6UmiMXRnAmAdEIqonacMBW9Nlzc4NWNmJ0mMwHy8
rIJHT1zTAAKusIYuZk2SqpH78aaaMpqrARvyFs3aDC2Cq50CIxM3wfeLNTG8u5lv
F0BQlTnrBp2KhZBYhVhUA0RckpPy1K2TXGcNkFsO82kZ6ElJU/iJWuATrL1CCNW6
SNM0oenbNEsqv8k1Yut6VMKbpZIF5+7F9wB36zIgmDiIIU2gUeOQ9XLxPAy+85k1
NpIBjEKj73n+PSr6bM/7RJGocH1HrZteUjpkrOf//qP9IETy6yExg4I19HvpHyzI
guwoS5EobIGeFQPzcI2MJsmyja9zSAspx8C8ar+XmHku2G/W0VP6os4COpmGaVfH
4R9DDuDDJQQzaanixncS2eNjJFgz+UNm4XNQhkUppn85kXMwVbqXdRY6b8cujJlE
I0Fcy6SAubsIA8G794dwCxZJeauDi7f6zxR23B3U6L/aaldpGfTukd60kJMOriJp
fhRtpiFOFh44yZ+16xQF9wUFCxMiE8z55tGp5MvP6xfBbEG4oAgNTnX5K8HYMxTD
F3ZejBO3sC6NR0QW3qQNa+I3XUxq121ZJDn3G6T/hr72YoBLA1HegAETJHvbj4hx
zw9P3BJSsgljQkuhpNlg5GuojZEgBIBGfFp88a77a2W3VrgwQR25qHiJvt3y0GlJ
kEj/2b+hW+1I+1kcqo9Z9MpcOfD4okZ2FJOiqYangVCzlFLiYSfpbfuuJ3Cjtq66
XQJ3GYWz17DNH17SLtw9tnsvo1JAEoSUnR86Z7Fc7RLqnzDQM5NCVXsigUGWX8Qc
n1aMdmulV+ZEsuHUZEJEBTSAQUi19sXVIKlfCVxh6tIjxw/s6C5hidku58D942Iw
dQT22hhozogCAgdFezCZZQu++8M4GQN39Bz/gKdGaDcfWNtwijPIaNUV85vHGPIM
6xMxIe5WB5cuC8mbSzdpFMz8VcAbY4uSnZejfeNdbfCKn+hNwW/+8VVguShH90In
Af7TAaJKOC76NcbQmBLBxsRE7cITHBfqyHD6f25hiiWC9HgIcL97icv9lH6CRXSg
DirGZyYoMTyq+79J1OHfqoo2J00an/9N4RP+NElBENZOzxoxtpLvikDG/cd3Ye8i
rDWVxDmUqPWkD+/FuYaBXgHt33ZXZYieV6M2fBdk56AOFcaf7da6fQEUnwmCD3I4
OpTYcEZX1SssvtXsAjfmddD0XBknwgtiLhS+xZUDwvO5NpbQD07JNyaicMbGrtb4
XPueCzND61bzlLmsmYUh1Lib5SKb8kPs3BwpLwzA266vnxPuxIypQacoVb92lT9l
U0jEInmV4B2Azhra2rngGo3wz+Ov3xavImxIFcWwJsde6ZtRi7SE9i2ILMOX1dYk
/y3FynxcO7vEZQrqmCn6RkoEdU/qr4kbR6OkLpPPM5Cf5XP8Z/uzWqM73oqHv+bQ
z3ebAMHa445EIN169yd4CtHqeXK4WvEGVH3tDrzUascnPgf1TGz7Ezn9vBqBBu1G
SZqJ9i00Fb17RV9PeH0veWe5DkwjTIS557/NoeOROdPL3tUy0T1aRQYpY/Ae0jLt
rTVH+OIxTJrGV7/r+qTw0tCwnPPk+wTPNZ1qHZJB45Np/FwgqpBfkqoUQxDV4TbO
2GA7P6HUPtdIx7g+dfPFS5qCqbsmgjarnPgzmGYsnrU8Ka7YaHB72KuapN53R4oL
77BYz3rmUYW45FLW27bRTZamAQLKwoyXdUDnxDRwHA00IYaxp7Jfhs9zMj7hQw1a
Sp8rmItTykiELnklulx4OqlvZpo10Awu19AXcRs4MbGH26/wJKiulKKiAg3OCpk1
93icS4RothlsFQExhDwI0da7XDWQL5hjUFSrrWl3aw0GHUgLO1FTCEauyKbJXInL
QZ3Wheo0jS3SjqE6Th2v5i3gWT5jaO8FBH7nRyC14BthuK12/CLDKIRMR6xaVlgN
RYmPmtHLjPU7Qvi2x1dQ9M5OIZreNQzRjEfBa6/rnBnNGLfCLppuU6JHUe7f6y80
y9wQ2v2IsFB0sHu1kl/Q/Yv3ZV+6co3NkB69ZPGXTX/4188F14A1MZa/JaY3rli8
ZDtDRt7tJLRtJqUIAyNxd9t7b/JxfjgtP+bEyapRbVAWEPWJK+9x0IzDyaNR5J4o
abnybwc8iUtWlZoao/Upkzehr8/wCaWWLK9qLPNjEdzJfQidLw3VrEd8xAQjIobc
JrviDZbr7nrQU51B0VnZPqJesrE8vP8i4B7+k9ay6RYLl+ifdSLf42+z2DjCKjO/
jVLnaY3kKXtsXQrVcipLT9/raZW9a9xyZdokGEIyTOi+LYwZArAqepHY5QIXZw7V
tfZVsamta/aT1+d+qdmEgft4d6bS4Vy06AkkNJTivLVDQIUAgddfeG8sfvbaY8Vu
NmI+dy7tErjAEX3zON7w+rghBdUkHq5kLDI6zDNzcGs1w5EiXAfu56kZGMo2FC6Z
Af58on21n0QBiIvfd96MMZxculcvQ33HObqVV7f3+CK2XjzdNQ2m6ooJebHsbgLi
ctbTw09zOHXOsyugw5/0aRGLILGoZp9q6BU4l66z38735pQFtGBX/nshKXPVi1iQ
g/ZqarG68U6VLEE0lUoemx+chgjfRqvbDR206rSHTiZl8jZHg0fL9wo11bkwhcAq
iKcc2ctqv9/hQU/TeuyAtzdylF/6gQTSRe8I4bCWPYNt4Xf9phwHK5h346jc+f9D
1nU23082HbjTHqDpC3MO76eQTejoBeo5S92rB/JS3VPdFzzEYEJeyr0fHqJe9/La
iI1QnrbjF7sGrE8IxVj02bxYnVjzagMDBvY+B1BPvMxuLBLMfrBMvRnGY2n37XCu
awXEOyGlevnlj9965yxg5j2iE08tBQyOpbeJvumTM5FS0LOrzPtqW5U8Hg3eezEA
nU0h5maV1pmBcgqWg8uoagOlO7i/2On2T2NrfOC23wUXWlYarBUSM0gLnwqpy7nl
JwgOWZLu3gMYTNL4vDtKyk01bzCqK+9Sgw/nLNS18B7NmA2XhPc5nOvS/HjBKyCm
IbG9m4uq4/irGAxjwlRiASBeansxoEl3DILycjAAtPIW9ACM+jbLxOJ7HfpdY1T8
JPSlCPYgJ/zRCPRqtmGQQVo6VOmUxTkKuUAGy/UK64o=
`pragma protect end_protected
