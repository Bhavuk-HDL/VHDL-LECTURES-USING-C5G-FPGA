// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
veHvtIIhVb9Fr0FZRom+kYMd8ZbvnIzsutPwnjcU9bJiFm/BBOY3IssfxCGxDvFXPvoF7D0S+dz3
ZPp77ydHes6JG+YlYxmZsDHN+IFuBIqz9pi/5cj7xErm59NwL+1XyA2RBNK5dBAfLPj02FOsps+w
HIuP49SexzdhH53MPBfrjJ4oHLUvZlWA5l5k+HV5MkPCuZ8zP8HVLxpW8fZ8zEfk0u3AF/nzpCLy
3M8zHGJuBe94rs4fzmJqkt1DL7j8kI7Ujt83YX9/FTHgwD0R+swRnzMRwobVjwkF2ul9JOgt5fhL
iXbGMSBlG7wPo9lgADEgr4GKInOVdMmtffkt5A==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13744)
onBMyictiubdFkWW1b94+BpIzDhrBBPDWOy1AluwLMmprZ1x8Vo0txyEeitmZbdCE2+IOdNiwW5f
9Q/xt9tNqSleF+4DbRCDPEl+yMJnSakdtVazLQfWsRSjHf+CYKHtl1gfrEkeVOiaOGGy8vUKoshK
9RMZv6bvrcHTHaJjLKDp2sh6+wRBi+GBAVdBKG4pVyYxKa1CpjzfQtkrVWtIdkIyFqzcw5td7cgk
QY2G/Pcdq6uMM1EF80apo2CCWxOcm70XYTpIMO0eqTSAkBx2tgcI2Ju2TWUvTtX8CtaGz55EuVd+
J5Xw+bXugqZ3E00G3GsUvaX2+n26OrypfLGb6AIndbZMxd84Yh2btGaqim8XkkLmqIXBZLsIDHFd
iNtYRaFy5hrXVGueW+Kz2KExVTqTHcQ6/tcOV4NPBl4Ek8uoBOKOqv11GzJ6pRKMzeUxYgZ0o6d2
/NPFvq4onJnfSvjJcYsBAGOzo4zd3TQeRKMH7sEkcOdUeo7jNv65mwSHo4D27+sXuTMwboQee7sG
Am8ewIb0cse9S0pQ0R/sFl1UPF/TM4OXRBVs24mJxR6tu8jyOy6pTOIhdW8pPtzIMWRJkSGBbvnL
IhaccFc/yTQi0TYhWmFqeczBICHNo7NIZmjcjZyG9JgLBru9oCu595fVBeOsa9ShxIQZsZNPIAma
Smr9A67E4IuS/7lx7dPULMT5LRnwjRDBCntHIGq/DOlmdQjw6uuzQY2EyS12Rt6xf/wrPwYHUd5m
aAHsKE7zcM5NYharKr0bXEoe9Vzw+zM/XgA63Vrq4bJi+XDvN6D//4N2qguVDXiGkUFbhS4FSuzh
btjPXf3HEXRCP35QU2S3fwIbjHCMrwZdxL+ERRV5qe8G645ph/ft6TEfGVokTbwRHoshwPvk9y1f
QrPf3peFPSXE6YiV0s7a2HAjFEfGWvzWK1kbeFHNyLhSytavwkx8pNZ/4PDf3IR3IhMxeaWguCAk
uy5V/k/vw3bI14cd8lXpSZ4br3gqpDb3uW+PJ84txWX5d4n9+7oVwhC1k9Ofm+0isiO3bwL10zRJ
U4SRy1W4WlTqH/zAgnJLWzBuUo7yXEqeB3Qppshk5ckkf1WTN7QEGKdIF5D4A7I7vSAQovazI1oU
7nwtntYiwQA0e3l6WdYyqD5u/C3bKYlDFnYWu1Lxk4ORbh8RAA0rXzhESFqWiHfPauk/m5SxPs5w
KRl/HOYr2NtinKfyivhKCl3PVo+26zW2LMdjVN4qU10d1CzcM8Ia5bPrQdTdwGoWkD01bkxqla2W
Geg3RdYzS4RB0RpjZIVGqM04CyUImfs0SQrftBbigXLvoHSrNuXDX/Zb89NaWary0TPUly00Y/Va
ecpbrRyCof9dyLJarTNzw9zzcB7s8mAXjYI96LG+OeA7kjFKDTKgoZj1VOg0B2+zAqxVDscrcr4Z
cG3Om/sYcCJF3LgngzCQSvQ3taa1ElXh1cuiZVQbgCuskok5EHQBbQVZadzyyemGCbDby2KTX9AY
NvYDSbe0dVyqdYbXt/IXYPRymFS1E0zHV2uWOpKKdVCmQY+G3z4cypzX2B0qTD4pGK+vQ7slzCyA
Ahg4c41/s7p45qG50VJVCunOOzEWuTRTPn1VwE96ARKztjfux3BXdj086CgCmxsEQgnwB9P8yV9V
NpzBrTa+BXWisdaH7Lem6Dzzm1PGEcgyDplc1XCQgq4UwSyHpxfKrxsi9O+4FZY0DS2LN4nWzep1
6CaJS1COtL6wN6ORMqDEGeivgTYcWATI3ujlA8q0SWFTcGsg9X3JeJdfxHnqgwJQbebghZI8P7xq
nIRSmLmE1RUyyVqEQukFTuoK6Z8/3paUkkhWM71+tc6zXIbtWxrb/smaVWid9XhFkMRyrxmKB6pN
JqiF4+q/NnqwnnJLx1ok4ypUeJIhwTlEW1ElDgQqVGmlNlx2dikphHNd2/tnPKPeHYXyNQdB9eps
CNP4fsQvERS3NOeXfTUtPHycA0Jr9AK0z8Y2aOnxOcIJWoLyf0qF5vbSKZRt0Y/pOnRYuQnZUbKD
ChJ/XIaRLXPrKDWt87rQ7VrNyaHbtlG5YZSxl8kE5TQ19YpGnDaP7M0RAHFVicxjQUBhKKkk3B0b
YA3FGPV6J61Rund63oaPh71XgRbFpMLvzQ/16Hn+7VMpp5cHKcipltDaBYY8NH1wy49behipNJ3Y
WeuKUrM6sJHu1lgSfrg/ax8//ldzOg5gdhtvZvHaX1KSRqoBKoUcmiKt54pZ8THbQ3EOeCsuyTsu
dk51WIkXDEgYfrxKr1EkgXo9Nidjs0NtFW5BCCuj8n4z39J2iPLeojZ8Tl9+YpfwC4959EXFN7cd
ObnUMvy93bjFsbJbdxU9d/sUnmH3tOn337joOqdKXn1I40oxdk/S3GhkNvyVMpkwNtLK7cmF3jJ9
dA4kkSHj6nNphlZ3YNPJecFLpPX7qgQpszteAnIOBFv7NttGlCxBY3WeO7MZWoJV1g3Rc/xBox+B
/uPjlfFil5E07d/kYnEs0sZsFrARAvA/wgL/d11u00N4cHKcr8Ip7oSRAiFOCpxUVCfqVcaE0Gey
hQG478AyutfMZgcgsQaJJ6T1xcQCsgyEluYGlk9w/vws0M/Z+TVmKtXFc8kM/VaaS6BUv1rbUIMH
M52ViCKp9ypHyjMVCbuWHwoz/9fctsn86IcdNznICNV8o7Sq3PzBspB0lWxYjwqW7V6F2n/l+Tp9
WsPz3nUANOb+qF0kfNHf8DRYItoFH9GDO05JrCi9nQ7kFprp8khlaQypMGCoHksv+CVoQSYztijP
TjaNs/R27jjCHvjz+xNMpQ6ieY5NSOKbqf6WgkxDUO5ywp8Myll6aKMQQNra2fXr/XSpUsJFO4jB
/5q6RZw1eNRVjOSfO/u6v2qnzlxiM0EMPUSlzl89IRt7ZkR1lpgxm0w02aLFPaMQNXwNks7TrVbA
2ujy+x0nYBnJbL2WUCV7umsg2aNwGnNB1t0Ie4kbWgsZP+xtFcpZmMbH9lz6pMM7NK4yMpFIKV6+
MriBCR9iQFr1EPvbb2jD5rZxpcA4XwnLzOnNqAVDj/TWOzDCC1OBLJDvFhcS3Fd3miK936XD6hKt
Njvs+s5JxHPf4YlvKM28kOV6EkPHA7AiS7tvnVnRZUgl9c2vTQ9GRsT41P+ruCOn5pEU682IR0gP
fb8wycNDI5PFGIB1dfndtKjrI9TV7qWnQ0Y8hetKWAdtc7dwEqu2z6+vnRdNOCqQEn7K8jhnqgNq
YdMPSR4bojU7N8d9xBvq+QEw34rJm0/DOnDe2IqPZnzuaRDuLuMjUIelmWqzkFKKy//UPT9wMIrm
6iHtUkfMjXIOnRVGO11mdRl2St52Bh8/6apLR84WKPw15LnfcLeHjs6wuZeSJqnMx/hM0ZsKN2vK
1fmU0rFcqe9n5e9MdruJMRpZqohwaXvP+0QBW8Y9seuYDospHbOFBhrPxJpXk/ZaK2heiODvO+ix
czl4r7dg4OWFXSsZN1mxixyJQcZjZUmGzZm+mxPRieut3FiBNGOmVIrhLkbxMGJOa0t18LWVH21S
vr03Gk9YsLOZk4iL58t2K6LXGk/cdoFJB1Y1PlRsdkNOXPPITCplDJVpn71oX416CXsQtfFYDVTB
DFfqGnrO+abfwXk+V0nyrEd5S5fDGaU01uYVoec1S1a76w7OcIJ+8+03IGrSfnXa8TlRC/ual7x7
JW9+BWTXqYsD39u5+hXqDa9rhukSsZ946j1eCK+w18hGW/u8UBgneoLsvbZQekTROImQbPeLVVKU
6qCPM+zoZWHs7cPznY55IacnpJ6Udy5/imz7Rk682n3YYUdDR7H16tfj7ajbZiyuWIKZVXJqgoUA
c9lhW1JK3J2MpOI5TTakT2GD0fjJ93rBYlIIqccoqGDHtaD0zl31wz2ldBfrz2GTkG6wwAigfMra
WcEM0s6r4V7BLVCURx71fCn/sQwSPxMddUD8gkM5dzaK0wIEx7I8d5vTXfrZBHmto3gTpqUzXGuq
D/9xlRuQzr26naUBB7RavvHQTKaxkthI4emPqQtyXWRTZfH9pJTu2zT+ue69gdZLLk2nqfAgCv4g
WSxbTpB7Hoa9TdDZCaf5wCtaY7Mw7oW50I+ugCCBbm1KVpf3iVQXbLX9vEKlGfnfVqLoEFgVXYEc
1wFwOEgfcnQWTyt2wKcAGdEjSj9mBV0btKesBRK/ltbx6YGdyR55X1GzTXxAgVmhA/DPOXFMsOvh
0eTbj9E47B+T79T6Mnzj/1w6Tiwby1c7KAq6NXBYnV7s1fuR4cvNMfQHJcEiMyHerXr4bFNwbiha
VFl+aaqWhH87utNkCYCVndv/WIgqu2b2Bx900pW0RP+Lnn1vqaEHs7vKQ2iIeuraTmZGe6jMsQ8m
CdAyTEw9E5jRSKOpzCFaIvxNpGAvhJ0PM3ZJdmBNTARZD08HE9O+dLeCFOzEpne+bI6pGB65p+nV
J/QlE4h8z2FgaVkXjq2ZHgsEpFz1Z4Qib3iM+nl1oHUA81+cvP2do/aP1FhBKpCcImqDg4nR3bda
CG2p68wIxAk+gLknq1wuonc57fnlepy7EggbwKMfxwMeMZa1UEetOwYcwdFqiQL7GdQMeszlHDtM
nC3uxjaXO+gmC7rKs0JDP7k3Ihr8NQC41OwwL6m82V/D3Xg/7Lg+JABcoEWbJoImzH37pcllDb+t
7yzImUecKhoyOz5Xp2aHGZwaZy1y0b1hPbarOem4opzY0wLY0ILmp0ccBPRwPo2lZu1BvD6uDefS
RIsScYZJ3M5TiyMNMYHsAuI6RnSWx8gULPluNkj+rkC2O7EjgkwLhy0TferK42zjhfO+BohJxCJz
mfuBA4DC3Rapau9vNVVTzfrze1ujxNEXpbChbAsJSl/pmsMdSs1ByG78Qimhf6s1sr7RUEg7wtXG
SS1Km9OK43t/I0XJ1Iu/2DJyzj15GXa3e2C41/E0fKzGGzk+g6N5Nek/rfQioboffJWl6RDNKaMi
pHpiw/BZ5T9+QDpZdEdlP4z1hTpBo2t9hHR6VpJivnbrhc0zvtH0I4Onzsyl+3Tm1bs/nn7LpyVO
1zw+3rpr/7zWu9fJYaVtrkz0DYzwrxSAfMZpSYrkY/8ZepllUmSkRC4sadXhKYxf6LY1R5MR6ZPe
2D0n43lV+CK1xq2LCja2KSCqhPwv29syHTLHEMzEy2ZnUftPuS06i3gYAtoR4kx/rCeYXwV3zY9r
FqdNzsUHyqJm5t1n4XW8+kQOoHtuogk6YBYZenpbRQbyOnNrpTU/J7VCOmUApEmA6TDm869akQL8
iTkDjeX1QNl6OErLNtYF3JOXU1miacxzGlhGtsHNUXxPwn47Btg7Im2XZYTQmDcNA5ONWD6d3/mc
Lf3kC7T5YAdkakX89M8utTp0bJbH8FD4f0DrLRrNwAJdvoAvJGuAC60qZ8pY5HXH9ajct5URiWUd
m2P65AogCvSWcxXmXfkqG2vVD8y9DRexe55c8sTBP+RZJfvZS+Vz0W68mRUsDJyrFGLSX+Uso83i
9bW81EFURGpCS+JmPpjyAOv5hBHBr96nl4I956b/+MiL6he6FtKI+mvGpwxmfTYVO9Y5BTxNO0fE
2FyeZQxLhIrCnAILoty7QT3i9qmgC4Ek6CLvL9/eH3+d2Yob9BLv2i+v0lnJ2nRjE2rwfokv4HwH
yTMvMzE2yBP7W1X6a7syme5poRzS5jVPKaXCskWethoxphkOp5mG0k6lyvqy0hneBN1W1pxfc71t
txBJfZfebERsxLmasgz+YpH5h4iAAWtAnyrtHSfZqyRLAbRk5gvUWpUD4vsPm3CNgP8Gkznzv4M7
YOerg0OEPvNYTxMGZTXs8ErQpRlf66Liuju/woLuBQvbcYRAblG3d8gp2q97qaa/z3YLNYYP3jXW
l/9lPUGfIcZUAxP0KT1IQed7zqSxY4aBGgH1piT/cB09TYX7AgD9humZBrYGRM0jZtCODoUxqMdJ
pEldL2gqI1KZ+VH5nPhjDCIor71vGnkGQ3lD17bWgRgWcfMuR2EtGdFAjn/9uVFatbvo/ec1mwW8
+Fbk5TJ4iHE9oaf0YbodVzroMUNJ4O1xJY8xPlU7jszHDEjMaTS6iLLgfCtFF8hpzZs/IhagdwPb
lBYB5MpS3WApsmglne4rslVfcwhMKsi0JGioEVP0NIIQI//DnwxsWOLoleVCBzgA75dT/Ca/nD5P
edyRwoMZiuCYNAFZVsKQS2FQnCkwq335p5Ll/b40zC+MB1NRx5BRTB768dSU5P8gkivrx9BRWxyx
tRgDhHqYxt5UKuEaBqQR0I2YCv41pNmOEa3QLKVqeYYj5UwVmSjsowOr/3jzbbt9Pddn+ebIqOHU
/hRO/1I1DCZtGDv1qZyW6kyPBzaUSxOd0zLn1WC4fVAMVP/0FNcTSoo+mYsIzabbZ9fhzIbYppoz
V5v2THNMbq9bs9M2M9bg4H4XZdrpMp/Pe/0gpq0ElqAOgIezEz4XQeNcjHuw/DsGIQF+0tmmVBIp
C++6rs2WTKCeApgubX7jHlbD/tuNIZLY2QEBesWeXEaurQcgqT27mizzf1s0Wt4sVD4fsI4CegcM
q85ceJsjYFS0SFEbxdQcRne7yxDs+rE30T2w5x0rv40/5V22RF6l8vfZHxqpX6Um8gDNQIZndq5O
FvQa8sQE18WgXVi6N+PvaHQIn9wF9SeV5AwXVeE37Bc562hI2DPpOUw/tln+X0U1ItOse8yT/Dcn
KyT0U8K8D6IOPkwUsYdRBL17et/B+JSuVGPr0d9GJCUrfH9XTn+3vf+CuC6LL/DSdSbemGjSN0uJ
fgDZge7ZTs0qPgEQu4P0ULgYP2J6wJUpzCMDWJ6Tm8GjJLBsl+7Pdg3X+hlVEiZZKPeT4owzOjX9
tDwkR54j9QpVi85P5MeF3PASJ0FF96tJTsuWvhA3UlR4gDMtdynn/B4Ea2iuoXhTZlf1Ti1O80c7
YZ9JgCKMrIMai+VMuDAzjvgzsZEtHTDMZld4QsCvJFnDvcqY9nR/SNcBL7nol1aa+YEdmpDmtT4T
vRN0sXWU9tW7d9zgsVaNp1n/xjbsNaINkecQQ7rN2LIe63XiifXJmDP9w7u6bum2llYqWeYM3GEa
41oXDmQjFGjbG8ln2djaz70vLzPj8YRyjoCT4//ZFjeZpa6GX07dczXLc8CXcr5e7+iv4nz5N60w
XMfNwba1aCwmzGuFcYBMnn7e+6ilCGgF+dDxXEcAm4ZzFEv7oliqYk6ke6F25WjK0ZAyU4PClFgM
WLFTx35UkC0XMmNyc3qUvvsobLkaaYsKWsd1SYTgvsQLifSsBlvGQ7HgT19w97A9OX+EBJ1u2XIi
89qrBcuplmh4P8EGAoNWGY4EpNU48su83X9mrrAAoOVuyk3Zl/BiCmNZOmCoGkhXUFogYvJV6Olc
0nKx5FCKia/4e4xobU17kPeMN++KbLVZjvulCsuzvNHNeVhiutq4/h1RGeRc32DVcnTHQPDlCe5s
plSi1mfIyM1zvrcnxyoMDwUsK1D7fNRrtX1K/KDkKFIG4T9IYDsPdJSYdnf/OEYAyqMoQDSACudc
Iozx4KbFgLNRlPk8MkGoZ/IAZK5k0hpOmqG4/utyScpm592QioRaAUCeVKaeCyGYXJi7YFkLi9Sz
UkrvJ/kOIkYktVcNXrEIrV7aLHI7bRcW9CO30zV33kYt+ddMr26YybNRjV4pG3SuDceykmpTfeeu
0w4Upe3v+frbH71dSNaAkAiP4KwuGtkthUGmKRviW1dGN5VUS5udSRa3wQzaNU5ZHoqYW5kz29b2
fkWPqwmjJ4gJexF+KZMCdBOjFv3LhFYHt00ZcjP0j6quzOUsCUea2/ZLSDQf54iGp7MB7uJxqIw5
H7jqMyR18DslinaJe+SYuqWHLf2enKZ1L4CVT+AkzRTjpdwZZCc+18EEiYA1tYvKJhBKekSLijJY
vaf6QT37s4OGrAY8LMaw4ZnjsKqQ+44Kgbou778ozRidp69nerkB2C/MA71BMqZCNkJkDX9t5XPo
DA6yMOCKEWgoDymTm23VW1OGpkZdI2vFS/ltejVZdEfsFX/ZBWuPr4AOQoRcC4WyUc9IpOpB48QR
C8Gs4sUji8mtm78Yy4BH33doKTtuWECK3QD5CoM0mIRudSAoo+MsSOJdcuLywtHk3TcTR/mWLwXJ
+d1Cx6YSQ0PDzMSSYg98tso7i+jfrBAZ13xeJFc2lXy18NX0debKJw/MZZqVFq39b5GF4p0v1hhz
6kuH366kj/+ZzPtZsIyvs5EXdG6cANSO1BTotMOtvpD1QLcnGMBOLFZVORenz8/xRAjlMmLmyXiO
lkRpxmYCTJJXnRawcAMmuTvmbS4BRZ5hMDb9MOXAEdeYHt7VVl1J8gT5kqahA9Gxp4noaw6E4ckH
5rlyP2e3hQouqOcTDslAWjKonVzh6fE/MrzEU8n99M7qV6pebIsuBaRx2jRlKefrMcgrsPMeFw4U
9tcws48c7da7BbaPvpC5mLOI0sD8ak2kQvi6Tn5Q4Lv9nDfxT3124tknukPQrZWaA5Xoe5PnCAhH
/ZIa0T9c/9rMk8bkCgjgvj4EzAUKymAHJu13iMjl7dgAy0Ro7ocVg2/eeqKNmbHZuzaZv/kJDJdf
z926BdlOsA14Z4Rpw3w6mr3DdmAFudvVSYlw/fnwX2R+54S+O2+Lns0eecCjsPgolURxrw2S1SCB
hAr8AlhiacKL5FPfqfw+cI7328pLxvQyqQCKJXT5QYkwxCXvslO481w5plpjN3mmCkWZ0sQn57v1
RyD9HH6lNQrY9rufeSU8SxuuKCYbEi4seEYfyKCq+ovcRCFh27OfGeaMOu5zWr5tUQWNblFyo0jn
zZYnqnC/tmxUHIHDKBEzz50ymKZ+NDLDzzwYg1rfeUUVm4rIYF2Y9AYtSAKMTD7WFGhr9j9dyeOL
gvv1Rqxi/IMcqS+W0efXikgFtNpQOsToPBSliE3js7JUj9gJFcv+OTGXa9I9o6lh5A/CtzclS75f
KYSqQsBb2fg91QYCaJCa3FL+HrOoIr3YU57GL85t7tZ7/pPChZs+7DovjCo5eTw0ctlCjGTA+IoJ
bRQ1WWEma/TANLSnC6u7QTS2XNL/6usAquXXPRie5G1c0bFK9FWJzJ6qNzI4Ak913LwPI+EGm7hw
c2CMMOJa8O8Y9LYAbeqBP1ayaAKmLZdAK2LuIL69k/VpD12RiJ5WVe7lHu3sbdD6m6jV4nZfleWM
K5cAzuqjY64nLYzumRRWgPhW/Sx+1j64Vsvx/DC6CKfYZh6DPnQqeUKlMiJuJ0RZq4BNwC6GX9H/
IsKGP/yYD4F9mXHEab2m7d2MG9VYNFXNcw60Cbjt+Lg9WgndQNklv/58ZJfdK/FpaNJxQZMkOwyS
M1IddcHmUoqrkpgD8Ms/a7pTkV92WHY9tMoFVRG/Ufa62mTe2D4NcGic+DTkDSByIW+CyHyaFFi4
y5rhjMAc+5yDMzbL8fz3Dl5gAkDHvxdBSF5cCHRoBEnUn+64BsyJKjSaM/9tfaHFKcwkrLBw5DIu
zWtQdLMs5vY9bsxXa2FCWiHavotmwS/kKIqPo2siAf5EUdaiFxpQhXnI3Es5NQqKBapUue3Z1i3P
KhVupfSU5A3TcRUy+eOT+NNjlZq2PWDk+/SA9zForv3IamRQ3/Mno35RdlgotTJfD+XiZP5awQFx
vDe5ugFyAIx1LgI8q2SOOCQy/ws9nrcaZHrenvb4xuoCn33PKcQSwMfhQa7rGZ280LfrHvHuQUBy
zf5gpeI5nPmoG1Wz1oVdwKA5wrdmoH1e8Nc1zL6lJ7rcSdoAG0jjwyL5fIZj+XYEhbIAvw6UsJyX
U473Aqlt20PDYAWzRQvx2L3UyLa0csFyLNN8CmlPJ+phRYwNrhq4mLsrtJUaohMy3ACH3d1n8fZu
WJzufpj2BLQdFBxpBfzD/OmjL+MhkJ0uo/K1VDL3wXduBj0+R5z1ZTKUEbc9qR1jBCdGJ1Itjlb/
H5SPlXmREV8UnQIRWh4LWp9PXOTZeK20nS0vKdpsbrh3NTsx2vC5g5mBJp3R9f94gFe9LFaCEWc+
p0iTNrBZ9d35IY4jWLtcMXUElzSyHCrUYbLSEteyX96qHLjaZsiWfbiXoottuV0Y+kHjtCrvvpyw
lNTMrJHEe52Mt0ljG//G4blnzQUmwMj4AEfFRo+63tmErI2XPdcjlNKOZpzwjHw6flmNMQc/z+Z8
SAzzi8RQwK/dl8SaqyPf5N/6qHI9k6IBEXWBUin1cVz5vHBtpsGTedyIPt3HBlFkWHnTbO6Bmfov
DXhKdxwldnSQ65Ve7X9dYDk45eXV4/d8Q1NlI1jNl3gVDkzKlW9JAFe6kR0jcdja4PzMJds844eT
8XPewcxgDSoa0zegZg2rLpQOa5kEDnjoKW6Gy8TIMRW/HRevQR3gQfvHeOpmnFNHPKhHv/Gu+np5
1Ji54hw39REBIa7JwS/V05eITS8bzIRnxJ0ZNuCk/mOBAPkg/j33xkXPygD80u3XymOISEddSM/t
i1EGcS8hAdJaogQAHXEc8r7FIO9u50Acor3ZLbjSTmYmE9WUqRAmsD6v0cHdvWEOtQK26gFzX0S7
dOuk1dJL5QIG+8vXXl6SSGrd+W9mj4GnbGtXY8+slVhya7UwQzlxod9btXz56IonFLhhvDD5wFNI
3E87qlyBEwDnC8HPcP0jm7TOSTq9uhVlEvrW7JxS+fHTdIa3eNEMj8Ut6ejvfk+nq+KwtYzOm6aY
lEGvO7uYRkQSr1OVPNlPf5Le7laaLtL8EQAyHLOkSljuw89SWlcV5texV02HVnozJiy1CDn87yqf
H80j3JOIcGjVqiL8GpQJpD6e2N/toBzRtta5Ak6275eE2ASmgqvbKMbecE/9WPixi5YEcj1xNLw6
A48fp423EVoNOq5yS1q9BuZRDMQY9Trtc/NJ4Z5KWIoa26YmWv2LhoV2LPyaHFEZ10jdiziSr0yd
x4JizdpO9lYOE57BoWvtNl9oPAl40iKSKcFDvx97N5VGH6kRngGWUl7ZYoMN2sjg7jEJn5rl64ua
irNHZ73JiE8OYpEw73HCebQ3hcNwBFGeJo+ZtsaX7eVP6Ii9dn2nKIlFx48Jq/NIhMZCdn8vdniG
oC7eohxp38bbbZDOcUFA0U+mRjh9ahXYlQqUHB3K15TOFxQLOsaU+n6ZNhNJ3sJf3PWzCK4/e6ik
Oc8+e6183/Ou6PDnxM3WtBkkeKuGcCCUSBTAXZzoKzirkoAtLBa76DdMifrcMV/UHZh0QOzuz/0g
k4M2QwzY/LGh3rYrm5PDFPB/aa9Dhjkd3xGKGSja6nVkeHU7ZgSY30k3IXtHEy94PoOW/0hW2tgt
sWrprjjZNfWcBMzX8s5llmDhureNM6Xy2o7kx2c7iiozbMvDHcGE9/HZFbcmeDV6qKDLUfV4YklF
zZvpHoA9Ma1L2hFK9b0jIMHUXLlDKXTWYJlZYNqCkuLDb6WLIIx2V2XxqKtB69BoavnvBA2w8T1e
BIYbFC43k3PO5KuCjNlcrRlIDXKLNkOn8khFPHy7HaJ7LjzTJsgHNk9g/vcoxmuNTxFNmKeFaQCN
Bz0CL472dGSqUcLjdl3/MOdvuQ2/DeHK06us6ZGa2vgYRwcP4rwR+5CGs8pVSHYr2c9t8CLV1OZ3
0+IBx5H6exFV9zFJuX9bVBFldePfREubReCCtSq9bJGZJBQ8NoGIZu9sbp+yJS69VU3rM7UJviAf
0q3rHfMPiUD8RC3tm7VOS1LoK2Xb+uCU0D/Kb7aHj7tQhRBPX7foovMwtLjjD4xGbqFGghg8yvla
QdRHRVroqfThwf3qVi6D9hV8uXWTdT2T1H76/JN7rsiKiF6vnn7f0sILjVLz3/dTygZNukzEdwJT
9fcTieGNCH0lb5gVtznatsMeyQSFrwr5fewL+zdXeAuCq5ToqImQpUu48+NH6mkY40dSFBvDnSsP
xIeLQ6VD9ljglBamg7sypuvomBFUqrsq9rx92Aqw1iZPbBq8ogOGDJNVjdBhKCQrpni92Cz5zLe7
LHL+pGiJjDCSxoLbelTPiJi/5Q0cyXbChgMeuvYB6rTFKdh51yb4h8w1bxuNDimBhpmu11Ewt3RQ
KiU2UV6czOXJ/tMHT/7qCn6b4ALA4zuwXKaBNjuYFGJWgJ2ZSeIdXfWut9HfKZEBnM6GEC9OpN+y
1elCcX4B3bjhc2OuFJ/xHiwI+cxbJd0ELqMZDpvAIfbYHT69fLuV9t+PMttNOK132w4smFowE8V+
jvJoOHncwwXou6jjkx9+9Y27DvaiQGTqFr9RpJKrknRg3aVCoHVlXgE+kWatN7MKnyAWAz4xX1mW
9T9Mjz00PXO0+YEn2+MQ+pMizruiUC4niSWjPaAax3iT1r5HIL2cotDTnR/ipIiYGu5cxB1/fJDb
2QBzWcXl+1qHqIUNeASfG4Dn7g1S1BvKAa0WhhXJYbn8Nyk5iLoWMP2AuMwWK7oXiR9HM8Q1QatT
QqD55j0BiLXMya+0xGRQxbFTaA+lIX4A8YrEgSl6rHq+mluNiakyzCEWQpkM80mICoaTi1vlv/Ty
3lRx0i4Pxk8k80gz9V3XY1bEirVsX9p8PqeE/03aLCHJB6BxD1d1fh/McDFyAIHE2pdv5SeoXnYH
fLAXciz9Zl2TXXZHrTeVuWdK91giqq+m30yhZ7wjyVnMIf79vYdAeMtBMllkj3unN9YLaODTarUo
Z14Bc2/siU4JpOqVl5Vpj4VRXH4JtxEqlpydAM4jTv0JR+DIfILzP0/Ump4cnDveYMh9waH2jur3
GfwU5DzOH/bf48cBrwBvl5XUHaj+dRRa5M8KpLXpNoJh2AU1HnDAw7Wb4Q6apB6TLvfPrjS8ep3d
g0als9hpIpnVUScLkzrlzh9bMKo0tipLiURdRKs2uwWxWMP4/+dn7pbcSALdrJ5rMOmt23UnsDS2
WsJiW424XQjmlTp+8yvaARfw5kqAL07rwENgTCRj2Et8ITZk3Uuz5o3IHp3VaShAtHnYnwbo+Ohf
aIav6b7uPJfT7qyTbkLgrjXSvfWfu3mI6KXQ5R++2sJ9IiDQXCIQeJl1u7bRLSt0ik1HHNWFh906
0Pso65UMe2di13YKZFtkiJZhnxX7t6f0ovHgmh4HtLpVM2UNAnt7UWy1oL3UQJpFPJE8no91SoLO
7oB33yB0mBx1+NIa/8MRrvQylJGBLUtfbndrA7c3nGvHE8yCjtlqSHxz5Q/AloyiJEylOhBcMKnn
yaWlQ/JbJAYr9yrW/bAOmEokFiL7Ob5HQ+fJOSXAA5ycH1FiTvE72UAL/Ax1SITsC4JcqM1u5DRW
F9c3YFWVZFIzwfQd7sB7sm+fo18qrUzjx+X1e14V25C++KQdXlm6rQNZFJfeW3zPA49Z2n1f7ZaC
MTC9hXeOlJBJe3X3x36WCbk6DPaHSE+yCdIDnwLxXjwf6fzEAD6/KSGMO5ygDM/ugShROVpY7RaZ
xdTYy/STrKlRbVFzYkCHOLuod8UzwWvHrlsJaeapUljObgypFGyeyWDv6CQw29RQr5Qyaksy8DoU
Eg4LSxeOEqXnOFq2Mof717zKM8eQAt/nk1MUCG54B5umf4jPFA/POc4uxai4ViEdJzSMnK+3X0MO
wuHJKmrT7ouafutKmfLIStcHRdd41LLkoCrBS5dxGW/g2nMlzZ08vixl7LSGCa8EAKXcpKxsFqi/
Zf1wq+J3cWD19TQqte+4zz/y45RUKRAgaT5VphhGeRWWGMQ8/vefhknSPmjs6tXzO72Al9sQ78XK
LotdHNJEmaFsxom5jMjvn+I0XsDUwDuFa6O0P725TU78p+ErhSrcKnQczIP3soPN1wDpgaBeySXc
+AHGs9FmKN9JE7B2AMl32qPxKdViQmGThaAxIh7XwmtyfcrXm/4IKKCKEKdX+nFaCdmRdTM+Z6cf
EVf2ntmFnfgRKZZWrGucSZvXXdRfBB8qvXmBByCIK+oMY5cxlquI4LoxtNiWTCbyoZ1zDyOShRRe
CWy6eZ6NgbSSOT7uIjCCphqCx00cNhExPpzRIunQhm0jltQWVF6CwX0yrPxzthPhlzHfQaCEsa4u
/SpfleHry4/L8SU/c81CCFKNAFBcZcuJOrwi4ayCB2NcT9XVv4mVzD6a4Bz06lyZaNMCLy8sKKA6
QenJW4hjNhHkU/W2IrsMHzfVAUa6V+Wx0tbknWv1+uuzgAzWevVgBYAbgkDMSD8//mjHAyQXtGvx
bJbN8+Ei2z/fI62/5nehzUTWNeHLH2SWUKzKRUdL+9mu+nR+rMRai5lg+gm5NjKBQ91fqSU729Nv
aL63KI9Bo8lOhtdxtOsCZ9EyP3gBLc8yMawL79CDCR6jnIf2MVlLveXEW/3XkHYY3UHhUWygqxtL
Y0hBkq0oN1XoPG9jujuwZnEr4Zpq7B2iQWCoG037ouLVNHmatYoZi3pIzZayNHvhGIlBvt01iKK3
dYibdY1IIevYiAtI6lZBWT95wIHCqzJf/04Q/kRIIxQpbWyMW0t497s7lfNW/Peb2jDs+nHR9+4D
fNL/PqN1a3Y0gvNDakjM9t+vhA56eEkySm1Po9xnJz/JipjRMKJS8gFIr9d7p7me6UGdOrqd8oee
Ea1GzDJRBKxt/DIwQk5ihsWXgf4QEr+8qQvFyMI1TELWE8UHoAD4DoZTGS0mYMfzNJVwen4hUChq
ziHOej1xLlKuTJ3kkpVI1C2T32TgyDtfv2zMgDiael9H4udj/IEb4QVJ5HYQi0KouPS9ZFP0f7pl
CBgs3pa/1nJ9kio535cXq17VG1CtD/Za4mfF81v+tZW2nshbrLe9AZiwEq3hyXQz7xbIx7iewSf5
iSyVjZqTKXN2gHugfaFBFk2Os69AzxK+K+HBlPFlOySOXpPZC5PZZNxytRgIGKrAl3Yb3HIstv/C
edszzh5s4jmyWTQMq3IxZYGyMwzGwGm+CPFrQo1lSKM41qWQfFtUp2QVheKssk6YOwcYqlLS2tcT
CWFwvbSpzWxiCsjJmoYa/JOe/DOEbsvR+srsafk1YKejZdqG42FS6PTKOBqiR8JUm8KWjCID9Zh7
ZAbTEohooJzBoOs/hPZF34L4cZDrz3UiqsBJOqjNWc8//ZcIMV3WrAxXMbLNCpblN3J25OdV2X8l
ipDjDcYoNPc5shj5TmDJcZat6E+mChd7fjwc/JjUyaXw3xPtmcTRTgbRakTAHrm5VzTHIGnP95g8
+1ExnobMkZlzY9LJ7Wi64pQpT4n30gV4G5iip9UzUN42xzk6hGV/BVlvJ0wCJYoJaYF8SFZK+hRW
w7Gw//n7gJljZp+wf4WIRCKbpTZHQG2FoZrrYMTi0f1XD/qmnKGDaZMS811zzn7rma01UQonE4yO
YzttXSrYCMl7IvcPZ0eNZKp0Il/0NYO74KNRlQBsDz5xqRXb7t9H/HBRemD/c0ugbH2Cu1/oiqaU
K6tsYUZsu9mqG6hAmtz8hbr5oKo7YRpf4PokWffG+BGGdtXwCAvVIvlNPTi3B8aTfgH34drRzm7d
oGPEVp09r3za45kIHTrbslIulbeXKX4RjHTiLRYgRsau6AOLbZ4ajEoSdu235YEAo4gDlldQfUsF
lL6Ryo28Ay4nz62SW3DN0QbIobUwlVcU7fyj5OScyTG/zvmLxhKgnKaTSlveX7nNOLsmfGoq9lOc
492CKtqcF7qC/PR/jvIbzf2Eh/SOhp00PLPrNm6BXW6kcEsCag3C1I5TOEv4EUDAG4Auy5GuZ9r+
1nbO/HuZLHvvvscY8kBH33ccEyT1jUUWz+b9elMG+0BIm7hNKKk5Morc6eV0Gb6J98gkQI2DjsWH
DQF+R9QnNntEagIjKn9+DJcgyyVeY/UilQunNTU3nuTk0cXjOO1ndChFBKLyaw2/A3DdL7JkwNJg
wyaCEVWXiLmXG5OyQwcGjqvk4cB++DpNFLynmhB5WRWWk/RXoEFnSdIr6y2cZZmDIkaEXxQKKlWL
ZstAul9bTglqKIApCkXtjNhaRGJ6eqGkoO94nsI2h8x1DJxlZ3ivXTXADUC6vM+UFpfZiAvhNWwk
bfJiyMp1TfgCn1Cf3XPMD+kjfJQkAyKtm6tKPv3sN++2k2XAx9wHrKK4FRU49xyUnUG746kvDTx+
QYLhqBJ0stOlQyz5CmoWffFSrSlnmIAoSmlIS/FpUI6u1f4CAFsVXtHPV1sOw4kxeaj3fvz5ptmw
4kuVKFnrE06xun+7Mn4XK0Yk2C5ebOT1LwPMwVadN5iwX77sJjx0TXXlqLeX3dlQIZQj25+ORCKu
ElMvNHA6Inl9qzMELR0nd1VQ6yVit37SjYGetJ4dUjZAML5p3wOnj0zmQ7mJ2Mz/sh2GtU3KEWY5
NUr7AyuWWtE9Z3ANEAVAX3knkSnDJmxumVdyxPkwKbBXd1ztnqJFP512q7zRmDWtjJE9/ZX7Q3o+
r5nDUQOD20bpwEHO9AQfXeq9DhIBBsfmuGrcEWm2BOZG01oYgRoaxzVr3z6sCu7oOjBtVEvZXtDP
C5VQ1p0uKLYEw+9fuDTuqNA/lFVdHLBS8RbztfxYHrO/sPH520DZfvWYRW3cZ02qC0TByEG/ebCA
gGXxCI0+cExYZvPpE+4VzHx+bppjktRa3GwIOdb/U3JH2Gxb/8L1Z8a4TjmUW3c0VxBSehhSMmpN
hSqmRJPunXlYu8aooXqwbQRmjv+f3ToEzwTed5jLcKm3299gk2hC2dutWgwCC7lZAEayRpkI3tAO
50xPdUesplJ9y3NyiPgt66atkx7jhCryK4Nm84SNO6vWz5WWN5teX5Ynvk7C4wdtTKx42/8RqyhG
G5ODuykdIoN8hiu9BGDn2vhHGcNZZAM/63UhLhPGsTnEBt35tlQYA1HKAXaCLNVcQxvuvZ5uATwm
Io9Njj+EigBMb48KvwkRgeMPwsWi7Nno4pB8ZpxB/fndZgZ5PmTkmJPGr9SyOsE8M46RSJA4Fhue
VzTvxm6POnDJVIo8Ul8Pkf4QF4sa3NPEdsfDvePE4TOv5NXj8qyu8cE0Hb6GoSNBkpL0Cxa4Yfgh
I/o8DAnqdVk7palnNHEl/70Dsql00dl4AA0f/3IDD0fjXPQR13ciHa4IhAPrzkFwKD1gO1uvboQD
bvHWlmivk6RFCnZszsZERIv9DyhyxhqKJqKsS1f1VPwjb7WPDqGnb78Yjh3uTARTNMQMCvVnHipS
JiSGAPKp6K9K3+0mJSCnGUlGrlRRSOjgZzqH4fjVQppK6OHfESfg+aX3CLQvIBoNfBm2EXg52U+R
QyG6eC0LdjiOfelZsENA/oh49Sg/fmjldDfsv5xzRVKPZiVAITrOQDW+JboGYjcwiHdUq3X4TgeC
BrZSUgad01Hn9lYi1SrW2jrFR8YdrHFxywK2IRHUKqtXo7j8njFRe3hKxf85KBiaTFODBg3HgdC2
UsGByE9l5mFUoVEBbft5iJ7vmseaX/hJFFB7BgPj097JNKin1j2tQMvFOOoponbXGtWtMQY36Lvv
P1YclqIpw9bWTELl7DNEb9LvI0vCmhFB5zFEkGZThbXOEJc9ReUOftTVMBWqLt9TQ8py+4sA6Xct
nouYH+axDFI1kPBKjhBtHiJ+wwggr1bmOCHT+ZEreWgTh2RpuhahaoqvzFJszLPY8wXGFP9LRrr0
t2xpB7OUCMQN6ag2VgKp6WCVu46Gc63Pj1tb9u7YBWWaE2WR1qGhktfvfvWOEUSp0wzxhMEgGdmM
jaK3Z/H7KFlSZ0q5Iu7Lkq6GE8JyRWp6UKAz2NujREObNVbOTnZndGFQWvHmpcJTwm6sTlPgRSDp
ehFoXlFyiAEBhOfEbs9lWCk8yYybs38NCmr1KNJ6cia5hWcq1db1olZcl5vh/qLLE+TykTKkQmZf
raRg3eLnm8co9wGshybQ7I4aOBjOIei0xrVDHtducFwnKh9gmNH8+Acw2gyo/2S3ie8WIfUiJ/5m
zIrYAAtuP219nMW2vW8b60dI16laKQwdbG4Z0FJzvEcE6xvMQP+GrGtdGd96UdSAqjBJUaX7s6j3
kceZjlTCL+wQW7+H48C3tXMndo8W/9YTkZidKLDEeD++xdds41S6WBJY/3YTAyp4Ha89v8cUIZh1
e+zRxoN6PgM62I5PPVk37pBjfGcHvH0yNLe87z+GRY1w9w5dCLHfw85+m74+f7rWeIyajLHidQWQ
yBTBREqgRdlPp5encZEktmvR94gYFMR16fZ3dlLGc04YxyuwqNBZAjsiZ5/x1pfUU6UGgS3JnFU+
CnybYPf+OQ==
`pragma protect end_protected
