// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
LtxdvMZ4zwmNGwbit4XV0x4I/rVo7OSrHAsi8WMw3jgM7f7TTx4Cp/9ybIjaxfA4wgO8l4SMCoPq
2gTrZhOOPg/vfn0tPj2uiW65WhYAyGtCoRAXWRQTj9F9/4pUyOHqSeTU7eBrv/du3m2n4D8TrZ5V
hHFil6MqxrqBl6rw+lxYt7yIP0O2ycdcMKsWV8WLj5EAmJ9wcVsHEQyDX1g3KtSPCbT6TBsET4bF
i+l8M9teOZyOJT1JJ9G6PeOqZWrhxDEd+ZMvcQ1kmyJhQaIieCOYOlUvIaHm5etB+7ojHsmB/g8h
OSEKrXGlYOOKdEVK3SUQxS3X6NU0LNrlHyJMnA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 17376)
8YP8p+hdUdaIwWCd9XlNh8wRHpS/YhvGTNvqRLBU36Fv+uKS7l7YHuTgbK7AyMh4blcVdbV4B82u
toEYeKbhkCFB/SZygyRao2G6M0qh5jZn7hMj3zmLnGlsDQhrW7Qa6lQbD/SHEHkRkA7DTyFYLcss
dg+EQ6Th84ocKduHLQSy3BqX7sPmrCpmbZl3J+ZxSw8N0316iCy7o8ru8Rqmr8+Yf13q9WnU2eX0
akRAqvxeW15WkgXjcyb/QyfGdFt9S1mGILxaKht7GXG4Isgmwpug+vpyju0Av8JijAUndoO1p096
or+q4wnGM3XKjCtVFM8/nKUzX+ZM2x0DIR2MmfjRRHyblcthGx53kL0YGPaKI0rN0EHKfrgkOX+4
hTjm5RvdYP1jLLnwG7J8JRXVsoxknf4BgnaKCO4bqGBFgDgO1hYvbusKr6ojhTbW5b8QnuirT++f
Mz7cRmKktsaLTkss1gUl635JpDsW7tIzk0dFEBMMcjDBxhEVbENa7vRsg6tzSF54gEMdkRabVyjd
/wis3+KL/ZiEZKbilNZQgkQNjBuAMtFHaVlTbf+0+sngxjjk12sAktIVcCfgZXniP+M4ZNdAjymU
ZwC/7J+SdRyUSiG7PPvSo1epIkgx9dmdzPLtbwmlhdivMwWU9ukWfR/6TykHJ+E3j5Tx10yrcjXp
EF1mSer8LbK+s5rAkHDGlzokcannA6p2TZJSfd0mZ6ZduE8xmfFmoXjkHm0UqJ4M1yPqA1TmvkZO
YQagBxNXTM+nlIf0oLa/6lO2WMzyaOvHjMqrLS0T5F4+GcZPHn7T62bQMlCcBJFY0JO1RUyzblTk
RE469726h+7dSlpaLEbXnuae8AeiwWXHMIEvfvdP6wPM2ALGX/bCZoPkW6/CKjJnr8msCcxJA0k7
Wke/1dDA71jcaCB6XZ49oyLIDqjohNscI6K7qPDtobwPNHbOimezEoR1jeXJw4KvxfMAd3LEa3br
bGKWQ1tXGDagW+XZ4sJglKbc6dk4ght86B40PSvq8LUMrzcrKCOHVyHvagkGvmz8DFP9KeQtM/35
FyhyWjZMhUEli/peSbDyPvT3JZFFPHzKJxagWxEDhlUN4vc3WtkqgwReaLjJI3LL3/d86WYr4SLU
+zKRbJEXCPoznrdBgaFTt+w1XRzTWWnUM4yEr7M1h6BUVYzNu+GA7CdVF1xZE0fVNmAWI/RBXvjC
Q9Duo3pYlU+ATp+MArjk00umExoVIjdZSBzdgLX6Jgs3gswZbjy1JADv0mLmPWP1be3UDYG1l/2T
qzAhBRjJniLUIudwSgeOh9Lll7UMrEyIaqXcNP0SOKi/n7WLN6WJk3DiFhUTVXiGqmT4bULil1Xv
ELjsGttrbnQC3V6v7jnR+fQaI5SR65lxiQWp+6irbYGDNvixfNBHc7VrMnaz1beR8+KDc3Hmt4QK
28jj1FqoNz2aU8ot8TAwzpee9MSzTI8yLVh3wkGdPiu2NZcrS63+4oCbaXahtjkMAAJUKvxt0QCw
Lc23pdz3Qj6abaNqOH8XCa0qN6pjAfSBHKTbD5Bw16YovKTEMZUx6XSoBlTuU1IXVD/RVMVaPVGk
B2BDZwP+biqzXeaRCwCfArO2zm0tKFImQ9wqX9bbdRBwVN9+t2DQHejh5QaF//f5rZy26CuJ5xK8
9XHCEVrOQOZeW4nukvfWcLqmEGSC/u11FroJtpu7tl8I4YFWYQy2shfwJ1HIPGNXUjFYbZIx9wYz
YYE+YPZ9FHL4EqRLnIh67xQ9kh+8rxUw78sXTP+wa6XYKaSZecjhQW0kvcJIUEkfyF22coAezzU7
I+BdtPXH1bQOtWqxtUHMg+OlwKaa+tKd7KVoxXglWDFesPjkWnvqpuBQ3bGrjt7Ecx3zccvTFLj8
6YpfY2wz5RIPZgkKKtvuUErV94FYX8VNJ7UmiVS8whyKotyUo8Ep0xqCtWFWw333b5b3PrOPurL1
r4gdz2ZNBoi8OZTqIGtwFpr0X/B6QZOlZ8jxqT63AGPs89I87lvEMClYNTneyW0r6CqNf4sLi/ph
0+BmTRiZpqeKTvD2OOFKfZwP7Y9FZJf+vonULnmZrpOjvJi7c4pBH62zYFgmWBkkYIxI7sUCEULF
kUejxHiQoTUgHpxmI5iCJWd8UkJemM67v/WryxtphycwsR2tAeLvFsoPTAuZNAH4WQBR5rF8oNLu
wOzFnvMNtWZDB+drNjZE4iLxYDx6VEbC92FfbAkhnuiHfeYrNmZyz+jUwhFKsJHa106NBatX/6CA
H1TtC9ReLCvJwJInUcUh9IHL269VcBBySixCF4q5HerxqCpCzpBEBnkKngrg5D8VqMF7QUYxoZbq
KZgi1zB7AS3jbcRHFQMc7aw7axYZ2BH2VODS250/WxoAwbwst30cwmOqrWOyY4SwzL9q9AiIzohC
wLvQakoRoepIDJ4P/K/20U67bzQtfr0ODmsnyfJQXZ0bxn59mk7vcc11zJquLzmJP9RKcYFHaQLy
6pfRjVymy6LICCOpPD1UVMg2dSF6XPF+VUOSlw3IjdvuN0H+77wdvMkZvhOZ7vAdCp9GEdkP1y5c
jRsXRIx55hgJ3otGZTIVnrykmulUMSYCMik39Y9/wx0j8HTICr2FgrhmVFj9GTegiaj5RhtyG8dE
wIJOV3Id169ZEPwpIVASmaNxr0Tt06rYoMTmBP7YCq8qMbDzoll5uoHVzaYZoA6CRKD38E672MbQ
6Ve04RyBC/6+m1GYHD/IItIv6yVuvVUFBy1YjlGjHXzT7UO9OBomA+6WDtXybb6PslSBOYWT6o5s
MEknh+adDY1pOa574AZtqRSPmNV9yKMYHiCIwfoqHQkU1cH3NQggLbPWDhBOjiPQA5KpgYolPuVR
/RBhBQtcd7cONcQUI646SLaQWIZQPLONxtiRFc6DuqQ9pNweIUMy65fB2YCZU5NeeTLyk1EYRmq9
G/2lpnEOWUhkL6xd9W4BdftL39ztPl/L0+owpUecMMmL+NeG+dgNYrqTlM8lVZeOkdYmnQgHOeuZ
qEpZnv0+zunn5fXBA+d6u6fWIKN1S6et8zZVTUfHPJiYrTeTWAVB81D21xkKuoziGyC8MhHDjaYx
45mw+8u+z4rfpSayCxIsVkI7Ys79VAJxURYFzqOtKL4ZZwg/yplVpPDHF73KC4AzGtY7den+nojN
NP4R7+8511P+8K8zPO0TIBTW8sqo6JKhg/ir2QJMmg1CcPDT7SX+QUmFozo+Gzw1vifn+l/X3ezy
Nxe9EJPZyxpcb0R3jJAZ5P0TyoJsvuc7PTefnZ+N4K6tS5PxS0RTpHgGuw0CbWeF6kb2lNzlxb12
RUCQ4ZUs0Wk6EnY49cUDDaPFbWPsHSlTOE/HIgfo3HY1yNQAK784L/Tmprbb1lq+gFHQRcPrEdtK
TuuZX4Am+aoEMPkjstylJyxdOAgSV8Z9bNJUwclfZ85XVJR1sI8eW6odq8cHRnbLKlQ+tZqb/x2E
nhFOxkeLlRZ0yMlCjbtkfy2Q48uKJYSmYYn7FB789RcGBdN0eE4H3fa+T0hFQZ+CuItt13n2rAH4
SW2O+wZwtrv1xhe1imoZDA3E2Qh2TH7Po2YUnyrnhBZjTtEmUB1r9XIo9GTklHUmXEfSJSxd7cKc
d6l6ivH2kbFPkZnyAz/9a1YSDMKtijalZzh73crfG7GPihb0AZLPHEjvn2ZLdly0pB/1BJRM1qyF
OgOOIE97snmxMary3L46NJ2XYmQZr2Wb8yYC3JonWpVxgIU6vSwIfmYbMJDHRXi5knL8U2gC27FE
25lHlypV1aERstzPvAsWnEl3AyY65Lgh7H6SeFjhYFaucdPLwTzmOHr0KT7nbGi8sCsRLkj8k8zD
6JOpFzdub/JrA4qa8NdEOwUeRYKcZiftikDkJ1kLuGz6aIx+S6Rjd02Sy3VTXKWT3phq5Ql9tgF2
5L4z5BGB8ytAPPbiZFpzr/XGGFtWjZiNd+2Nas76kLTMbQgi1wVFXbSFKJIY6d/fjI44yNsrGSLV
PefcM3TSaVBWjuiNn2Oehk52x+lMY+4p5Qe8gkhtzaAUrk5Zjtypr6j1ZTWXibcFXsR8Zdpts3zr
n1RQQvRZOj/GkdlzQLirsCsAwNMI/8aeFcKRnPC0QuYdX5W22oyORMRQQASyWUwt78iF4Swddn2J
o2BO4Ulcyb18B7AMMSCBDhlx6iXdTD7rS32+3N3DMfHHaaqIZVHGAkbB05uMdeNmPqPFs3vZoZHk
LO2yzvPnFLdnBoG+6OhHZs4boRfhZIeQjom8iQ9trGF3kQ+bxYOtFMqLG9/q9tpvkNlss0uDHExk
r5UC5NTMOGAi3hndJ3zXyVLvP3Z+A3JchC0YtZOdZ4XI5BhdpRmHOn9goEjPEZHu8Is86I3fpxLn
kv/kIxzAuC+McaJWZrW3fP2q4dCiff0LR25mI3GtdYgJnTIYzFiLwt5YR2LqYMix+GmQMXh6l5cQ
7jP9i0gmWAtL1VgCduQMEbEyG2oqwZvBold0bEY0T6a34JRXbw0xXfa1dH1kYAXDWfWW5PxpmEHl
8pOuKmKaYIZ1qUWn1NktreGUjtap7pBEijRg2itIlqT1R6taEf0Nl8Qe0+rKpBXJXO9BsUXM0ECW
rofx+V/Tyc+2bJX03d5HR7SY5SBpQV7kAP90aQATLtObWU52VL2b1k2vQImXiuYKYwxm04uP69R8
P7lzyWVn3yseDNYFoSWAGkVhS8hzNdo5gj1y9MVxKECi8TAhuwE1Puojkp/zML/VBsVtaQLw/v1I
jP6B64bxomv4juLfgvPzo9Q5XNQ5/LCzV1c8GEdyiCZP9E2cBWp+/LEtEkUyPRoaCiREfQ8iVTdP
Q3v5grSVhsJgm60pCuWXY29bs7/WRDjhhTn8NnqjbmVKbGrFlRbpcLTowAhT8LhJ97isWAlUcM84
cR0qDQG00FhSfQpZimJSlfjZNTLlCi4Lv9t1cdsj/5gf/aqhKXP72rBTevs/Ua2FykQFi/Eozlny
FkeCRdMEobPtaXXCAFk0nhctOHjG+6Syl3A9wMDrv+3N64AgPhVnoX6RnGcXPUaUOqYMWz+eKJ7H
tcPrDO2Ffh3/yFjXV44ymBicNM7o5rw1AGhHnvf+Lc7GGAAJSmKrpBFGnb3PhgLs3xPRtZw6aldA
LW3FvPYD+s+uq3Ux7ZkZLLf0LyLBDI9ETg6Bpr9DTfYmiTRFIYRaQ9Krf9h4/qJMk0SC4+i3cj7l
r0g/7jOg8Nzpx0k0RYHmhnQ1g4j5JHkjMDnufh8v/A4V6yIDyL3nllfNKN4jQ8lGxUdpneiTivwu
upolrw/P6WiP+6gz92Z1ClozabyC1bIZLcF9rEKgo27IT+AhPEOd5104a/BdiM4uDNNiGd5RCqFL
m56ncO6/950KFFx1IPJ3oGZNNO/2HGNsycVXzSjBHuUrw4ZnreViGbd4ec8L4sXMsRE2BWfH10wR
YeJpI3SyAbi5gH2NUCM2VmT3wqFTTu2D+zN2YVR7K6i7ZvvlcnsdpAvcNMIbP3qzCLzd5eR1Aqwo
qYtC3rxuqZl9cTDpuJLnCDuJfgiTOOC3l5IA/5wKQbNcdVo1E3QucnoRPfHaV/JobBk+SBdvjYWc
hVxEbvegFXBr7fz+dXc20Ux9P8eW14JohrlTicY8AzpwoC0aZYJHlPptHpT7j5jQGzGd5UdUrZSR
YV9sI8FR1oJLk2t4sKEd9dbsllaF7+8qart9hm0Q3MssGMLNVA6d/TmNTtUQZrTgZR1o2QcUuD2J
nBwsdwLzW8MBRQl78Syuv1lLsWg/kt/dhhe4wCKp7OJNn2xRIj/iwHv5fz54fSV6czPl7PgbYTJ9
N9bbArwn896OYOtsRVkPeIoBLJx4zgFUynXG/iRFNNPuKRoPvm40R/CF9YpxwciQIGq3aOPY3lVq
J3sBxmZhdERe9ACmPo+ynULBXAJNhYszMuxLo7RXe+AsF4/yjWEk963aNxr59aDdDoKJ9ZO8RO7i
3VXLeGn0rE7pxV0w8vrxfpqp6B6KqGCJIqbY7bck6l9cDAlRei1CRfcNUZipuYj3/lUApM3xyp7y
t8Ry8Qg6LojpWMKiUb9OxxHGUlnWl/pgF33vySy4ubRuyghS13HnK2xmf+acp8p2KdAv6mAiMyNw
+/DxwV95KSSl5f9HUbi1ZJCKezjhBjQ28DA2W/n3DtWVVzue28dZWQqKHbJnTKQ+UbfoUMg9dWCV
zGzp/fg9b1aVdynE5erW5IMx/wJDBmcEHe0DVZAWCxz9rNqgZn/QoJMzOAsNH6k7CkXGPqA2/k7T
/JBKJxamjq82t2R9JModbdLmUIdmxSAz4yQA6if5wtInWVGajtLdKUCP7YSN1N6k+ZlI/p8nL2um
fqVDOzfzW9iEjqntuCubpoBXxYRWl95d/mJY3FWuoGhQrgblhNaC82Ocg5HrHLp6TBWDQEwvYJy/
wM/7nJCoSPwGeuF3gvcWvzfXLGP0W6Pk0ORgvyNGkh+dIxCJfP2uWphgpU3D5Aqm3KsQ89UPDkJZ
Ih0vaypzL97chGkW506uILU75lrMPg7vaVXcEGz0dyel00kkC2ee7pf9U4HbfqL5l/LsXqP1Vps7
HkAnSpnGxjAHR8oiwUUgpe1pwTLF1uZL24mx7x9vMS8UukUs6VtH8WjV4rOdJEFHBOeqznfm+lDM
NqqcF9yy1YPG+E1ZsMbj5XLsHd4cw0eA1mEG7pSSo2LnHckIWrRH3T3165JgzqacDpgtT1X1tVfi
Wn/d+56HWnS9jLpAGTOhjsfHodpVIo8YXzy4MBO0oHnLkHcFU6PC/lsGwEz12sEY8z8TKUMzKOi8
oCE8HcHjU9KKsxffiGe6oUNrGu3E7uLcwXZ3kMAbf9hKcKDmPVj5GwdLwPMHU4KfhXwupPHRfdzU
LYbI4s1Bq5YN40zYHrAXljfyf6YBn4wvRX7QJuTdiM3NyQkr2j+ZLYRPbqnUgeuVWmiaYlEioVbV
6gjqOTKNo00Ovw/aOrgHYthyBl8oCALq2YCzfZdCuxpU/UAQpSafteUPfEnhqLYnh+fCZd+dNQTP
U+d/jEbjkvyK1pu9Aps/dQqwJihtPG+qgmfSnpGdigftn0lseAAdyQzZH+DlnbY8NRkuCFdMJ11e
5MGe6BWyBPaoftofXpxUeXTQcI8ksNzJwJgYOcLoTmt2NONOMk6vXR9zWiCyI8Edp3mq4OGm3ub3
Gaj9zRjG7tPGGy4uTdq3I35SqEmpMAdPMxookSidEy/O9qK9QeNAGOthTHnWvZTDJEEanrqxdYwA
w2irM3y0UNoeQqrLrKDrmJU0NwNsCC5MwyfbU4P1G8PmptiTgAQG7WVL3InUl6Z2uuooLfWO9ZfH
r+EmDax2+y16sGzTqcNyXlmNDoNaoXf9qdVaMtMTbf7gTKuLFtqGusVlHJ8eMx/EWTZr4r6M+BNV
Pep538PEtff66B1bdCAGkOfAIBLyhN7iwGAk+61cuxJXtDKCcNx+2vgDCyG0dnclfU1ABBE+IAWe
QIUdwQ1tYPlc5hAODlvGZCi6Xf4qFN06O2LJ83zcfA9u1TxnuZJ0+4ioH75ENz0pBFIiOAizxVEm
QAe31liXrQJYxh0cZETHmynL26OyctwmnJLtOCJJ0A5HEOBea3UxhD9kk42Veb4z31VHHkGeDCST
7HJkZ8zyhhm7mN2wA65XZ1u4vmVTmCoa4JKcpXCJMNjrz6GU4dM4BkFTLTJkEEIOdZLuOw2E/pSd
n01SpCXjRESkngaxGedOe10O9tOqWkbpYkncgSOwJpfZ4I60rfK1LwnYWuhrMJs6ex07JZru+lK1
r/bnoULcyjLBuzoAcLQwa1CmZ4mXeQ+EHxitug9Ohe2y9KXC02REW26HcHHToJdSqucv1L8YI/bz
PhTn8kl60Sf9vSsItMogd/PjCgwWGcC3a5ILXKQImgeOT27r5qiKrcByX/KJn/ou3//Za6rm3iXr
4qgVLZE8mI3K9GoQM6aGodfBE4PHmCXJw/Feo0JcI8QE8B8Co58s+mWjlnnOnCyBW7bUZfIWzA15
cMUadPZ4b2y/YSIsMlAMwuxnzSzz/o+WJRofL+xUP0mcqArKvWVCpTzDTYRgFf3+Fv52j3dSg7jd
lHkNKrOBIXUQNxY+WWgyzTzfH+NcEL7XI2VK7x0eK+olHkE6YWv9lTf9T3LgM/2T6aD8kt6W1N9h
1F65Xgw9HuxbteGa2RKHIoqWTxpMy9UuqFHYuB+Y+gyfwGfmSGrynsnQI8DZAwKqw4WWt604Yftm
H6ONsyVkxn7D8IurpEEr+StjIHOrg3itRhv+BBye+Uj5ycQ3Yx4AjbHHcbbfIIXfnLVNtDfUQHUV
wtyupIUaRfpdQMUAywjtglEl9B5KAz3DjVnpo8X7mysJAQ4QajXFoE8Pcm1JDsg2jUUGeixl3Oqi
qBtkCILlG6h6bGkLYm0EUkYDTM0vhQEuR9aookHj7fKhFRnlJGX8Ii7LEhtQJPng4IYPSVmRZTk7
DrdLAFzCCHtznlK6hA2/f1JHZhtsiO0RBsZOiN8u95Mp1qaacF7MbNv2NftdNJApTMzCdRD+PYEt
xt5l7o+D4EPsba2JMwR13Odjl2r68q5acyXzQJ9W3ga5lEXAIThQ+Af59CWElBsG4VImOkwn12tQ
IuzgA/1QfpZX40oJUGfXIeZZCzAmDaaSffRPQscKXyJ8isZkwKHNSe4vOjtkGOjFh+PYctUMK3+o
0swqXb3mdLZCOeXM4UsCsKw4eXRvP2HONCE+h7NB7fUj850T1pVlk9I2MgPwMaSCppLVmWIfBjT6
AymSkasBArffx7byylkU1GiMMKMrSi7UveChBZ0TOe/xZck0uavA3Bn8nY0zjOIVDgw/yHELbw/A
BikJ443xPYFMHsGF6GTYJAwWBOCF4vb//rXmlB3HKLjXw2H+cctBu++AA3Rs5dxf7FV48wvSKVml
9FSvV8/3+KbYjXrals3Aw/KSTe4Ob2RWXEZzipXVpxngN+CrfOtYnsKausGjEi74U39SEkAPreoe
QivnNRNuLDHqRXkqQvhCN2SHaJHr5Rc5dSU7xllZORAuX8LUp/C1UcmZEv/hvfi+u2qMmM2yfpQ3
eLZ1iaaQnK6OT3YGKxlBub52QZHHjxNAZBQV+ULIQR0A45sgTLTqdmfQj5IUC7UNx73T3sJqHb42
nf15VgYpN7sPFZso4K/kBsPoRiDVXYzhZsuz6dRCMfGVYGliL5YKvCvBE13KWJAuoVQtZNi4Y7/4
uecaZMvijQ81K0TL1aFpNQuN+U7n5zMIjEVgYKCSx+MP4vTkxGY8EkHs1bQzcFeDAinqUtHSLUh4
jVIYlqj2kLCPe4dXfEf/6dHBPetrNVB2l9I3l7kbd0hKssNiKt0q0T4qYF1czZQWqm9RGu0loHEJ
y8ygypXhy9YJLZgQxLM7Tgvc8PhCJpyydNd7QDsplI29jUIkSHGCrmMJ0gM7UvnH4t0k5kQzleih
qbWGOGDy1sFmkYn16/GeCQQePiRf3i1gZC/P11vzimfThhJFk3Im4zb0fkngFYm8lUheZwPhqMiL
jB8XBbSJyKxXDhFSF/XLd58zakIuqQT/eSRw2/I+l2NhJOl916i08Af7MWPj6l9J1WQCHtxe7SvB
a0Pi6P4saBSCKrjpop7i013h/fyh9efIQTZ912LC3SN/BBIilGK0UVILPCInI3J5n5RusCHHaead
AWja8SpWt/j+I4UMP3kcHW1TFDXmAuV1j2PNr95GESUo3bj7M0dTE81+sHJphfvjNzrNxfReG3Mm
hMJC2GuL+kdORGt2dYs0B2XRRFU9z6VYus3mrU5/O3hAOcJYppXlHjfNd6c8XJD5ONqRYhhJazCp
bxfQsu4nEHH9WNxBFhJ9QJ14aiYYFUbaVfU0iKLL4yZ3cBqkC5oxRuc4W7zCXEXNX6biqrIkb86w
P2GUbZZ2ZZcTycyabY0PEKgR87uKDTA0H7oYWkZjwwA/0WiTOSXLI7gSTJa2aUOlMiRk3QDsqhNR
fD15HB3rUUItx7i8VlwzBiOdWNv9Yr1KWX0+yBEvGm0ivKi6Mfh8S/F3XKm6KMVDkSbu7bo0jF8W
NYopreiCFtAwG0WYrcUcQedmcGkVgFnN4yNc9c/ovPB1c23I/1eFt3ZT7SlR9hatlKyRSbFUg5L2
nm+tUa5PsbziVsDgdZsIkAPEjOGdxJo5JQ+yjhx38r/AbR35zwGx+nkQDHjZ3sPpRjm3DliA9gOF
xjkl01wc5JH4FBw25hRilCO2zw5je7RDaTnbCCjdJRix3M0si4FtPyQIeu2wdmYZ3oipU4l4iAt9
shDczSFu8ScHfsJZzvtNcu3W5E3t2RwNp1HY2FomVc3xtNyFxB0yA6M0M7pEjlNCgxTraHZHWX4Z
ddz3P7k/QeCyWPy06rsI2UnzaH9eXObtIWDUTVqJXYYH/wgzW9d+UmxVM9ZP/HtIBx2idFAixsG5
sSjqHN8pBzwCqXCxOwK5lVdxZYUIYmZG1ytFVDPrFRUhdjFcGXQNjoa/M7iunR2JM+L1f1sPaGJA
+20JsipR1f7dhDduurUvpAhQ+ZCaEjj4iKInzVOuNIzB7fLPVlGhQuv7LoIg+LNdbIKQVFZjBJlu
wMAODUy1BovmboX2iWZXRQF4b1RorSUg+nSLnKRs3kEgj28spsZu+Vr/8JnGCwh8C5vNTEVwVh0l
DuyZs9rDv2L53wp8ULKgnWHPrSbBFDoaOXw+cL9OERQf5n4wnUImHaYcodAVyb+I8l3YMxyFb5BT
3eG9SIKezRZZJ++/nki2Z2HXivwK9c2zcq/MT0WcVApGEKHChanfsyUyX7Rw4/eWDeRvjeQP+dA6
sWqIr55zxXw1IqGATLQbKgC+e5Mhmc7bi3ZduTOi7Hihd+ZNqCJhvSITBufJn9GCblNq63uBObfa
LUR8OAvRJHAGQdYvhelBhFArp65H36YDSd1TfkZbwI4g6gO4O4ltJXSvYJm4uOMIFMuBlkTb4fc8
LOPmKBTr1rzjD5qmHZYdzkKZFeagDalzx0nAQKHThIlOnMzu8bO6aMj0OYXpBfo+ectQhi+HpSIW
Kavd9Q9YPmK96foI0UgEzCUGyO6Y9VjXeN4QkhTbDKjXeW/4IbhHpz92UmlcujUBpZ8c04Ixbwg/
x2b31FddoW4TtmeVPU3YAFPnacJ4SjTD1mwb9/TGW6rPr3r68sgtj9xSPm8Zj4j9KSTTaQKOTi0o
spMkIQx3gkIppYDkBCxf1ck0rWDU/BDsGX76og+yFTEE8qlN/3SyD7Q/U1Mn5qI0XrcqnJLmxW+Q
wAcasUaxdggipxontv4/RBnM6P7WVaebq4pt9POej6R1ybTOhkZ4fDx0IqQdOi4n8RMzSWNlSmPO
fo6gGCSQHK6pOPAYF0whFjEIFinUe4DIlDKHGIh/7xSCdZ7PWCBovo9GuD4nfkaepahPZ1wD7p5i
9lq58P9hYb7e5rYLF6vS/Qbvb9csAm57vQ7rm+O5qTSieXC6Jy7Xd/FbBOhz0YIoINsdRihu74EZ
RQosxctEfzVeGKGq77fY/IKlEzga6PSsexZIWOD26NdSZka+sWg5TqeOjDG1AZ3mfcoriL0pjgsu
cSmyNaWWXx7+lTZ9JTyCT/Isn95vsWzC8rMNeePF12xHvbuLO7pwP5OOOtrJc9VraCPs0BC5L991
uXBajR/ViTlkUJDKa+1lA72x75OADDBVy7b9LNv+VCHENpkXM1AoFFTAISwFj2RriQsCzf7MrxFH
QH1UCfQVsxJozluLnexF2vnlCldocn6BOJ7IRDGmrnmT7MtOYzhfUYwCR4uQZZnH/3NJKB28GnRC
xaOQWdaHAf0goIdgGMnCT6iXmbPPLug4pj2yt8RdbtdojCEClMHKwBnoyAW0WnwoNZU57/9UbHbq
8AKKWxDTZ1cMQcdYqnV8yI4SOsHw57cCrJcjRHtmdSky26IKlvX5Bbbns6Rn9lFjUWhhBbhneNwI
+oknpMOhpp88AvopC5RH7MnpwnQd7IDOBzrVrbI0Q99Pq3Aa0h/fb/tRi8/kJcpcBRJgmHKYlefw
1r6wJOoXQ3wkppHVFuT1s/WHx5J2O8ZxUiVjPJsiIz/AZKlUxF9IKrQiyg/8PCwNsznqYXU3ZW59
+fh1JGKkCNTHotcX0Ishv4aivh3wrsQbBg++7VuPo6qSQAxxCEL7fVpn1gaEQbqnu/o2n0VJ/x/D
BxkW/dYcVRjaSuhMGqkAmJYi8fMUj/Q3eMbhZSmdr9KfykBZWhQBZU0felhem/BWMjRVauLzGIkP
0Taj97db5Y5AoGOaKh8vhcY2CLm8tohcj+062jw9lR/rlL+gJ1dytXAFEylE6pOCNzAoWhcnZX8C
y6mOferrcJz7wDtofENGOCBubLEDx25ylqCQG+CAN6pR5eEi4pAwIt8VIfhvpAbJDYbuDqSTFLfi
tSqX98EPHgkZvdxXsiGYfHBGrBT0lLkVEAX01rCBz5tz3cw8vndwsmxwh4FMRuiNGUUNjzJ79Lsi
zy09Cff2Oj/9Nvv8xHSZ3KnebFdxbHAHtQVbuJYzww0GKwvA1y37zYeSXSYe0m5QRAvJtJNTCtZQ
pjfkhFQmRGx+mmfgzufmTSj64JYChT7h6aaP5EjmlFyesMVdp9zhdQou2Di9b9qckAl4i0w/ds1d
QhXUlxkQCk/krEFeABpLa0pePaFVqupVvJsK+7Qgp9nzfOinIpoQRg+S4OBZtw9JGdzO5IB3IAZ8
V1is8jianrRMjRls7fco0ZfDOZeNhgh9xiHnOX1M4xVe+sLcoXWHIup6oFqnRbonG9QlQY8gU2O7
MIPeeGEvE0vZ57F9Hh9AMAfj2wlFZGgLGDOu1XXgDTF+V0uBxBi+Rp+Y7KItSb6hCQMp253XPgbd
hUpdCLNyBwQkLaefwoPfiNNeTcmq9wjH3Shxk2n70fOECLhs6NutQARw7agKRa2T+G4XrKr5UPI9
jrw81cDfP+m4FC6kX2F00Bi/6x/DRT0GE4PNk+VZh3LeGRw63xMQLSAl2ktmiwNYPoSgnJTBpWFx
g28XTWotSQPOwxslxvKBSE7Pbccm1idv0G+3j5y4VkWU55bTIMBdJLMgsEzYCuRkktM8TPXmbHdQ
ebvrggu4RsTChdVjxxAHr+Ibt2exdlqIsZ7JT5knrXLEWtB3LCtB+8mLqdujSejBXh1u5O26City
xPkxdEvx1hlKyU/qDIw7+WgmfOY0kBSYY0CfZdUBLNjCD3CN5P//3E2cson58U0M2LQ1Z5wgLTR1
dLZllEM6FR8alcrLLRs/rB5thJ7PKrXxsAJH1LxzgrJsb4ndhF6vTC0sv5+7m3YrblSoC/jWgm0v
20j2ye7l+c2uioW3mDzQPnDuMYynicFDdZYJISd+GtIBcgI3nPjBsI3yzqGNJhiNur7vI+N857y0
S8SHdUqC45jU3s3ssSy67m1qcYn7Z03u7wOaVRQtRXIEalX+LL9OlLUTgbeR//rI+CUkGq3+sYNb
zP2UZ1++XUzBlyiHu+X7hadeMKex7Yq7Op4Z787LdlLMc4OZG8iI8crMjY58YiT/tP2TWvmopxvr
Iyj4u+eDu98G0qRmBJCco4e+Ts12xOpCDBi3BKRCFfG3t1z2kmEwcyF5t3i50wf5WqT/Y416vZld
Yq6WcTv6uRb0ElgMcJiUNfTDXPcsVIiY8quIqUoqQqpVMXuw0PwkOsS0C5K16toAn8CIN3/20e20
SJ5ZsLUvqbOmAncPFgRvSQp0lBc5OrRd9mX/YKFfwUe1uIPPtGY4aHMh1qg6SFz8zoccft15idEH
uIq7aNaFwtPuXtFpH/ocVO33+57P7pQyUMzls/hJsPWGE6aqEsIC3NVD5J3gzorKJ/iNlJ33TOJX
qReR7OGQkOpySpHjgKMAQheJ7Ej9TPDhw/vFqNboGnBoxbg7J55vfg+GkVb2PYZcJgL6jQ8qUfTp
DlHWZYAROAf38xHQfF1NLjzcRoBtKTRUzPgvxTqaAHxEeNv9xFJ9Yg4f4rn9QbokX5AH7b8aD7ZX
FKHlZa7NPew0si1vsFtJp70ffWHr49VtFvzSkCA2sSL+qbL9l3GKgBdmIxp1l9yZJSOYNxpoJneU
G89u8yuK1VmvQApOw897hWi5aCsyTDL343iRLBcP1pU/YwrAQQ9JS00M79+9BCakY0dvePXmLWyQ
8hZVipw/ZNEj89FZViRa5mw8cDjb93AN1lyxGtpvtbZB6Ukiu39ogDdz7eU19Pus+mAvqmPxGjh8
hjLba0sDD1nrat7mRnBU8wTmUEeYDzwOM12KEuhc/nCMBt6Jlb8tMEWftVIBuQr+RSqyplFpsxHL
wVQSKyyz4Cir+ZlhYNbSTTPAt9IOtnbakKEbHRAeBDHueZO+v4KAfkYZ+ZJvx6xDeqq8V6AiUBfJ
t1LbQFJ8bz6veMxYbN2HJ0rK/erE9Ftv6SZt72x5N+dmMJ2EzKi0K/kdxmifmPDR8S3ewBXfoquU
k4+fM/EhmIuZx2BmEp9rfece4qYRk332vWZY3SPpdSl9DPVz2g2TbJAZevkox4mHC6CoUN6Is05l
Al3t+WD/B3zqYdgWQM64qboDBeklG8uRFbOgnPA3Kgq9sz2PonAPpK9g1X27EKF0WXvKGTQT2ICb
oBdZX/3oDwAfP64dRxmSbSh22qsX5KLnlERehDFOWzid5Ip4qzQ1+FF5VbIJrxwSucVDSw4SizYi
KDLWVAcpm5CYbojZPGf1BS507CBjrltQk0er2niALTOvzNIsq3sajxTUehDIJbZLtNFrN9uyCk5w
Jn+uSDyVXuTQu67llj+KCMrHr52YsFjnH/gCy7dQ6m18jHKeE3QI1nqAngJ14bGLpqM3mO1Grh77
6jYZbvhiI6X2JeaNIUf2VjeXa0LLc5NnBPBE7KSK3D8jmEBioO0cjFcqTXwcLkndAdrA7C6/4fCO
XEhMVbqIxxw8uvkr29kHQLJn9XSzGXsZ0Noq75FmVBay1sliv44kiUFxOP34WkdAcfVa8IF4t4tN
IJCoATwAKArefCj1xeopu5Tslpu4DRq4psbJGPAZn6MSeThcJI3ejJOCIhb5HiOVRNect0kVcntK
0medeejS1PgkZ3K8olpTmojpOriA/NKMTo+swRdp9V5C5i5YhRlIlbrijT5uP412+Pjf4JmGquzX
hk/NzHcoESQKn8+rJeU4ZKCKSNQyT3UFELeECBzWO+t3j5zxUrJmrcjeRQWQgv/20caXje0vPHyC
mUyPiYLzX8A8CS9sQCWioWos9o8Ty+NGlNGjrgjXkqabIQPT9VCiQFSyl4rcFNYMayWlEcQG+Eqx
UcZbtNfAfOZlbWTUOarF95vt2G1IwevrLeYn5xH7enIL+cz7MKVibpy6UXEZ0xRfy73DoF+vQLnh
Xy22b1F/dSNC1+TRgz97pNsY2d1cqE9k94cK4m8sUKxqC2n3HbnFLY3L3/3/9zJSDpPXkoYUdbsU
MWRSwGlcqgECH83rDbpcxrGr3fm7AQ6qZnjzz1V1X7AxUdcvCSHuV88Br2LaoeG98JxGpivTN4pM
04QDLG7HUL8gdYwtTP/X5C4ax41s3zqZhTVFDPqoKXSLaLWMzTUk5AYdp1aHy2t25Jl9QAERfeEc
pHR9MsqifrPm8GSZuqJTOFpmMaR3X9NxOnKiXHJ5tc6fCE2ckoLiP0vPLSnlqZAWQMyVKJnGSZ6n
3AlTkIR8PsNqIY9s8zSHQyWOahHgSbmir1BXBbQ2CBrtEcpMAEGh2IFXOuKGV8sEtgyTwWJ5g9Vp
7BdJlMBi3flCtPXem7inLWCzPWHEekNbUu9Cynh4q9TOOpOMRRmy/QtkovcKFrWVH2D8bkHYvixe
pTRb5VN/fwusLMsiRj3qsRY5URTbZLrwo6z0YZ5TYPy/C+x7x+NFC0LKeyRO5dn2cAnbJxG7nWo7
oOoFD7MY8iqPK33oxl4NEHSLYv96RDk890hth/4Z5Ex6949GEy9xrqx0idhGbBJGkL080j+m3Zet
teYZf/doaz/2JzbNMB/umUdOUc+KziGExYVIYp9TzHPcqm0yH7mtSh4Fzhb5+pkyjM8pSFz7YeRf
jT3NVB3PTwPILVGa2joUINdM9aktXqoloffg/g/E2LuSxNOQZHw06bF2vZdjCQBh+vy2+Lfk3CEv
PkEk/osnyo2CMvLRZELETYq1rU/A0NUUe5fhGfS+A+Cb8m1kQNRBG1KhGO0taS3K+wBM/WpTdcfN
hGXoB8zYVCL4Ixa+wxxstGAnicY0NK/er+D1xZvq+25NUyTRdkFikT9INwtoaJzIO8EF63BQWjIL
3AH+RHNkM5dn0+PkFJUWy14koVjq+LoacRO+6ATAv92XrvL4AESKyb6c/j0dqS2gB+k7+5fe/6HG
705HplGO0IrjhArQNwAPJIqLPIHbgdfgtC5KnlGzDuq92fGxsFDBEZH3AI/sAwDzDlWyyF1jEpGm
k4ehdVXW0NAJNEPcUlmbB4K/i3JCc68P08XEPUMXOouV0ogGETD3e1VzXVVyB21j/o7Kl7PoDyPT
nUPVUUF3A+SfizVw+9M6aoSVBovFpWApFj4X+18ng62RaCz/CnhuCk0Az8gZSv2vwZImXPMU9UfD
FCHUM0Q/rQJ2d5O2zBLTKRA85DX+gPAM5d647lUeVErmXMFIWmQXSZV40h0pJLCo1d/KCH7MtOnK
Wfz9ZdrPMoARfaWL6TelO32i0j+jA99EdfOhHeoeYhz3ujHvVRV6bdw569lzd/rKboLHHDLgn+SA
ZqF2n8Qp+0a5UsaDIAKbJmI9QLE2j90epSdQFghXpOHzQyj9n06wHENwp4JGbP7JjpiOyfV0ZDaw
bFuN+7MdNed/yH3lGo3DFQPamQnLNxzm/rNPwjmUM/rEG/SnWEcKJx5fMh13zlEc+cUoKI4y7Hk8
12r/hQRnXt3Bz0pGAG6vxUpduB5qam1F/oI8yQTX9gC/gCTjGryKotj5jkZ5fB2D4nnSQj1L26Wg
SU7NjWaLfSwIJ/TnY/kr8tyWb2bunT+O1cLvTJN9/Vg30clvUwtBCV3+vw8kypbIDlyN1C3HfYvq
Pn+8uL9/mZuEW9+eZ/50tJYy2MUqJjovbxTzyBglle6uSkDDDQgRU5zyy0u1cRjejd94vYiqld/C
RgdHx1l+nN/9nAmMlvS6tG4AECx6hxmNjGgD3Axq0NqSSH+m2egtyyOyQld8w9qrjKc+o8ME6BfO
5DyuGsPmkZj9W4lY1E1pcDZRWosu++ZbdfBZAMuXIqNabhLtH0mYCQhgDdts2iXi+c0QHY+3ypXN
x7J4VzB0uKLPK7saeIP1vBpB+oLDgBu5W7PILdXczXcBLQPEw0u+EDdDN27yZIK5glz5GoYnSPng
e+4OzbEFi8vUFsZTZatsaqd06sAamb2i4A7HnY3Ohn85LE6OCxTIZVsZ4SlyV61rwbhVmuL7Trgv
7suOh/vr1YJuRlrdLQMpxunl4tPlEmnRcn3pJ+M3RFGkyNTJw0JK4VNN2PcKBzXJH1OjJ00BpmST
NTXyCZdk2/RA0Xr0/GlI39/DRyZLHpirKCsA/4XL+9jaEeDg9bw5AW0L+eOjTu1PUgmG/nvHHBxk
RTT+vQ4rTnofds/iQz3JZFL8hNpYVVcHA1ujTdUZOV4fSYLteejsby7D6y3rdt7OoBQQ+ED3HxMF
0+KiC6u/l1/cflQvWSYQEbtJV9Z49VWBFe+HFLYvgTXAtbIg1b5HJL1OPLCsVFwtqGsKMTWw5gM8
L8TiV0R79QACTTd5UzoC1lHaWhBM1grTb4dnf3Zc/AQc+KX+wYurjWsOR79CZnxlTU00OPwdwtJL
v3lBdNScNbuJDw6t413jwXQvV9yqcX+ilLy4jFZiqS5OYcPiaN8mNdVUwMbslOck87EuXNqob/ps
x0k9gbTFOQIr3ceWaTS1ldjbf/aKJQnZimDesAQdSiwxpK7wQnzUuXFgB4vrgt350AsLG1j1B7tf
hc/g7GBoD5S3zWGKB/kUzrl6cHE9Wv3b7SgTKt1OoHTXlMqzBffQ/Y96rPICvvx3HKoSzvlpopO/
oVGlUh9L0dcVYDtECrn31F8HjkiWXkDn4zMmpLMgycofgaMZHNYMDvvw745LOgp55k/RlFqkyTlD
xX/NKBhiPYk3bD2ssxvhuqYCisaWnT/9KpmtDDuwGEr1VGLovpIvUV3g2yvyqdEsT/niAmpnON+1
gAC+qj5iiAtIQCcdZwghf4jUpkPmCh4Wm+gzc3L3UnCaCctAW9o9BVyfB0thmExWzxD4zEJ6lyks
CKwHrp4xfxWck5T7tsZIPRGiCNmZ01pGbyMsoexO5wF+hZkl6VnJYNtN3nSyEA4YDlj/ILYmiBHn
qgplRDrFWJwzdCnApMwfiMp5zu3/9XyMNfm11hHEW+VvuxlpkdXnusQOL52xVfaj/x8Qfx5fDyw9
mDK8dVl2hBh1vAc3JXiI3d1f1yJKbu+XjOukuTTopawiuareYqOUYKzqKdEOTW9csay6SXVtMyDy
lRBVL1ZzfgFLvAnszBWybs5F/Dj4NTiSBFtLuDOFvUKHfU8PuWxk5BtY/CbSJBaHcYacwAdhmtwJ
c7Ow7Pwo6TZ64xVZktefbQDRJfXa4pGp7t3BV1INKiwTp2+x0H/tuPMNy0pym9VGTdOp/mY75/Mk
nnHGOGZ+ljnxrDL3uLkgYH1TLFpllJeqhGdznW/J0UIhJq5zDdR56xr3wAoH0n1yRxPLzIv0Cwjk
EnlqtFI0CgwUJAH/d59fy5irTjCpwQIyyDBk+g1hF+f/ZqSZBCI2IsW1DLuoFeU1Ybr4I/HQxtJ+
tPRC22OiyOJUHNSyn+ZzLNX0sUDvNbVIB6Uh0q1FRexJHtW7KfCy+r4ZLGUrDKIIcq2EPYx80nAE
XO3igTNxeooU6knSXYktup1Ugu9VpaDi6L87B17fLvQWRZdU+1DAhDCDgI7FkSW3FQStQ6Jkkk7K
O1cxxfEq9BTWqSVzEfa7lSSehmq/aYTcQIbGlrLf/bMEYnohJt3JWZdZf7mgjEac9FYqYmnhufIg
bqVQlk7rXsE7tQFsYZyAoaMPsSOECTnXBZ3BFOmnnHOFEVzj09h/ATRxKuFeKyE2+y0YJHs1QEEY
q4AvKt6eph69Gh3nEn5+w/Suu9f3QKSXFyFiSqn6p0ByTqabiw4HVJ6k7iOCHu2ti8zI3GSYq+tP
VGHloGNkl9UzPo00utnkpRN+BOYM9jvhCY84HkTBsfuLM56CjMdujJw5VddJF4/2t0Z5WBsHQr20
Fy0hn9OmZgZ1n3kj3mmSXATZlWqiLp5cQE3WLTQBwF1DuTLzzA/5Cigxai5h1Ei3MnwOOQRZBsK1
QjIsLhH4WMLJ9xheihNHTtM1OaWX52i6HwHNSwcL5TDFQdn/kvhGvU1SSIc9l9AZJ9eoaTodo5Ob
x7eo18fNQK/OhU0NVsvzEJmlFEHcFuLHzNDb5uv8uq9oZtfpM9OAS7lYtoo0DSO9LjTZopoKuLpn
VruPN4gyvIoRTEk49K7XyhkOpXXDpYzqYGLsTJyIsB1jCOaWoAACSbw4B+ijyNMq2k+M8dg9Bljk
OkIh3Ug6Gw+tb6Dda2X8C8+xftyaJbhF2wbaal6+NnGs7UJVezLWFy7LD6sqfxPf1nzFz9599TUs
9U8ClWyyfTnSlCV96zXWqYYSGLVt2U4LJcvCBZGIErJls2DAZ/i8qQ5mQIEbbXaL52n/NHwnDqgW
98Qr9h3akoUG7KLCa9SlM9LrrXSpW6eZqHLLU2J3leL7DhY52kOn5iL3EbjNL54n4ddVqko1S+vi
YwE0rd+6AYHWgLoRzTVtiLSjB3nvbx765OAlGHjqFQw+SY1a2cTEXMVqH1+xsXiWmJDsYrsX+afy
H2hBWV/ih2QEUrtS0L8FlAYJjtOpvDw0H2/ZXg5Zg+K7LF83j46W5eIK9+wL34CvyUKszcN7Nlnt
OfDuuybdXTutLwsMHFIcWiIbETO8E74nJCkI9IzdbhOPellX6ywkhF3Wr5aAqdhmRodGm19HqXGm
SucG2R/TQJ2OEhmb5AkVGEXOPkAlKz0GICnmt62vFLGC0ovZ6SxxgA5+K7Xi7A7hJGdgWsC4+ekU
2FRLVFoL9kpNqNM5bQSJqwwhJxhOZGI3ZCwLxkmDy0kjzbDYPmdqeEv0Tva80uqwIwBT7WhYnJ9A
CbNCUFdLKyJ6KUGQ4L6ug0L67yS2NmowDa2i5V111kv7pYdmt1mQtN8iNTHbn0uivV7y7ORg8Z41
ryma6uxV+ivrSK+QhC+iu7orfjhk7xczXHsf26WShj1x5O0DO7Tq2Ihc6Fgbpinivo/Q5HA67CJp
RUCzwcZT+w4crMb8wVvo4DJu1hXKNB3LeYGNG8xn4Epxd9R2g79d4J62YKQXJmZdLBIQquFBrxxn
09ta3mDhFHG6laB2urxlKYylHMJQ2/k25uZuwmBo0DQPEo1YseMFTSa7HWBx4ya3s1javzg/fHX/
gO7etuxVWtiT+wGdymJq8dr8tWuWqKILM+Dxrd2wPuy9EA1Ovolix+BZgrOKGM+xGre/YaIlhDvr
fWrbRsI8G8/sIKKxOpJIPBjQh1AFtcU4rBG3IlbpbcFzvBJvDj8c+7y0ISV62ryqNy0XetjXdTPw
eQZMN0FzMZC+pKF2GOuriZj9mLC5mH7PJiM9aF4AHn0khc1JWbumrqSC4TpzA7ZDrVedE/NFJjHp
I4NXNrglji/E9B+mzTDC4Xb/Kp76gOz/P9VOABUeWEdpeW9ApY+ieCW9UZROa0eFtqPWEWfl20fi
9lZYVRZjybbBE1tCVOna2BdGGpiYO1fHXJGOEXsafNMt8utnbwWkR1c4TjPcWNKMPzR/RUZg1TT8
Fk9V9FoKWsxiR0dnlopk97SH6KDYUqWbBw/2PoFzON+v4e3Tp/BwWgdpWtgNe8RFU2I0iTLkgIGi
vIjeDa8j4SMSpmVztP748+b8obJAgmDcq+LqBIWVsFN9B9qAJpBr+WxJu3BX3ck65TiUkG2ZEFKU
BnS8OpZtw8pIkZ9P+XaVouewgUm+ZSGzX3AvQ4IG0QcCxoPQax1QbeTZV7tcHweSdBOR7X1SEb5f
+biwmSQAlfm+DhpQWdHSIwctAQ6UzsR2KnBm3Lw9I7EsjGyjK4QNr7n5UrMa57WF/9h24a8HOuRG
u5ewaGyWFZHGa1L9u9XyQHYi48rrdmvLOTkMaA89Z7qpzjx67SF2B8h04IDkasSdXLkgpdO2jB6v
LHhbaW0frd6FrQfx/F3a8bgPk1NdFRPDkYUh3cjkgJqwU8qyJ51qmChreMsegZX+7gM4GxfiHF4M
GzqMCSpJwUFnnRe5VczcZoJb8kMLX9M4OFnZeDbadmBqeJ9Pdvx66jLqtZVk/F+KDjEXRCz2tc7i
KvQBaW6lnXadU74qUSLk4flh3qTfhxB37Tt3WcISfPG551YoFmEwOLwPeAKqQ2apRtC9NnG8Ec8i
rW7lhAvqtROmtolNntjO/Eu/YvcokNkLCR2IxSRdwvx0BsH4oy/VWfoppBBWRK+zRl5/Vosgel1/
BYwuofEjaaMMDQcxZXOdSJn7mfICRWSWLagG23kpTXKxSlIda0HgcQe7kO7gDSOsPFjTvzAJPZM2
2dTNSt1bCJmvNFlCBmfKyls8ECY+4N/u1wyZEfbukY2ZfEutzUERjpOHQxj7PIUhsVdMyxl7iMPl
PBMC2IkOpbQBSH39Hn1LASEXsVX0sKaboqkm6sJNYXuYsThvb2sRg4A5rgzph6rCzZaVvurwizxc
k+jrJG4XE83JLlZgeJdcsrjAe9ZcXyLkNRoUhUXc7MnUUs4TGJco2bdwJeMjkBvFYsN+TkxbMWb5
SMgukPLJnOGAaOm/ANKcitxczBOsO53jcY1YtvxqMwTRtkzmkktpayegEUsK+ker3E2/U4e6qVFD
YNuFDlAAWV8osTfGp669fuPogLda8pI+KtKx9/VwXBa0VMR6pY2mbLXBtqIkqq+KI2lN0YsV85TU
zf3/11nJZ2dmm9MvD9dnyVfAKjooM+tGgjMJsP7tUXNrpISVXKVAvsLP8+d8zdgSAesElEpUFhxu
ExirgKdZS2nSo2HnJIKDIorPWoHmy6wq5sCyw1xdMaij+gmmwHnJ8H/pGmqv1jfr9VYD/kIeL5LF
BwPhytqeidkhS0aCi3WzD8c7lFMQyeGwdftvegDWgmyIxx3m6OGkKn+IzMqqbM0wIeXikxT/hwSR
0HFPCn0dRUGr0lOH+Pg4+U46HKB8kgvqgcm96Tfj97vsjHi8mwjmIcmTnY1liDExzQO7k9xOlw6z
IBluU4XjdSyCic4Oj41ZHzKL19yHvOeyezLDcP40ReTLbB0rfYXEuJkk+BCl7BQUMdJlI7nNabR8
zwDBwlxhJGPXufVMLyy1CGZB5bWCMD7Ym6lHbupbiT42FogcsL/a3bTmgoKrTN8J3T4zorqgAcSG
1HH2vPz+dV+OfgDbG1weiWZXWk9A3/IPNMJrZTIlFsvJki6PfLyV5/GP/Lvtq8bf+2JyuvHZQmuv
CvKzTTZHO2fKQ6p5Swf0rHrZUNu0I/RX/8oEBGy7fRgvTzuPPtLmtRXAuHUs/8WgXSnK6XqLNsAI
GjckRivulRqNxLES1QgVfBbhZ1R1HKXHunU5/LNAr7kH6cNT5VzozhfQGlT+wtMsEjwYdnu9ZSyJ
HuSMRTk+EEI7q0sTd3GO06D/NrwHVfyJqjH5EzmR+Vr8ARvnXI77HsqP8jBGGYUOGHN5f+U84U+2
1kxbDBrn0bOowTr5hgBvfZVAjjj4PBQ6X78zx5+aACkEZsMxX+MqgwSImKgb5dGb8hGUTJNJN6ca
ea1vvUoQZZrF7iotsE8DsN72tZBg+tb/9BVFR1ir66i9oC9CpF6236G9MpQlqMrqUQI8Tc9u260V
NpL67hDD8Ee6fqk5dZID3at4LwB76FQylscQH9Gtlg5XL0Kdy4gACsSSeN7C7ti+0TC6Yx4fl4u9
zlzOnqPiSe3vofSjoyrqskCY56/XdfNHDkfsZ47OllsO0Wy4S3nOq0t37xj47cK6dsqD/S57XkV8
VdDIiytCtfIBfJcNMPb150QpZdxH0FcUY5x7exDX5aHBJAb8v0Wmqju19TnnAWKX
`pragma protect end_protected
