// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MRsgg2YBJDYvl2zgKQo6zZ/1TAkgISCJK3jx6XP/FdRptt2GNkOYJg/qz6NnHOMp
/t/knnrlUGtwvnLQWvd3ZGbx/RAdUv9+d9TCzN1SQw7O8COWHldRCxvL/VTlVOtG
+KrxyFRoTCHLLMDuincn1l9J9JO6/k6JBdgSs9VHjME=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13840)
ztT/1WtBrhvE54uyR+DT1YG26wbIOIYSIMeU548siL6SpB9dzZuJ+ghMcwPu2RQN
X7/wuurXT1aXX03X21F7+ZHwa2FEqjKFRKSqA9p/Zikyi8ZcqLEnuKeJrNgNf4vz
lrwS2vuIYMX6S7x+6t6apShGDQNY1iCJcMykDRW/nE637fzpcX6DjVZ2HSPJGJ27
q5zlfAYYjbTfAHiblQA8yr/Eno/JtnynXqJz2iWVkHRtnfaYXAwxxR3DVa1elHVJ
CqOltdzlTCPNl/nvJqzYWQCt95WMBlxCggHWR4ddeyQxm5XizqKPL6gaxCQDasdT
zXsyYPYmG/QGc67KSV41ETljUiPabTJJRU4HhiY4roI/tQvxzFp0SmPgKcKuFG+U
qpjsBANnFGY54mv8dmY3T/dtsYTOc+1MuJ3IGUaR9KSfAoyNLjPqH1VBNZjAyREB
4PTUreCiDKeA0L+hC58YUF8qx4yhxaWP9QxxSxJjOYhmkrQ1ln4WGDJafH+p7qnr
UY5l+MrWrUnqLPqbCNVAEvwWK4SpDBMcfZ5jWDUcOLRhSu4+igwSOHjSI49AB5ho
u06spD9FEni29rSEZkMnLH346Ew7q+sy7zMAb3UcmCWPuW+4LJ6T8atn7GMTbN3F
W/GMgkf5chNtcoxaxhFgTNVu9o5LIKvLaWXgIqBOTGV7n13XpMOzCUTCp7ThZWGh
d3D3N3Ij9gxlvtwkScJ1wfVA/q7k1Y2HNe1uViRJa2npxphR0kIqyDbHWWycdr+H
NSf9qRzLO+NmctUSYpKV5eC4kYG50Ct8eIjSTB+BRzllkgAmckaSdqfeIIYvA/NR
LMbPO7+wrNqvrEIREogm/Q5IfKugkWzkt0KzaK5BUi8VPNy0OmXFf+KJAUFDFQVp
2H2sM/kJUEUilOxAgPgczheNt6buJPDODl5qV6VEXcQkfRaeLO7wzUXb96iBh6zj
65GLkrkyvC+W4JhhU6PnqyVkPJ2uxQeIv41/aKqKDw5Du5YbK4ze2VkiTzUx4Wfa
pWxZqdIBpjqApLcx33X4wVWCyIZ4uu/+/pM2KdjM4IdiZCEX0CtGRoYDF3DJRc8B
sSv1YQCh/R5JyRmiBqv6y3Tqiy91Glpg1ivAazaPL2xEN9KwlSIvM06LFIJ0q0m9
JnP1NgqCj81jeQ/EIXfptUNY++WIlC0wkaa7uaqDxssf7GMVdm1DS8n/STEo4i1T
8OR6Agq28NTk+F3ZffdlI9Zgy+px5pOpjMy8qIhs5jmn6ZGc9BSTUlPWhYbmzfBm
klmuT9soCeFlx90gPS/wami5luDxwiZ7c4pUbQWFYNrl0sJZtvLIKb7O/AASa8fl
EX7/5Z5ObynBD4MZRGhRxKrhHHlH6uh1aKbulz6Czq9eLs1aQO3Az7sla3AHriW2
sdJdyhG3siH/yi/54R2xYLva72JtiUum8cSXpK0w8y++ScCbCwM3AUsH6RAql2Fx
xDydwaL2vAw2RhhXMsEzsiSNXxmJcjCbAGYw0tW0FsoME/UHRXLky5XM2bDsSl7m
Q3oWXO4Oi1tzlLXPzSOlotXpAeiGrgGUgFJlVCccZjVov24skdH7J8OZFALHUP+N
VV6e2yiN/2hxtDBWMWMAcNwTOdv4tBqpSfZ6wgGjRVDr0Zi6VH0kiQmWs3dB463H
4Nl0Xzf7iezN9bcgbTUHBZMIIt2+i5ZbIbpI/lwZNdJhse1O8OuTe9QOcKqLWh/u
ftMqzDTcaSLJ70kcNuzyhKx6tsw2Tb+mG7p0Vfq+a/WuhE//2fxuwdMMeVbdtC9R
wYQu8HEykhdxu87O1iBi/QGuxm3s7xNXH/2p7Ckj+bqr5kb7ZVXdjcVUDAOnev8/
4aiYX4e2v/eJP6lAI6czAIq+W43MFvd9asQhr+LKF8FNdSazeP6yvVmFVX5SwknW
cf7TqPIEA/QEUNN5qlYY8RA0WgWOgSdVZkJavFuDXWNVqkm+jBp/LTYeTEmiCSOn
+hjK64LnrqZGW+UeDfcqBsgUhdMiEpexnF0Peyjbre158UYMhuNfHOt9fYShudHv
mueh2wjj3m6K09WbY5z2BqKfhJThx6pZCwqY0RyFouh/nAkMUdkU2pwpnrGAQMpO
e0yrrIoqdJy7fZWvF8q2G+Ko6QKQb/8WlLClv0+esZsTVrp91OIyvvS7SvZnHTsf
79XI/pXJ42XG84C9VikWaSYuuJ15wyHTyYsTH+C4+edrn3apsXdvxfwVNghaKCRc
CYn+Vdb1+oTU1unDcIuZbCaOja9IPILqOk4LXFZeBR0ULHBvww/jASobvUymx3Cv
8h5XvYYwwlkikC5vbx4OfCXZg716CsWq2b/9RLZ3dcz86UJ5xNjm+bqLpCIKPgzL
CwiuPQzlvgwb4rSIIORkeae+HtNaciypQ3rx2hMPVjKTc/GTb997EjQ99uUmUJ0w
qzDUCP1k3MX1Zku+GzVWsgsGSmQc44RdKszBpNleP8LruO1iAt094SsF3KSnAZmL
DLMQ+wN0Sk1GB39wulxbTTBRendqpyv9kqEGhHjQgXypMa03xulr+dra+AmbjPgG
v70Mg7i4HldzNyeYOf7R5Xu2lKf9upmL3NxDLJ89HU+6Oz0gdippB+tAfTWILKyy
55QYeJkRVbfD5W5bHBrVHd5d1Dc7V4ziUd/kP6ImsIl2DNevQn8Q5MZzKC9S6jyZ
xyIZ8CVcamXUHpARSbKnQzeLxb0Gj9PuN7DiDkXG70HpStFyAqKAOLOLdaih5H66
zT+a+cWIIS/XjxiPsy8vPYDwMPPIrIHngoVImFCVkfMdjE50h4N1JW4Qo0mlqL7z
nQLqtuDaxlYPEXVlqYNENU/TpryJ6suOof/BEMB7p/yF73gS29mAndlqSkcaH1fo
eByhQtJPVa5ClQKrjzt9rA6/6xO1z1AYV8YmBWKPezdXHCfGa5+j626EBU/Kw6cW
sIFvdG2sB+8P3nAyruX67iUg+D2eterEPKgTb7WplSrSW8XEE2u0mwzzRh3rMOW3
qXHyuCuxqQsBKk8ybl+AeVFWLwOqVq/gPB9q62aeSRF7IaiYuP2oFReus/lmE6gB
wR5UlOrixPRK+B27xDv1/mjcbjyy1llaMZRG/47U2IrHYLRrM0+Y0ovlJz0ZesRS
uiQ+2SD3E81GMjAOA/oqYT41EtYkjIYzzn3hybWuyNwZthRIlkZ+4yPY+0qhqGqF
VxZV2TgnY1tIH9IoWZV4FBXtLmtzD+TAshKLcfCPXVxrP9SYLn8aosJTPK4S/L4T
azLyJnGSdCsBGA5/OpS1nkXDAAN0VjygiDRNv9Q5/FEz02mjvzxQJ9emELm+7ezT
RPD4oqpwpYzRYWbdLnhxodVsLvCBLqeTAuhOkr8WDJ/dl9RNPb4qJSnIbmF0bjyW
nXSCewbKMIGCd5zzHH2rC/94JWNy+FQXqhmRYP647RY90KYRaNH79sfrcIYwls9Q
F5JcO2iUonh7QJxiUWIPL6nlsTjZFbLz0wUma5jMtfPG8M6wsKeyeXMKSSrsTvRm
EehgVI2Pwzljcr7G5ho4VqTalnYt5t3pc4rCZn6Z3YqQT69djOtSAQ75y3IjjCAX
/UEEgWt3SUhrHoGenta5GDeheJUaT4TbCn6G1UoM9ZS3N3eMjtv09YsMcSvER7CE
LOhrdXS4N2iqe7nLqqdkhgcoV29Upuy8qWiyQERe56Seou1cg+/03T/q29gBiVil
HSrm4GGKPGFGHvZ5NFZQFnXAPck8IPEIHlpgTNndKuNiZR3x/bLMaW6Jb0iMeXfB
9V3c4N83bRUvh/7IEgmZczJHBPpaAqWWD10cPbmEHCPO3T/u+JiuIMTfO6f2WYxD
uxRlb67Wb+58Mv3Ti1T6EdRmPhE4U/CzDdBZz/ewF7j3JCaqgYW8YlkWPQsSBibH
yMOAzgGm1ECIy1dq2D9VGMa+zeT72sMq5F1+8HtLjNea1Ti1nJ/6VN88Ty88bv1M
i8GdJNG0ONtceVDHiY3G8fr9T37EgAh08VlU9W18bdswifPIcjTzQtio0JnEBB0J
X+lFvZVzScmYQBzgTFdHmZI2nzJeDp5X/lR+SFjuYsmOdFTAc+pUu7SLP7z5AFeb
98WPesWJPNnhhqeUAkleVMm+moRt5bVgRAjHixNUss+3yDHwaCwJqnFtMO0PgSJ+
qqT4rhxj9yNRbNyVuxOUckPBx8Y+5/RYiLdmWp18RQBaJTU9n7nshF/mJp+h4Siv
0Qp6gAbAaLEMS7WWLuKsCeY0m0rRxOjGJ0Hf/gZUkBv6DkJ3RuRMx34UYHe7XEkT
F+p05ERLtQA97zkmclVWn6X61k2JhcYyIw0yIUNFmIn4ifa35+L81wD4Exe60PWe
1AQAYi2NFUsIsdVaazfRdcxNIBu9zPceh3BgP6ZJ/4tKZnRcouC+bkoB4S+XFmrE
BNBYt5R1x9lda/CW+R3SqKmY36Lr8fGECC8s9MddKvBpDcSQZ0kPp070d7xfYKua
e21zwe90GLbMPebdd/+XIj8hhhxQXZR2wf+/wNo80sLEUlx63cEsU1mQwZiDbfZu
HlEhg3p6LUMZCEBo1Hhsj2Eelol459KiWMKaHGbiIHMoxAjO0WVVEyBv85KU9uIp
F8NrBjTyezKnOK61jJMN+0hv7/gndexKxEKu4a8kX9uN/39M5oCM1tiix8lijiTe
apZRO4V3YmdDw7nb+LeFpXpFTXylM66g/kFHBR9xT7k1XtuCORUQLsEJFf4Vk4Im
GcJ0x91EOY9BYSfhrmYYvZELcFCycCIXS27PTakCUAvQzrAT+IJsS58CzWokhpLy
gcXXaZ8Q2ENY7Uxa+AU8w327ij6O7kN9rcCeBhLTO++lL3jnzk1cxJG8GZvZpkPF
YhogPX3iE2cMOUwI4JSVF71bIU5Blx+mlQmQ2tOGQmL7fIJ6R/jawiu+979v/muy
lJU1AgYs+E3RhHqe4qIIFjFphB6EzWiMt/051CGKT84JWpHl0B/f6gs5HZjiqLCm
hXIy1sFddfTmSIDDiulE+gNL61dqLybHMhuPzjjpvkmYGp/J0Mx19kuA+78vxYiE
MNYcoXmr9N0p71B9hYNOhjCwxqRUTFIEqOKj4XTGaTjD+PEBXjxPLHOLigWANtTn
av0RTbeafJyJemSvuIxwHWmmCFMqQgfJmh5yQCKDImlQv8cumnFM+N/8+VJ3Owhj
oy+XuXhMRMOHZ/z+Gd246U8ei35byiTQNxt0GViD10pIjeDOgFpQlus2KdueHtEN
w4xccqfx+u+RqVf72RtZG/HMMUanXrftzQNAmhosY/dedfD3TXTfCBmLEaaPwOPY
zZjC3SXMOd+jCgVgbM2qoakbsE7VIr2yS7KmCaH99UmxWYHUoDK9Io+ZRyQOp0eB
4cvCpHIu0puVsEP9VPjE/VsmvUEdE3oyKq/ObQ5QZh9Gb42xM4jSMVmSmHIh5ofW
keRJhXjxxZswrhz6JphDlQjIe6I/inb0ekVzBLOWccVEi5LnHdOZr1yyPdcMx0cL
i25WKOKmURnSLZZ/ECdkj5l6i4ot3xukxlnDPyc8RCAY/g59LwzoGdER6EM65iOn
RSJx+gD2/7d3IVSWzzoMHENmskTLJkGS3xxCFERE8h4Ep7qbDX7KBBuw7iFd36W7
PJNB0OLj7ufyGFPfZHk34r5ftGD7rP8RpgxC25kqgECEc0dgwfkNmsLkYWUhLkGY
X6doTC93jCtjG19QX+sAQ23zpU158dOUy7D2VBhgbPwrEdFq7tEEPY7r0lUEoS2S
/4prIhp9wXBwgooA1Mt0LXNeEE+4ZaxbwsxCNN4HLwZWxS7TIW+SoXm158ZVPnoY
ZsCFn0qWCEi35Osry0hg869cAbWSXvD6ccMI87cSWgflb/q/jdJkd7bqavzIONZU
Z4GA47GtAvYjwWE8lJ84P0v72TPD3aRU0hgpeSYla1sKESmiE0emtDN2rNwVaT4W
b/vQspnGFJa4yawjT87ycKr8vp11Q6uBuQ1SFEHsorb2CySaR8DQF/b72wm1gcm0
EItEd0Hq7Vxjnm01HQ58EuwjKMssqmIlH3a/focRwKlf/bfZBwkhFbBMyKWwmczg
8jIAH8BvuwNk8OFaCvdtTGoR1aW/WWE1YjE8fr+MMXgmxS0d8JA0lqbGtQs9o2o0
cM09PX+9dMk+NK05v7cMvETSlNPKgW3x+ctxNZt2vxo/hX5si4eQGZh3FXlloe0J
1B3iDmvlpyHtO/+/kKB56ggEPxADsG8jlJToFNDeRXF0AGy7wc/U78CSOvbpxWQK
68ruxBfE7boVUxUkm4FACgrGFq5R3GV8rXt5kpOaBI5G/V3012rlDEFFtVKlZPNo
7yRFUBBANuaMIn6vRIsLuWF5ShYCRZwy41E77/abp8vJ+5OtQLFt8Ov0ifv0nBih
3gzSbT1iUlNfA7eP3vkaLn90UiKSO12sDrmiTXvN97P+oza43FchFSP1HC0BdxiJ
Mzz/QjlIue1ySxHf9/xfkm2HhHsL1oNkczG7zhAJxBbE/MqILgkEQFHtLPI5zu1g
un81q6T9AdrL6pcdtYl/T5e20kqE0VHYvm69wxRraeHzW/UzUvLVf2v6eaDqaK/y
yu1WCvYIkdzdzVpbHNEesJvlJgrs4OFN1k5oOgiEYgKPNYtmCTOWApBSt+6lI6Qb
2OpNtHRXBs3OtV16J4s46Y4DhjilhlMSrzFr5uJ5VxIAdgcbl8vL5P+s5b48LMd3
XWJz3GfgBnCi4NCyOEDdCAwfVWjTxuNRjTxnhptTVzxa6R1CCJMW4HVMCqITlOyS
iJ+0BIepFS4Rcj6xGYx334gNxQ9e2HC1kOtD8uOny2YPZ4R7roQcK8ptaHwqYq7E
r70u4c5QjZGDWUCVj3mBo7153STtl+5DYTAS/rqcRSaGEWooq9b8t5LNZODzfu3K
1xDFPcWQJOLjtGd3+vtFoi4yMSiBp+8aOJniID8W+PzzFEZPBrWUqFukwt7zhnoB
Er/ZBDc5fHhv1UFCtFIZuvM5VMbgW0R0nqkCTr1SrMcMtx7g4etFEItNeW6nvPUI
nMPa8S72TV4KE2w4g6m/auIKm5sLqxhEzpXbYODxfSSSDrFlsCvW5th6XUJNDoBw
YHY9mTT/DPh/Lm9ccATsjdDDpqWZbiqwIfdVfVdpcgNSe8NkilEcoLqRkJ0x7bo/
CJieyqkNNrmKyBtkHGckwrCsqcoAqI0oP2VgaHZcjU5w0gsGiHzSg1/UP7T0mgsZ
xQB7WI2td3Ot1JPQXTDHl89nYmK5hmS/QNCWbWOgBbKnlpalDo51AfRRYpt7rSEm
yJ+QjFSncSLkJrY1yxmBzozXm5TaM1r6534YgZq/2VXchLCcrkiYvHdU5VMD9IK+
Ut1RI9eoa1hT+K8SDmu5OzQqajfM9Ujw5mZO/OTXjCSuoWgu+PREsdlortuZRTiy
LMvFgzDxFKKFX0WlFmKGX4FY7Uz+zrTa7MdPQ+8eOYF5CoNghtXDKJ5FedLhnvCs
yRaaZJxiAgAymRFQvPHbNqF7+LAXqUufejn2YZ6RPlYWmh1fhN+3jZsRFEquUizC
BY7U0smGc2ErGVHFvtwMB1Tnqn6ygFdSIuJErmTy+CL0WAy4oELfROVN1r7Czb5G
p8XxF4SNFuIdQRbNwSQm5L1RylTt7eOcuuxX85EM/Z+jde6j1zk5LvSU1gWJnAus
pSpo7kwenvpcCuaGjxKSRmxScqx9+IiWfF0HugXRNbe22nmn1bNrg7mI4w6OkyOX
RJqcikQgho+Oy1YkEwELKZRklstm2iKsyEOpXw71I5WNyvPPCEJ20o/Ia0cvw0Fe
a9+K8Txu5ld+M/DnzcObJ7mN2pVD8mpJz5aDqvLbb7c1jwNiBFFCuWyIqFIf4dTS
mjjzbiZInaDAO42s4u5IzUY8lsesh4tzn/PgzgpQLZME5iooqDXKCaWsHcmD6Bm7
joXHo1CmKaLYNTHZO7bl3cLfvTC3/8btFYe+HMPgw3hpqVmdlK355FSlhdhFRiUD
8Enjlss4DxUgcpNE2Tn79oTesomjM9l4IvKHdL11WRdbqQo/z+9tcqFRouiH/Gvn
ZcZbB+1ZyzsXJqFiRhVlnx2GHfezUWAnGSNw2UbUAWbETM/QWx+R2vZ+TbATbZhE
5LDE8H7Qs7SJm6Z3Yf59lSYNYdMHmLBOnAPiKmTTtLe7zi40QIxosnu2YmGUS+Zk
BmUu25AiRlNZFYfPviLY1rkb32iovaW/7ubtqMhuSfgHZXvoxLk2BA78C1HqKiDb
LyE14hzQ0oGV8iU2PWs/rBMe5YuEYW1eMEpHBdBY7LPH6mH33xbQClhC0e5qkvLI
JkIXw+zbIFGcOWXQ+qqIec3zECZQV5LJpYb0L+VWDQXm1YZN6aVBL+vfiPEy61lc
HRqXDJpBqjYJ1axiVMEp+Q+GwN7Ah/DhJFeB0F+VlypZRw/Bx/gJk0XhOtLW24EV
sNifmt49+XUhHOSalRPuMw69Faa4cu0qMQGVtzd0PZJ9l6gZWHftqE97q7iKagud
m1w4cPIO9YLTshW/34LQwg+WbcN28nGLxwkL94vg+ESGNuOiKkj6+DYWccengn57
g7JzkXO0/W8oCyR331cO86bfoxqnjG35xoY9J4dANcANhQoIix5y2kTEDC6cOUV/
+qvPoyTb5VI5p8+Ysm51Hrj3UsDEEJyGh12MS+kcUAoKv2uQLPEmirNHujt0c6Ye
a3jduoMZ7uHaXLLUtmyOklvIrrIAyiE2t15dppf1GsCp8T06uNTYe5Z0vZ7Zra3o
CFyZkEM474vGpy7hKnmDvV2ulfJh+bvYbPAlbu9b/JCJwqn+36A6N+QeJVHgX+n+
UL9iFamHAZo4INpqVlfAU8YhXNj8V76pUnBATiLDvTYDWtw8uqeOlvJbvu9bvyvb
yy1H9wIKI/pzV2H50Xs1CTrmijRmFTJI0iddE47UC/A1R57iVZyQDNNY1R4KZbvM
aKLG4C7BbkD1diivE8QQOFIgpC+ghS8Uqyka6Dz/jUHL1O1Xmoh0pYMD3sMYN74/
WKMFf0QsS+zfcFcY4m3u2pItWDIxtwDeceEVjZ8UMAw2lxGQu9LyuLmRJ2mw8t58
inYJgbygl9ft1gsScmsNmYjK1LbNzS/QUIDfbXdeVcaAws/96kY+pOlOjU02EvYz
2qwbtqRiBfauwkRYeTDhPqPzTMyXkqENnN5ie9QdegkX48Zg7Dw8SttOsmYVT7tf
fp/GDpmOPLNOpvi/rM9bf8p/KMRL+DA6X9qxBcYX9r+wYVZ88qCzhvAygC+76mNa
3Spr6o6GwnHnWhsjnLjn1AInkt727qnNmNlHXlRv2YDj6Fk/Bax4NdDbT3juR5Vr
phFzcTlTlDT2l3wpEPW3iDiyVoVuXr61HoMXawxzQ8WI51HtAL0RMW4aSD1vEGq+
UECJSmAEVbM8IL5td9EtYzx0nkje592Waa91yYJERVxm8gojAkqQIblAOAfCmOwN
fzEt37qoCPG5qHxiAIe0B9+G5VN4S/yFuzXJyB3umnWD81x+UbjQS+n1VCHIIxdX
+Uu2uBe8qxmHs84NamtQsFfs6wyCEyjlC15gpFDSkdcS65XZ2Q8himHPUBCAA7AQ
rUXwijHfPVuhzLokru352u2wmoS566C0BQcTkSfPB6U2f10BdUZVMOv7ESc9Fu9p
c/IlKSzBi6fu3ScZ18O+pOkAP4Waef5eHUXDIpL56xv+2Nhmu+lKV8WplDl5DVgc
IDiGdJaBejjCuRb0rcUigGNSlk5xUfef0a829SwfquaowED5B9LwRULkIPyJgHqJ
Md1IA91g8/7EbjhZBGEmWlbvgQK9TmsQA911ZL3VKbRx+fpw0pS0kIHJCOrAecuX
hQDriXyzBGe02mCAiW2g3Wyma26RAk7U/x9Bbu0so7JighVoc895c2OdPrN8yVXF
/zHYcRDK8PGfXJphMEFUGZKxUVB+yJTgBBDA9SqWKc8KIw4inCyK9GQnOnJq99z3
VOlIt/biR0XgvzCcGv4+vpg3IsB4lm+yJNOcEKyCQUXZ1h0O4P8gbA4i2t4WsrHD
RsTEQHtgFgobG6sWVAWN6+4H74boqGMhjhRAK4MiEs5T9lkWMqKWyBwf9hqco8HN
BrLh/diMHlgtZ3mIzTUTrD9THkU7ABq7FO+MA0CnHZu00VB3dPSWQ/jDp2sxFNeW
29zimSiBO5vImfkTU+c63knj7e0Bik3+jnWGrqeBTrO6mVpem3+khRcK9D+PQzem
zFUXj0MRmgAptt8T/q21VWJwCNdglxTRIHSLiSAnY9NG0k9wAmpwrElN2dSZpD7r
2FSLmOEd5Ye90q8jsh1G/qV5W5fbw1kd8Equ2IKNi/a1O4pWcoE/O9e6ypqN5sb0
7t3InMESkKNxdjMom4FMRTl51ici8Q7gpJb/tB4XqWWK3BhlNVZ9EQvk0JqmW9ue
fGkiLidly5169aFA+SleWZtNp7jFNeHEQvgFxW/z4wveeOUe6UzqZGUElLOz+Y2G
vKCZYr+TzFtX1l8a9tQEkSXkobQNZEPJc+lEuN0kGrplkKDI89foV2HnySlkw6Mr
tLMLG8ykTP267UY+d6NIujc2ZEGUnrHdTJomAoh/JBZGVWwDmgHQJJiskNAmGUD5
qqNSttaKzSS96T3HxYK/OPLyc6NoTZ0QbAT5Wbh0cGBYoip/3AybkaujJv7G8F+/
vjN/L988Zxe2iDgirQ85EkGZopG4kBhqYBzZJ6KAYxlh1gDZbBvZnxSEYya3TkXg
JW+qj69TX5y5M1MFNgkZHopa/jrR9XUHNNJlMkLbiE3IbHziYHqh9Roy648Xc9MP
d5Dvs5zFbF1PZ3lfEM1jXTp1ljGJjywLCha4c413lH8G/H60kx/k4gYFF82j6S2s
sEuQczFJ3W7KauHVyRsZle12C914w5NJGPEa6ssZCTxrI307LzfuLgIYKyE3PVsE
/i4WDZP6fSo9pbDHLyq+BQ0vAO9wuvfjqcayyxQxZ8ptS+KmSINgiPjeV06nQzk5
mttz2Ik2b31k0qQw1DS+q5ixN6nT3YLPGKW45VTzZKxxIW0SfvAlbFBx/Ha9d2d5
rR6Fl5fjjpMqwrZ8fIEG9XVfMkiYq/92hOZT0bzyAwI2xLC1ECYn7vL/8yK5nrEW
wVUiqueeYGqkuPzs6sQEcEtbHb1/qQ+GsmPW8ZsuDotCY7ZVYINDy8eofZgldQGq
SFE7CJVOyCCBNDsj32NpUMfcqnHQm+67ChUDMWt9GYvstYXXdAC4TWcboUz8XI0w
9gJVSlL5vZXUgImxEITM2CzBxdcxFAkb3UVpDFIhw/AYRJ6yfrnXtdTAgSzX7DuN
EAWURB/093lklxB6K+kUNVGFBf2J5bctv8YOrpM6mtCFm55k28NFFS5syzjdLAtk
mZHeS67SU+LMSPlzQy6aT4tNGVIU9LTw4gnG/LOUDs3UZsKW3RPwlhVNd34SiEEw
GUDbujRtY8ge1Xur9F7n+3+dSETg+/BuegLjwdKbq5g6wIx7niB3NDw5kGbeS5ta
v0F6kd/Cfh89iCjEusoBZOZc6BZXbjLjshflJdoITGUev2fzIB+UZaDFX+xLG7rL
6O3H3N6WUa0L7k379n4GTPfe8cCjk4TRqe9SHPTIZc4hq8Ktt4gctnQf8J3ga4f8
5ZVwRnSQFCU/i1+f4pcjKgLZWZ7taQuLSjnCjjKk2mHAbHwHGRv4HPzmdDjFezI5
HzJJ4yXuE52YsWzZYdmgZkEjRpc1l5pPl2EkWAs40JSN+0wXkKok0JJzg/Yjjvcw
andGoZwngmuzHK/NWCSfMz7EWmSmb5eox2ZcF7Iyoa76Idm3k695FHBWWTWu+jZv
qJKVGksix2MtLBWsmFYlPv6sx4Rog4sxz8iIvfGaRCIKKkV/kO5j2Y5nRmhc8vjM
C0/HZK/jaG5iDSzTOv7pEQYykBbOhduArksZ9DD0uSxvlPtA9FV73+sUNl6r/gX9
VI4v4kl6C2dA+H7J3wedPBwJ15Gg4Dt7VF9Jj+WdXCRnVhu+ywm/FoO35ggTGLzl
xvw6HOIz9w7s+R81gUtZjBkZpEQGvCT3Pz9nyiRlHyH6Zvf0BX0af4srCzqNO0zF
XBqppnqYE6XncXjLhhidwPOShWkYMmHIC70Wg+gSxBs+tkEzYFyushSxSjxFQ/9x
hp4BgMKFoY4Rkep1VWbQ1DJKFrbuRmiIzeeqZFfPMUifK9GSdfLLqx0ItiQRBWz4
0CILbGnDaYpDLUqXHs6+y8yDvzse5pqFY/e/QzqhlwB/v0yiVeXSpuh7lpLOtjyE
4Ap1A3OHSeTKO0oNeRHyyZZqMQSHpu4p4hv+rK+hI1kHwM0PpREorEkkYxvzLK9u
7A8oD6IkI05m6J6Thsp3ymtYt+qktpBQ4+JOfEEwJV3jwJPWWsCkfHfeevJCnc26
j2psf0YwAWz3KfA43mrHeiN+UOOgvkeJ3JVGv+p5awP1aN7J8tLTZ4iM1gD/Hs/H
dPePve3974KAfg2gFzlqx3r1YKe9b4dAXqtSFuqyVJNp5Xk9l7DWcJlzetH1LTlO
kC+XRR9qVseObeF9O977+QUgoeG9u4PFWud75bf1id4pTkzXfRA4x2CwonjVBqrj
zxYKg7fLbohc0cJg3Fh2v5bjAsiOJ5kaVeGa5tyWNQCU9tYKReoozOPEKXhrLJOO
+pd2RzkiVJ/uLVCf9h+5oqXEujG21+7rtAPZtLB0sPqPWkhZKV4a8TFwUdQh3tWz
9KBa67ShXVy2JuiHRbuJU/gu0D3FPAUUcYDtfGrK2ALbgIZlJaGLS+Fek6VYNbl/
GQ1RsksdkAoyq1HvBmF8GDPC1jCHi7qMPLFdF0OndUzdjLkPJY+IWAuK4TCGmhNv
QXdG996fJmeYfhd4NmUnVKIZusVgB1Hx62oGakOGZ6uFpWccrpQJDufoChFTTMeb
cPLwkc0LL+ceQ8W/q67SA5uknIJ4aW8PpKRSWMKIlooaStcsK4ozcceiLUmfdx1b
44fUACJtBMw6s9BdiOPpNeMaCkOQylQU5xZW/R1BogH6BORWMf1pGLr5gyROkUlK
5mJAhimVtk7JK6tEhbpYbrCdAJgbf5itYajVpH+DlEvzizZfrhe/TTI+ZVrIzAfo
nDAbVA4M74XBrzkfy8VcPQUS12tennsNIi/ffv/TrG6g/LUPodABxYR2tUvdoE+e
jBXZuMcQdtzr7Vb0MFtCVt2WIpbwK9p/WMZD0MjwjZmPYZfmBYRO/Zh53AwSR/Nq
cx0es9BOZg0AxzvvVFWHB76ANXftVV9iEJmYBNGXvvbXi+oZMYBK8hvUlvSrpKfu
m1Fxpn5obt4GJjOfnVpDABYmuD83axvhZT5EUxjFMA3kXPUdlG6nrrMJQhtlJ/R3
kZqd0nXy8z+PA1VF5bEXCCzQl83AsLIU+iv0jXK+T2djDjDg5SIpV+jfu8PASKZM
zBbewZ2rKGtLY1OfNftB6WBMiJvimP7lc6+Jc/+xNEa7NsKarKgAXnJz5ojrZ0XC
vetfW+Exc4xR88BGcB7Ny1HOOh+wI49swY50OdRsZOcLdlwkpRlS/520HiQsO5bP
ptzjAn/kff+h7G+0aPCwDOu2Jya/xg4NsR3fBjUM25Ka9c30a7sTT7GZhJi0Qfi1
Gx5WCFZ6fuSTVXqzSjRaStmfbDBUxF1HS5Q5XaRB9YDtAD8jGC8/GyjHI9aMALIG
L7v/wHTlR+6q1/Cajt/J5+EPca+BbR80G/lX6bPbC9sZDMUGN3WDuemXSNU5ZZwK
J+0voIw4u5mf4LpezFKYQYi6PfF92OFc6Y/O0kv1o3+5spZnWlEPPcE4sv1pS6PC
nwOWvw2W2lCnm47kLq0re39tVS70aEC58wO5HTT5kSliA1LjwzuwKnbil36LQu0j
x8qITs1nJdSh6lNtnnMyfoxSmqnUnk6YhirC/qG+aJW3Zpj2gPDG0oVuJoz198Dt
Gzy+secgLoBzV8c7WyHvORJa9JCqqziZCUxHP/iAGGGQyTE/QrCcQ61AzbOY4dkL
od1rnHANeqn/EYTQ5/nFU7ujmVUdBdCTVbaa9cEJFRLYhDMqDC9FqCSjvfP48+fM
W7d7oiMw6B73Qt3CVVWUxJHJwlyHckmz3K3SWddzbUTVj4GqGI18nK6A4rIw6y6W
rok+6dtf8cuQkzL4HDhfO1pgH4LLS6Dh/6R+ebRAc2MZNEhha0BOrUX9TGd6l0YE
l+KHyspLwiGFT1j0yMbgtI3kfcSfnQGfv4SKZXBppaqMhWlHOoRU1ipOKq6Nq1YQ
4Qy7MchdrjtidlxX30qw1Qmowj685EY/lc9LcE/WP8QkKpjqaggSqjjO9aECtDlE
scuoN5d3btvSuRBaDPxMzk47wmRPrp2SG1zTzxXDuskQYePiLQIHAgLcpNgco+IW
XTddrJNmCRiyf9AQTx7/0NM5Ub99hyMguNVSo9z33Iuwdpf/pY5aiNDOYnN31Byg
dCO6hcKivU6/cYFQhFmnylfhTIqiRYggEMDB0y/QvyTJ/biCoTPmpHer4DSOcnIf
c91Vl1Q67hH1maHaiu8pvAEq/t4M+LMXGIgeNupmEWih96i6JeVkEbwuBt4jfXog
oi3VQXNm2W+4cRAHkFTaTlfKV0rieoQ+xJPEavUuk/3yGqNSLHQO1VoYRzXO4ABZ
j547PgJDkNCbjuYVmr+I/3etkV4D9p4We85unsuQfi13j2ATE+QE1qedPsxj3OHF
m+lKggi1Sp0Nw54eMU4hMfjL9fPAPZ0eHsmjfDhE/KsVO1fx5/kH5BXB7Gn0JFzW
eHtGcogBe+4TogBDFPHhZoI/0t8FwWOFsuuqeJxylGBvF2ziUKlf72Vj45zsTWIr
AHZudPNP8IAl9h1VPaDXpPuIO5q5FJhJYpdDHRUx6ZOJMtUUVtef+KlVb/FKxsQQ
7LBRxW7BtpmXTd5igxLfPNNFyKJMI85jznzeiMTU0w9VmJebSVQrP9+pqCoKMHUl
/NOKhWXTt2UzK7Ve/LGbX/Q5fI3e8cLfAmadvrvcJSgcMfZX79/ZaJRCCwn4Wiap
eFUxs6oClXp/33maAQKNlc4sf4inLjqZO81Jsqo+cPLDH/qj99VdnRdObNJfstfd
o38NQWa5g8u2Q9v/8hQrD9PSnsi160VKfIWr0A9XYUAQPTm2goom8bSjW0Z4v7rV
DPZ0ppFYmQ/chsuCBGtNp8nfwP2dPzHnEAXuMicLbUXrkFMUwY2X897uirnbPEML
mfyupmLregg3xIofH4hQaHEFc8x5HHUhUSErD4QAC5norgzjbHc93GCt0kJrHmwz
zYncib2RQbu1axWsNGvphCmXvwnSzEHXpjcshA926Pc2QlrNIdZFO2b4BL7YTbKl
/yHF/zrFEimt/v2cqcAtqnkK2gAMalwd255SbHw7Ti6nqHFlbb7YUWrz7QiNl1bb
SdJ1J27wdgUonlRT9JW0VDLunPUZdzUuX2FytD1xIxK6+ilhnjYCDEH9vTQmNoNK
v1xVC4dM8F25F3e5rX5AAc9dZ4EAljNFy5WS3DMMF3CMGgnnm1Y8p8+xhif3Uq+F
iIjXiY4GmS7IYeDkQ5WHlKtRvlEBrMpWGGdVZHiPBxB2RItT7krKr15T42EVG/dq
jSjF1FdAxeL2YYBoVUYvxFJ/QC2A6cynq0uQzJo35IJm8hNZUQmB42NEleMZU6EM
GFKovELFs/wzGNjjh4m71Ft0zNcqzb2c23C4sZMXTHLOzuqLmgoBd9F5LC/u36xJ
nAfQzq3obYNUrKnhL3fYhbNqswOe02Xca/eIr8PIb5iTp+NPfVJgcEVJD94geTMB
Ck+wMHjSIUVuz4rZL6FAQB22kpRkO2ndVWgOFKZ+MT/y0gn1j8KAH1JA0cotm7+U
ZcY/ubHFj8S+nSFqsNtv64vnOq6mcvkq7F+he1xAOEqTOmGUWstNNMh82sH4oTGc
SvXacAfxCgIk8DgRyBCaz5CR3aykkykiMzj2VySzipxH+lQufMVAE+GsH7csCc+D
Fn78foGSphcPwEmbN5HkH7jDDBEAL/78QxQt6uxXTV70vdsbHdov/8QlRb5aF2ZJ
QuF1SnqoPcv/Mp0FgNRGZ29eXuFFdHYdAxfZ3BZm30DXLuIBL8ve8Vgl5vRSNrPh
yM/Ga1owCSdHuBFuwx8Hwk4EvCXss8yrZSsmxYKqGW7rnBQDO8GmDEPYBElIMwhF
3NdOrPjO2qqpdPrSYEWRmwhmQO4a8Y2yNd3KLHuh8eJxhPFhWb3v7UeTY4C4oM+K
OQJ5HvmWQeSe+aqG3i1w4ruEP7NTFCQsNnCiJFR7Of0Pv04TFkgrDcZ01bbLtNfV
RvUKA/Ebey+ZR5mvWoutnLevEujLc1suaniLKuY44ZMp9FKMAfRJnpZR9VWbrXEF
U4E63XNbs47PKRJS/Q9MUSptxSOCJUkxFFx7R99Em1sUq64b1wlVc46DKLr2mo1P
lpYfKA8PX7lMx7+oYMrSzLNYPLhjIUvbt5hXdA6FeoOi6lMWNgogHadGR83VLuUu
LEajgO4mCru+sNakJtr6x+Y790z6skkXCFK4qzUdbnj45DO3776N96EizYXDIYnb
abuRsUnPFJ6r5mNphQ023vGDdZLQWjlmHHXCHux+vZwWBCgG2qzti2+0+pG4BhUO
E80dJmZGsEMLCnHgebfzAom7IY9dZRbyZy2ta1kE3NKTPGBE1BDUQvUwWyD1BVQE
mk8iDg0WcnC7Ky7ZOHqOY1yxhw60IRQkIoHSmyd4Im+twi5cNuqgbcwId38XC9dq
0L7CAmyPAh72VcOUk+QEklSxx7UJFnwNjH/PePrxDFz5/nUM/3LPfVOTD0tF6qhl
yahHpJELcwkgdSMSnCwe6eZBuUtbcB/gDoSUZQ5O5DzQz6etG1iWlHR2cyXgsSYs
AEXOUpgCbb6MgNnvb5YPvmQSo7ZrOSJ6qiw0HuyEoacL5oLEuGPiEIFCTT63G6rz
8/+dwkIiAYnzvluzXcOghTbFkYvJ6GRxWgakWnBgB26KLmmYpU9Jvok5kAOeBf04
7iERKefCHyvdVffIUY0mshl8+jRMP7lsLK9zvbuzIJW4HvXKa7sBCWW9RnkVj+cW
nL5nnXSZLnaHWTpaK2zjG0UVZpSp/0XFygMqsljrZ+Un+P7DjugRoU4JPgu6VzAm
zrmDnvK9Sif6eI1UKmR1KNwSNQn5pgH1Q96+AHBJCltks+PiHBzrmN7bszg7NNdl
yqi/aNtZCR5pU1HdcYns+nEy6VwbwEahvjgHqAlLp5NGvgXA96M8GIOqlAuplkwN
99lL6J/c59DbXW/XQlquRUDdBZeO4PHC5uZN5O6NRYdYP5dR+GQbcLLNjgShrO87
XiM1/UkqmXElCOlCWkvmzZh1rKBOXXAUzTbQ1TIv9bIAEuKoZ0FxLb4cmkiYFC1i
YfzTD5PVsaOZkS4juaykgeQNMX69t04+hvx5U65bKc/reNkUiyesBWhWdSTh03WU
zwRGBFGG1beHpEFFFfHngwLS/oUjd7vQZFsdmCiRh4Z00YxdbKxe+WAiF275H02T
0evAmr+8kHnkLfhoL4pIQd0Lx6izjGlUGLDMiIJeVA+ZGrvTsUXHsU06JQHoky/r
tOfk8m8CqmodEyslLE2h9NnksmC8jc4TOdsALqUSU73AS9GP0X7Evs95nkC0Wz4x
DRs8YUe3EIpkjtnmasCOMdgxBlTh05+m8nOwKxIzNpYJkEbGGuV1Tav1aTCmPuZ1
JyD2P4WR8bKxZFH5F3VO4cFRlxQNHX8LxeJVYP3GxqI19mjD0QRxTayUMrHkPgWe
EIKmwGCwLx021Eqs+EWwEeObu/A64qVYh7f+eRzowUIkqV95xypFtCxsK/nZmAFG
lzxU61tQONrejXsbj3fyzuMIuBSk46dKzc+JeKn5oK98zPXsFjI0ZdlwU8+N+Qy9
zP4uOsF5N57PtGDaBsalt42Txb6DXYicHO8O/CakqXHfCMx84Stf8m20dzqmHsG2
9Vk6KwDuoSgEC4EjOMKhdswPuEWowYcH+PTaKQMQq6IzSlWvF0B2Pz9xkjYVML2R
xSCID8tLMKf6V1PoNrN3Yy+W12hxTFkHN2fAKvWv5DSTV0vnAVaLGM2M2vxIYz3m
9qnYDNgSy9tJSa8lAlFoafCUoY6+wV/dYGI0ROM7tkJBHG+nPaWS+Urzy9wpCeai
d2twwNWp2uyJ9AAoEOsvGB4rwjzP2YX1DumbEOfvAcZTgxx87V3Sr0FIX9pNiqRS
8X7C6weRSCHgruFhSQ6uSay6nPVb4ae9NlUm+05tv1H/avSpudL4XZnWhSg3ObIv
uFTaG8aevPEKHR95r7BDu38Qifh/XPR11H0vXGN1x+auVp654x8RmIt4KCT/bo1v
tOjQFRRWvNRM+sq1Jg036TF64gBqj5BhufE6627sVWO0hD0iHS6TJBvcWUHm+hDG
NJjbtgg/Ip3Oj32MEGydTw==
`pragma protect end_protected
