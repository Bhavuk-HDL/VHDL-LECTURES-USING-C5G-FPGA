// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
PmhbTb7SjeYxP5Ss4XqUSp+qfL9tUq8b/fmaENSPmtGrIlf/NctdRPN2wVzQwFcqvZM2lpqRB+nN
73+Pf/j8PuUu342eBL9geofbcikPcOL0ISyOrd492nGxVn4hLcjOtLb5FFYYQwoh8LOSK09gdb8w
r/6zCQLqfTbao90mCUcTTZ1d9iz5IZXq5FMAguFxgBfNVYyHS/3OooDlQVgRgNNAUOoNhHLYfO5J
N9mNzQSRZ2IAvyshVGnhllfCiWGdrpKwte6VWfCMr3CNzM4cLQg1E8/aJ0N/yCBmGfQ8RCWUNIkW
o6BfRmmQgqUI/+yvBVLKAFQAQS6IGtA056Nl3g==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 13744)
uenh9X94PnmfEBqLqORrqPEywDksPYKuWl4k+xvRAINPuEQ8BYmUyTyV/EMacbk73r4+r8Q80oN2
IYNxMbkb+tB/yqVG5qfuuKhm1qrYOTisOF+hWOtXuadmav0L6plzQyCnIVo8G9JoPdk76j+DJpL3
fr/4ikjnWAydxTgVn1viooY3ROCTeN+egIst9cy5G09mLX50S9AT5weFA819hHDHFRxthD75kBGp
jtfhLuJBAI/wFl4hUO7UhYuVPpbd9oqi04onz9w8EXzecKY0m7bFTwWhh1KBLywx8X6vNoYBf+8m
/glSUboEh+Q9e05vjR5ogXg/6oP3EYEpsVGvXT5oxkffaZr/E4hv6Hx54f88fiD9YwnNkF52fdwu
m6qdGK21CTB+5tcTobuYWEMcgf6R/OtTQ/MSreVA8y+S3HEOqcS8lEWA6lFIGznpCSaKClrsTM5Y
qafD2WQS65tGzzYPagf/ayXM1rL0HIgYpwiIXyB/3eC/1Nuze5EZmkAqcOplTRuA2OsBoEzvFe40
XolMaSzj6wS0p9vFwiSSd6sTrz4g/DzSvYGYfvGF34lJ+iFTmjzw3EuOf8sPbcVNVIwBElO40xsk
Sn6qR59dcdxfPd0s8uelvldyUTIUFIgK5oe54eO0FgKLfOWvWB5kdzdkwG4CVfYjKTy8NZpwJwa3
Yp5ofe6RFZD5kF5/PgiFUvlE80ybmbccFHOtD7krqz9TD4iYEC+Utc6anxT4CxuEQqT4dvpzUtb0
x9okVMIrsgCG0LsI2SxWC/nkXO3ysA3+xflrj1Y0Tlo9WsCg/Jw+ENiytKPtGhhwOrXvvEZ0yJG5
YFYNsTa1+DQJYONB7jHlQyoCpN0CDA5Bo/RO+U7fx0X0w17qdY5J6oZYJ6rxrEvERFHHEvUTwsIc
seoHu2xkM6rKyKmrpicV9EAWgBOmG8IjjO8BEFk6V/F/M+AdvoCHMVKsSn5WdqIGtPAzK3fHf0qq
LHoF1PfEl0mi1p18HZ5VSS4LjDl8DaR/3EdMEqk7oMvy2CkGXMGG0Pq4XSZ+l4uXhmag8IogweMG
9/b8JB5miryras0ZcfSgWLVJqr+Xr3eTiZHmtysoytOTByWds6XL1xKc3YF39WdB8NNLW27Yeaj1
V2RTsvF8vAFtUQeakzwSXLjEaFzkAgBUPZA0Y+ATNrAPeVz5lFyEGLoSe8symfN3GP+dcn2DYGYP
pgHuviGPl/1e19/VmyLn1Oj8DruCWaQNXllqN+TYTYjmbcrlEMRu52jQNqa6txv7bL0x+4wEgrdZ
R9l1GirbIDFg0UkQ9eCW1/rmaCescVI56x6om0I+m9az0ZYwZ9Bn1QSDhQB/pyLQJAz4nOTHBbBF
E78zC+ztX24JOv6mk8w06+PVdACuizxVadyRx0WCAW8yQQ9fGjx8Vcpd36+3KnpMcdHxESVsanIw
3xadYlyKF2MDg5wyJKg3m+FtuesrjnKqzFaY7xVWECzuzYHLo6IIWU5RnwrFajsjQBrwy95HcCyU
DPEinAUioifvI795bNR6BE7MF/RqIXtZMJIR7zRQKOjGsHmLPf0N//w06XlJ1rZaxS9LfBBuZOhC
OlatFRGeJ7i1ETZMUH5mgyrkxlEqM+PVvsnZNx86u5+X6kF99SN/tRu5jyNzmQI9Ko3q3puHszuv
JcFDKltoqRdaeY3mY0wXBzWI2FCVURATe4lSAe1jxdTANMEHziRk8d8iVp2CkxEcHOQZH1N9gtyO
1/IcWp2S8NVzceCh4goWkVJXZOsrESX4LefRbdZPpJv17FiaUvf4StXW20H1xnmcB72AGULFcoog
/jM10n9RfHPxeoVIyCnV91SqkOxBtKlbh/L3LKOIAvTwMHvxhUNMnQAiUfxyEFDxDq5FiluIiBJJ
FbQOBwh3S2QTMVdReqBcCJF+itkWsEV+ht/jKBXjybXesg3AwwnN6BxnnezPqIIcwN3MTcU9J5j5
xVqlvK1Tkuu462l6XqVl4ikcRNTFOP4FYCWPXQxsjccorhYvXDoBIH1/5bDzhTiTGgPRfJuNDYU0
9JY9O5twF5J8X+gXY7iZyt8F2yeORkex52jY2E5SvBoaKGGuusEbDBZmUvK8v01Cuq6ZdXVf3qZn
6DxohNDd/cAAMmI0XT+Q+rFdUb6XdtjljQ7b0NoWFk91Uf1rZQ+KR2hzh5b71JYYCgwzls8/7s1D
PBstNsTA8kszz3/3K5ETsg3TuXxQN/XrgSJcb6hnEpZW55TCq5RDFTvleuTPwS8E9M2h6kwFgGFM
Z/as8O0aK+zaGwyVHZOtPh2vnW1VmgeMzNBGMztI4A9Ga2MVyAdfpaxg2q0CO1O7OpZwTPL1IPwC
vBC0dqCUp3qBezzwlM3FwWld2C5kLN4deBxEx1ZeNRDPV5ouapAYdFmwMaFuceihPvzJUrBu9Nt1
09w2Ay8QQh1ZkrAj+iUJaEZ9BVGc8Z596Qk6mrQ/xPe/pLzBgXY57q+JHaG1RqTHr5EdGWz65a1/
v9UmWmW/hLpD6i2B1zPg77k3KguoI9xcfFhsmj6IVaVZrA52ut/fNImB6DyJ+q5z9LIc8uqgiMBm
AZeiSdxHEueFU9EwP2RgVTl6PLY91yMSqwp2HCQypsg2dityyoY8DLJrIOaAGJU6E73r78Eq5VKP
mLGIQER0b1xArsIQ9WCxtuAk1e9IiS7xLKBHfS8q4Eaqy4pkdDnfs7QvdNdV7rcAcpCDORUkTw7D
4u6NbTwXTj4qE/a9s35vp3ZoVwbuY/58H/bvE+H10s9xdSY8kmD7Y/4ciDyBvv1r7+onfJK57p0n
n9ySR5OYI9OD3XhK77DIzvAO+rtUv5RsdLVVvAWjF9KTKjz9xtjAUxOTNb4WYLbKTlrn/+RJ/Dul
1cYmqU+lA4KL1FQlcpc7uVKAbCa7R1IbBW6RZ7j/8VtNO8EkdAYQLAa0SiTHHlbIph3isJ1Uin0g
+LEmtgQu2vI356FpyuoeXs9+opqYGnuCvxW19htrSGRZA3T52FN6H7vsZVdRTh7cyaQvMliAAm+L
Sc/HKom0f8fM1JiLFFSCAAD8LLncI8igZ6jpPTZK6KnA/PhB4BRHfjYzigy3/6Vep5L8zEx8+8eJ
yHmRNymZq0O+hEqVfVkGL0zh9uFtaoRnLpyapC3T5911vg+lSAPs/ILFKy7q4/qrGPx0Wxe9PTVj
214gL6Ai9gCBAFHks4dvVS/zW/gO/lwRYTbLRG3MRelLiCB95cOlQ6etlJX/dXr7C6rBpyB/MAce
9QMa1OntEEyRId07nSxSsbWY2EA+Bth5+PCDD8SUYz9bY/VFy02pI6eDz3HEqDE3YYvZcZ18ZNb5
fSKXPfMWPSmHOlEC126kAF9Ys/iz+ZX1u/Axccg3OKtVsigiZaukVI3uLlR1Jjm8TOxHu/UKQktx
9VsuIwcM7MZGbgvasPXj9DmmkuD0MCetxuG0xX8T75rHCF7t2M66sJatsruRfwnAlAKMA55+z7s3
gC0bwwsJy73aBOlO5hlTWFOnhS7dn/xUKKEI7YGGRJmLGmAQlkSf1yCobcqHid4THisAzlEI8eqH
6GLrK1fxxL334clm7JMpK4Bbu1TyqNEX3rGWMvclrrn/HGOpZRKJG60/tqPOgZ0nBPbY0YY0A+Jc
ppof1Sp0bjjaRYpr8p9xzpz/JVyZy/MQM67eC2o83nHWktvC6VJMEJ4cxhKONrKv89SJoTOYddDZ
f/+AJWAc2+6tRa8FzwBghKKlopIM0tRzyByRWkA7tfoEILSsOb61o2bYV7A00oCZCWYUaBA+9e3r
jZuZY7tzoS49qg9yv1xXn/ApOH0cNKj6i4vXWprLGK0FqeoVjF5TjaMnjqKKQhhzS5rqBca4b3ZS
y2B3LS6pgSnTu191X3mgOZiSzYo+Q6Tws7YvEEqI6jsjTajbn+vPcnrX/Tp26N2HcFcB9Yp4W4+d
ouRd9kLdns0ExhvhtvCcECr113FGsH4J2BKzRKbZLlYG3jetiiZkl2kWL2iD3NSf3WafIrBKt7hO
eK4Bg8p3HY+P4gBk+s02F/tcvp5NKIHB7JuM6WI+aNkVbNIvfyYByvSWb9X6d4DuM89h/fjtbV/G
CCZ15+YH/f1NV8WiQ/ISPdCIMbqJZh+LfAFfZiZpYdK3FXaBdGxMZI0Zax/Q1VjTZ5kbL86/BINm
N/YjWsfXynD1IE0iWGC/mzhseKUhiHFkYCjOcMw8NBISFRRful+UsKHtrt4/81M0m3QIIX0/Y08K
3hgUnBw8AoGxr+nzCWomfwS8Z32+BC8Ir8BMTDoS/w56+4VQCRASsMRWFC7mt1SyanNjILjUp6Pd
UVFj4E7JDR7O61Pgfe9s6m6Z3yjZPUBKcDJ/RtjtwJ6RBRSt02Q2kgP5MhO1o+Kg/l2A+iDs5SeS
UFT+KAVxY0Acp7PAIThC8rD40B/5K/Ecl/cDxT+pxntSp3XYDKhzinIDCjlZuCYNOmU9BbvbDgPQ
K115a8sUhPesyoH0t4Vd+DHwt7ihA+r5w+3O+dv4ZYHjsD4AajCGDHRXJRxoC38VRs5pr2SJLvA2
MtxXcXqC9P3iSSzXWVxTLvdlYwcCeSA7mg6WC3BietswP4CwUyjw2REGb4I62k6eFBsXI5yvaA7o
Ebj9RWW85lcSh1ezQGqAF+yScLXa01xMn4JxxejKSI5GwvAtq60C4UR7dYZlZjF6vjgJSI2/V1A7
00DT0HGWhWeBz/HTPsSv/X2qmgs/GVLAXbIcnlbez0Q28CaM9RVaD0iPvZBEVkSX5YlyP35PO9tD
F57ocrJVDNOf08fQLXoSc7SCdlkd0xdwSW7W+A//keKquHZajQGY1oosb88Z9VCse8TkX1WXrMPv
F42Kge7ZIfCSpCh3hLRouFYpHuEvMFK4B6qMGaqvmytnajgMmGMsNG0MfQ5suS+TGu6R1fwHKTri
X6p5eiGuFCzll7f2mZCq1HXAsVOrwxrHL55vY7zWhjF9wPuuiUTNwT8xFT1BWcqIB+rAtMRtD0Ex
PL09Ce64E+hfKnxKVVcCUouTWfhu16BT0dbz0xIj8g5cgNFoDwcrE/Yxz7H9mMamj+nnOWVuTNom
RZaRHb/uTOAyNH59FbIIaHdsiqVuB2Oqlb7EntbQbB/WcfDWc5xRpW/0NYGcXP09Ix9LCGceGN83
hF6vybwOukdkb++TjY4PIxo4jmSJ5KnQwx+eRMdoUzK6VgqlWsHxqZAPZ/9pqLisS6m0Epdvpuvq
GeU2LUNkebMWRVy3+kGTgnsDCNhyGWDRKXsvgIGYv01MQZap6hNPt0MmCNe6VxB2+V/uV5kA8HLY
qSezdTsjorOk0ZBt//m1KMv8QMKOgMS3a0SMWN1FJafYGJ7IrV6Rcls/EDUq66g5Zx9PdkVs+b/M
hY2931sS5VJa0wRWo4tW9l7F9MSbZ+y7JUmdz0PFMFvBOi1XGFXI6QbKz4+jTHZctm40ZPWQr+Hu
nNFh4hSeg9SUqHE9lh49jwXlkSK0GLnlskQkshTux5JuD6BVSBruIhaFf7eJm08JvthhU/dkDKEP
sQ7L/AoaiKL7qg4QLXIu0K+HBsC+EI7bSX1k5BpfdzysR/wIPrq7aG0drjzU5D36+GoByHcCScBk
T+Vn91pbFs1X2bD8Ot0Nj6DdQONt1Hu0MvrFwoNhjCZPWMCTRfNNhsKNywoIjg4xnZ5rpZMovE7t
z2eX/NLKZmFrJ8FA1XWyJ9RbGr3gcjbMSn/ZoczfWA2V7XwlWV8NIQ4epJSWLONqC4kiDDNvQ3mb
JiSqkYYA4ZiFX7HlngKTpFzbu3+4ddm3o5As02M1pal6YJiiYb61gdGSJlQQEbY31tRdEGP/IVQW
RItXu9cSH09KgjubmXzbcFY67b1GA34QRsn9j764JcRCLppnAHzmSqAjqNThsTPIDfy/+fjD0wIf
kUXzLtGn2/ab9qx3jJvNJHZLP4FAVCBD8q9+ObpGtkslg7ApK7SCti6pmppyNEWyNYCP3UCO9kY3
eSyypDRVypXFJsTk+xwljvMWnjgBRa/cdq/RPAISn3cr2JEhOn55oaNvY9ueTMuCpNEZw2GKOTom
3YOLwOCs+NpU+Jjr/M28YCAra6oMvTClvWel89hU0yIXmsvg1uOv7uNqRdpuB7NylvxLAKkrjmWs
BqMJi8DmpTK2SWeA2yw2NwKFvE3yhCB8t6BbQ+LQCkfAeyiT5XYZWXNhakOSioF9pHE/kpiZab7e
uSvkad3Q8n1tNafHr1/Ti3xF8oz5h3SqgNYmsLY5OmUiL6jE63LATrCmOeDm0CcbymQK3cmBhytS
DjoGLKSEV66txRymmVQYRsEFYk8/gZpLtB6uKVG+ByBvR8mrc3+WDvyO4VS4V9TS0zAfTzfQUd45
OfI7rE6Bq1z/tETABroXxK19lroXDX5+/vVtQjWkQC6bAPycgumx7DZvX0JGt1TEHjVDcY4sv94h
CTHlN6/mZXPfjoQV3LL+YY65E1Xyx9PzGoymwJ8mgUblNRiW9w/iI3jOC2+Rw1dXJRvJO4d0Xb0s
DlEC9ewDpk61+ymLQP5PUkcV9Ujcp/kDHtXGFgJDZaMmuG+zE12dyO2GU4vDWShp2NPwx8jph6V9
NiNnFrt7Mqe+8up3cSJbhtzLLVRO3BzfS5IsGj1924B1CKRt7e6xOjUDjbyFNMihZYd0C7ql0yrZ
McDHQHSIobZDdt9CkviwHgeMbrLw4m+IFDdOvXjqdegCNeBNbHn5f/0BnPfjLswmEc449Qimd1KW
pCERu2xRobghhvdZOGS628lWFmd2eSZ4Ze3fd26/R1/53tP12SzBoC2fYglhjWI1xBwl1M5VUNVn
R6FpTNkSZdQzpyfDC0dvOPD+KtLylh5OvqBY2DD4wwsiADg4pwYHuLQOEDSqZmXVi/SOF7dqMCui
IkSlwlkl7qDzwuc6vKsnkHYlnDsKyRT9Tptc1KjHEfffnju2xqpAfC7ryeUAwhln+vUkb8vyAu3I
EsArXkS1y7PdABpFmQRW4/Jtyxav30NtqTnD8rRTMVZCTQGqR4058kcRCY/l94kmNEntiRAF+dIb
e+dZgctMe5ZhTt8O2vQ3imNPcTCC2bTvOafrmxHBiW+PTb9T2kr/HMrV7K7x1O4DGc6HLyjoGixD
ApI+Mir4CTOdU8nSO1W2jFObihTuiHLSH+b6LftsAzAfaG+0QCUIaeqBuwus7WRWWGS4WvofYzfZ
B8M3IhQWav76rEWb2yFbUm0sTby3HU91Rka9NABa1h14IdHyyPQnVha4ecoBUsqTQ0i/Ny7geq11
uAiLSmgA5Da91rVVrLyYM5+Vb9mvBb6qhhoQo5Jn6Sq63vHvQBeE0GxWEr23X5VgbxbCTImqmyOW
KnKvQq6vKodMDBdE3ZnwsBtXxrZdvKQKgNj6RWGw04Nx8nWLQMKK1kbHQjX54DLaPGuPmUCsbeTc
aNOiEflCU5KijiEv5+VneKIM9nsYUWA8sri8n9IjlDYByOlPdwvWKTcO69OXPWRRj2HFjyuC1B+J
xmZmp4JR/36JlneNe3VBJZhjZdm6WYojISMhvcC60DLMuB5KWMFaLS8abB0wl7D1NPc79IWwys1T
SbBDJ0GNMhfOPWO1Sx2L7enjDSwagPmJzy+iz5CaNG+gRK3Dw8Oew3HGNAyBK2dcuXwxsDAXk9pX
yLi0SStQe2aWixx98Tdcv5LI9yP5dRK6wHSJZ/nSkU1A3DIeoVJbz2cqKbdCHTB/WMYAjiSMzurb
RxeK1Pqd1X+7kKNJrgEsF1hvD9QgF42Mt/dRQwpsC7QaFCYrnJXx/EQqGutM3i0jnND1mJ06bHlo
2Pr2nhWiI03kRBo11U808tD+R3z0vLKljpEyUveB13eGjtUdKa/QmSLHCMzm5EfskrGx9SHNwcUd
1pRzBvVII73u+JqUmXAkS0onToHP4DBaVYiHcP3aRGzYcJ9YabOnAxektS0Rprl2pf2fMAy1T8Bx
5wa+Pn0+sgyAF+xvLaPqqd7reQnBYVU4G2hf6m2BN7KvPJ5wZqIgrhwnKVZwGBFQm0ub2y+bv6H0
Wfs7yUE2v/8Yx/HA2Xtw4buEHPs8yljGJ+9LF32xG37yC/uaFOgnBpejJDMiFnPOqR8WeQBUDGni
qG8fbqs53haXEQ2HVcwsqRQjOAdhp0CltVZq8sPmBqGN4ZnbCErTywY3jYnWJ3xHje6A7bNDg6vJ
JwAhCIO312qqvg3xyD7Cdj5a7x92s8Vgrp0fKekM7HUCtz4/84JrF0MwyleynE384SGkLNPpTsN3
sUtxvb19MlfPqgGKKgYknXeFLXKpmva8n9G9p1X35NggKvHdcZdE/YOPRNqUZl6g/pK+fyhyIJpF
6tO6Fgk3Syb77IHJkl3qqI93XWzZHnwGKGQ3nVHrxTOB70yjRo8vr2LZsOLMlkSJ/3rwlmJg5pvG
6e6Ebll59Z18uA1wUSjf+hF27NGXdj0n41qqd8UKRDWoiyVI/SRvN1oFgRDPnECfgnSzLKwhT/0x
8oCJGyEVgsK8YaHcf62VHcIjRT+YXfMTF+nLKv7c7u9zeb0M0qYmaivYnH45rZJ8vO/ckaufgdmQ
9o6OkxDhkdMyW2pUux8ZW+0/HKuzczy2BcfapsC6nzwW48VM54TDzqXLN4SUks0HxALI1LUDZ8Dq
6F6ANPrAFjzYXSdgzcTkI4FHK/c+LCy018WKm/kGtH9B7JZtnhEehnW66PuvW0yN2vMTXsKIokdw
ByuYuH+/H49j/eYxW5qRl93X8qgpGFdaYBQ/vJ0Yzqt3ptOrReprX6jnMtsDB8R1E50ATMPUT3+x
T+0zQ8FZ0dU9KCfdOB3ZfVYvx8wn9dVsZU6GExrPyNhyPkR2J+cKaPmOlVnpi+N6KR8WmmYp7Lgz
4LD9CJsXhDGsbwHjU61eP8DSqft+ttx8VL81eY5rUfj2yOyBOVWhjdmUd9iazu3YvoWgarZCLu9b
Q6BjL3CjjMQ5Z8BkktVNpQ/BhtaXL9egPQiwu6gCFlzqlWh4buHjAWwXYdpqZzsl3lsbyI+Tj+Bw
0q8MuzM2q6tZYHP1F9JPkSY0Ax30nzfkR7QmaS5ZY0IcesNCmrLPDbnO/qffLHSOWUF0GnrCrIBN
1o6xEqFHWZTP6IIEZGxwL/o6s4DcMCTmZHAiOIJYy+NHOoW7359jr2h/P4z1DkHtYshUxIL3shvG
DeOktJ2HiPlYu/ucNIUV2dvv2y8nFEzVTEYKl7onFvF7FSoXnAnQ4K3gJiS9uwkKZy4nb0QqLQrd
hKur8WsfuqaJn57wPGSQrjq3NRGbcBjtoC32V50Y864P90RajDV2b5XjVROD4zfs6YGLsDs9WtBV
6bqdCLFf4QbEOH9RVXZX3pAAuHnEQjIi2orP25vaEDBbHSbwh8ccFC+piKKAlcrscvhw3b2T1YKY
9UOs3pPkbIXgPMhydRrP2sqFIbdUEdEbhWhtZcOZpVj27MFXoYz8Dsi8RKPpdzGQ33V5NkSlQmJk
wx1OmtuMz8dZu+CR+2EHjMK8PRPR7pFIePWKuXCIHP+qcGTIue4F0bZzVGo7xOHKeX0LmbmuuqgY
hNE9+gtK66A9goZpUNyJdz+YCA7fwVgaZCIAXbPmQ5mUhnD1Gp+52V52yFeOYXcQPRXO2ahCmTHF
sRUjwjiAi8bjo8+PvZihmyeLlk/Qdxox9cHrEp4d1AyrxzXyLxZuGJd9wN88vgVUxXjYdQE1+7hT
8KNNQOM9lIUFmtZfah5wKu6axHq1d3b5m6875u+fW/upIVDspwoUdke3zKve8FsTkS0652nJYDOk
+wmoOR+1Y0mbBcclRhk0TjhHlD/nm3iQehvwMUrctu2sATwJRNCGJrDlcwnbtt+tnEYBQYjLduXJ
H1HKKWY3J4OXiFOqn9bMdoK/n1e2Bs/sZDwk+XNbDeqwiq6uBstxl42moiUysxheTTmGYHICLWWT
z90V0C3FeNK/ER0gvhT38sQGgO598AS9qLqNbE7T581kzdcY2l0wc6zA/AmyWFk8QuVB5bv2weQf
yq+1DF8tzHIuMQixrV5hmR3AN4vpnK73rPr4aG1FRDEShvYnOD5P6Mu1wntg1KurUSb4BOUhFeHn
sx3oORRw/+HNhedWEwGf0NfMweq+v40pWPeL+2aJ7roH7oQitDufgo0lGLHfbnxhfJxoU2NIzeVc
eWC0hoK49qlPkv4raHdd0vcEA/e9RUb2FTY3qRRWBOJn2D3FwSd3raJ+KLIRLEYbly6VUBO5PzVV
X7c2X6xbS014lrUUev9lCSWuaNdPDIrdnJ2zeXj0UgebhVHyPHwuYS3LlyQi4T7YcM9XIJEId/Js
AptY+ZqE/E7ndqoVLB4/WFx4wIpKLVUH/wkpTzOo3mkR3v+znA+NRrJUeo/QGDNyqgesY2OjSfTC
OQn0jTn7DlUugrJfNHOA+pawFIIbs32CVGqZZ8T+TVLTvP4+bhjbtfjcTgMDz1MUtlJCa8H7dLkk
rctbq0s2Wf6OVn1u0k3W9vAR5tUjK3+x5nCk/bZUKTg6V2gkq3EpNGD1VRTWfxGQ3qhlSf2ZzXym
mitzrWuZgiZM4l8TbLtygrZzNHv9VVPPj3PxRzoqS2f/vuNB695gMqSu8JqcPDj7hKmrhrgux0YB
w2cqdDbMjLa+Vwt1haqydy7dMnPLd2ipUTUybNNG1ASw+2jwKQ8NsENFRhyHeyfXeewd/flP7XAA
sNM568ynww4HHccBetYcRjGdxg3wu4n/TSoehKIQW/vCbNzwGAoPwrchV40HVdhEwJV9P+mr1V7O
/WD9Ya2qj6rDgAF8G8dzymsjTxg63l1ebJtNqTAMvETLpjRj9LpBqIM10R87YRMoG3eiGnbqcdh/
ag1ysZ1X0uSTXOckCyfhTYZy3Sucvh2NbzFG31Xca7bugql1YEnCvby8HM1biuHW6HymX9pAGeRR
NzS+6+uI2qbtJllo68YEqUogMh89fMLfRplyL3alzGmONXac+f7Uc2l85KPjeqCojzemNX6a2jNw
QzyFdXnnFGtyJmXbRTtnZ+KoDCCPxJQl3RRyQoVYGP5AWrPVobcolQ/mMF6ZvU3NXhRDyDP2WllS
QKcAf0+d7TYEau3XBYtLLM49Y/KeqcqqPvfir4WCiP0ZZYp/T7Lvt3HrnYpywG0VtGlePDE/dENf
Z3tj2x66ZkClvqTEXZyRTvGdWpoLkyKUs4SKFh3h8+ffDmcBmroeYgnwDkRq4ApfGfNSIZUw0yPM
jEhVyLcjBnc8J4mN3WvNqFaNjDJBdWorY+3RGGgyapfm7vUeZdGwb2APKAVaQ/OSmurF0v8lyj80
sf5ueWoLL1dXGLs7YjyoosYbD4HA3GmtKCiIOTG3LsrsM6/KqRgQMVj6kF49fHbuB/oYgrmkOuoM
Cq+zHikeXXqPqrkZdA2IddRsxEq8rdXX2V+KIXaY1Fonh3HySZAGghFbeErxFBzmV6ujy84pw6bB
P5kx5k9cWdsPuLmOBLuqRS++6a6r7xEZuJqLDy9RFXwrouE0Bpfv5II7f+dQIZELTzhnx+YaEh1e
TXuQI4arCUKgZW4A9C15Ewo1XYfITrcCC+KjzGHTBJvsmMTbzt5wdFb4sEc9fDZl2/HUe00sIaWX
kpil/bqXtdzJeUKuaUa51ebiJqCNubXQtustTPOHLB8eHPSMyZC2PDYC+TPu97bcIGMDhQNbY4Qi
FyPJQfKhc02RUMT6ddTWjGruQpH+lEDYMUE35sHwVWvRl8SJwFL+J4pyAD1lM9Dk8O0IuI0DFEMg
wnfih9cmj2KSZZzuCaxMgL8psMhlnKM3l7AmV6vau4hd5X3MXO8scFPFxmQ4PwO6pkTwrj2Q1nne
hoCOyO6Tejk4XE0Gf8spsI2VG1HmWlVYq8RpyFsd98e83fj/xzyjaNLB82N4NEpoHXxHXPrZ3meh
7OB4MAieUeISIxTSV6YxC+9T52upI5re5iPHs7I6N8LnsmRcGX1ayFo0kkZlLZtXMx/WsIM2dlyy
FWnHzFnk+JonbL63bG+5Pt0gn/85aCI39M3RicGEFZaEFGblpu4i9vdY/jKyAZJTqtktH6aj0IpZ
nWRrDwi3qMFZq5LN0azBL64Hxqu4eGrRn+12MpZserp4j715kjJ+l40i3bvh9qkc+xb7diqC91Zd
uINxhUlquu6O6XaCqtJGCOw/19RwlLirw0bjbHRLIZ4fzHsxaWjh32HExIGoMM1Z7mlAMXJZa5KO
08s2/f4XF4OZS9I1CmwPKlp6jDX3QHFmWpwvVH+LoU7XOzUvzr2oBxAX8rkvhyKdbzSQHRUwBy2c
w+K43RPKMwk9yiUqn/NtqqB6fo7tba02en4f79DuzoTjz4ZBGOXbQ+eIpPrX7d531NnrUzKBzysY
19JMUy7N3ucj7h4j7gUZ7QRCwILH75Sl3KVIPLw6xEU+KVzcnqTWoPUZyblOTSN2lJnulkeULkp/
5dLUACHwr/1tQexRNF2tf+9tEX1UJHX0Fm4F90VuTcfl/GQLeC2/9sw6c0/8uOTAsFJso531nlsE
u5QF1b1dx2PE5UMlq0M0/o+9G06AhthASAeGJ6mrVkdtmKLwWLE2B2lVZEqJM001JMuso/MXWuaw
rJilo1Sp0TlHs9savCT30lzaPw+/s6IleEULrO5N+WETb/ieAK+r0M0WcdQQpFicZ2oAMhMDBAnw
EkyUTTJ6ym6iqgnfuQJfHEIZSIaTTKwzQvwvYyRp78FNOZhLS3w6C7iPoIO6M+M/bulMnxo4j/tO
WmALgvIGOT4hB1B80+MKDq6M4FWRf8nN+FoaLPlGOlSwi5diBD4lfg7mPhTKK5dd9kWjGNnF2Y9l
ZhqOgY+fa0CtZYW26yea4nByHoi8qVNre1Mxpl9wU/05gjxnh3sggHnQYENgSBPxn5DiVoLkX8Yg
zBTbuBX3G7EHKoba7ct7DdJpmV3ii8v1sQFWOhSyRPIBRKbD3Fe7fo/+0meKpWggxFBZkm8KtnBs
/yB3IUbIPhX235s7U3SeLWxr49QEAhZz40/cIfKLP5cqSecL0d1ftl/FkKxU79igSD+m1kCSSk29
1pX1Z1T0QZDzxA4ik/tYWv2qdAxietm6RUJ+kqRkCqKjLYW/yIPKwZ9xvbgSu2Vqlt2S9VkJ/7rQ
o1aYTo42Sq1LHmKA3da3z5L91hPtZ4ogjKNgMNCzB5Y+MvL0x+lz70HIXfAIqZQ8kanafEOWCaQ6
QdMf/nGGLSb47yFPuadjOhl4AXWM9u4hzfzJO2jNEBXNCfngdpQZW0KWPrtmziuL5xqczQz3v6SP
PyT6VT5HxlP/S69n8CZmyc8AAdrHMdXzAgNgzMoFkZJ38plrMfPafEJ3ZxLBXRRrT4ZuLc+BZOrK
ahIUTa9wJ2IW8hlZE01iXXR55jiKHh96A21xPzMHOZWUGvsDeSAlyZzfkhqASDTCEt6/SVzd2EEX
dMTrj08W37mLSeFnZiCSGprKSi2vW+8STTQWxWtluwJZDJiqG9XAQ5xGktuwfq8daSFGa3lmoCPj
4r4hFLELIKJZYPfpxMPAtAjNBv8CtyGSlv15XdID/e7WCd/yGqPVfkpzJum1rbvvw4dlqQVDlbbp
YHS/Hwe0C5yCuoyu3H2yx+IOn68dPZ7wQRv827dtloxYirM3RnvQ2gMIfXmN789TGS+1h0H2zDm2
a5YyRND3NrSNdt8lRxNJlGCp+TgP2JkiI7uxw+weNbv/wZveHrbgRPtaFf2xw18UPkSBW14+6TOb
/WwjDjKD680lCHDUlpAGukO730FwYYaCocDFyLWQ9zApaucUSfuiO91YEvgrSLzeWcjK4ihIkhSD
9FDFhlCBikUw3zySQxre/kKY+8JG3gQ/jWl3C/9P27LjMzzQPhOCL6ua5m0JpOLGEdQjTUymmWCJ
V7cbL6JkntQCMv5OEVqJxiwEyl9PGM4F3DwVMtkZxAY0Gr/kyYmbbCSLrPaHOb0OSL9+vPko7Wvi
gWXWys5zelqiy8auoWO60tmHrauAQENqExPZ3CdCKPXMrJ8YMbcbBAkCq04vuDErxRtwTK+wTrLU
rCWellte9FHuNP/6lZH5wxIOELhgeglsG6rmKeigOLc22cV/SOQaH0xx8fQipFIQmSvjItJmCWGD
p/+SpxRgPjddKFd8Az4UcjjMY1mMX9+rTxAfhfjFyJHcQIHr6Fn+h0DRuyWpUAU+B2MqLYUBXuKV
HcR9thDY6abwYx5CVbCDHj3HR3t5Ve18uVUZCKZhbpzVuVknStVSk21rzFtw5e2WFVOnYMg6x0hr
NTr92yAjb8z9dT0th+oHsEhygeo2F9PDZ6LeJjaMLf7SvZgigFEpqc2OgNqGVWuPHF+4ab0LeDlU
3HXlLxAjrsZXLTM8i240f05teZK6DfBmM7c5I7EkmsLFAu2gxc7tZtLXEkNFcihVKe1NaWeQPiel
UlNpAEwH7cnvpe5m8vzmLXgmCcKEu273B2nLvtmoqhwDIcKo2PT1silhXKNOc1nE+K2ARZopOGQl
d70z7o+kFkjdvgGnaXbWGwl2iJgRNNMwZQ/4rLDbUXaJo76pMJLY8eBDfK2ZNXveYsN/DcuH0oSM
luGNKUZOZWRaxLdQpge9zne1cHGe8W3LPmAS/CY68ACR58bern2fUP1kQTsQHS5iWy9dVdn+efIo
8W2FCjh5gPzyvo/QJHdsOgzxX/gedUWvelFr+KmCf2tTVaaRbal4xF5mnzjaXO+DIKABBv4g7FwM
+WKlzrRpacYYBEel6017ecy4BF5VJw3jpbW38DlL1oTeTDwOiPXyUHqxuke5CHpGfZ9XmjYzfu3o
MyW/1f1RAj/sK86rG9aVBG2q2bDsYIcXBk0L6X4zjhKVjcC4IPODfzOwAO1YkJ9VY0xjWsKeYfYJ
2NQpU3/05RvE6lkCTJUEJ7J9SEuCCRACJWh2aynuj9Dae2YotoLW3eIku60qJtvtKICkHAr5Q2Mw
dee44CFPF85tCebjeloS0d16e5fgOEcAsu/U011KhzwgPEC1V9wrOX0i0EChlIan4i9ivz4SSGcj
kejtfTHzW4UdlTGBDoYJwnDRVdS18Ig9PJcMYj3F+BrKJ0U/Z/shIb9UZhe/k7fTobQRk8XCZeup
a0X2Giae8R1jsXm4pzlm469J8bvwsm2QbNqygFMlGlRVmg2H/YPXKW8jpGLsYZ6t+plUCaYJfBcG
TDl0fc9z0zOfhkjfDThs1vgRShOQ3lhmrOhRnxUJLZ7AyR/uAuntf2l8jzIPZvPrWI7pLAKxF7OL
lBMPPtPl7cmWqPaHuLAPFMOOhCan9Kw9ylCdZleObnXJcrCxlqyudp94dJRGuxs81zhemK/Y1fa/
ZCsR2Jx8EpnARM3j5eqT0evC/AI8nSpBAKG9YHrVQ8wO9KaV2NMuswYdNwa8UbxB/fAZqnWoXq06
jxvXntBM8c23B9avnnKEQ1MnpyuqxazRNLIJUAVwatQiBKOC4S2bksbQSOfSNHkVD1OBSU0vdQuV
NXVoAzJD/Tia80blxksfgOFDUD4LFeEh9PXebsMXjXnu9fQ1MWwmkhNkiDOxqw8AEOKUteXjnSsj
Q3jX3LtsF1Sg07zgDUGlPV5Vj01TbFJQFiYZqLNLKInfiu96jgMx3AGVzxUGIUQWfZUmW3lDyYng
4PyNwkl0zXF33okscOs+8BeLr6IxvZtYwxJExzQKJlL/yAy/g7nn21Kg8v5DmCWCIYmMO0BMGEaO
qOYNhVKoqN95uF9CLuc9W25KEpMKu0ByphsbxuN3qYr4qA7XeSJr48ekj/8ZngwaAftWmMNMdaGj
03DL2Q8uODetxMJ2nEaaMiz/9muml//ei1M9/X/w0QxSx9/4v7lg487mME97f2gaNsv1ySmb6XQj
Z/kqF8p8yR+bKuk43XnURZuMJT/E8vDu2MVBQ4tg5sCCgNTyrbDeRXXMXA9SeiMMSKnU8ugY/qfh
gXHza7EIMlw5ReikihuzUPUh9b4f9ZdkcVsh6BwTXQ4FYgwAIFNDLhbiCeA2OWZaHiVHmeie/Cky
vaW5Qb1J3mCO/sGVmsexiaP/pFqBOFTMFgPOR8f6c3A64PTb1O/NMFSBKiKsEacQwhza/5IhFoad
Zn8NdpYp+FFqUuJSVOIX0IQzGozXoevenX7kZjMFioZ5Kd6yE8oLPscX4isqJspC90+3DdjuGk+y
4RIJJmLey+q1DK1xBU9Ds8siyNcrOdmrnXIlgwqGny0Zk2cPaWGHI3ARr/PvFSNpmHv5jMmkHMZk
H50rbaiQibI8l2uHEsOjHb9whf/qAVduZuAYh67G25G1eeaOY9vXuOvIe7AiZgnuvQkeevoatKMB
QhzhOk8+gIx7914IcKWAcpMhrlm9kAGfQ2/aAI18dWFDrPbhxh2qoiooKSDMSlbvAxs7r6Gyuvjb
0L60H8enCRF6rnkId1FKYTKyqGZcYEzYOy6W1oujyNOyVzKYaS+bnfOqlDVlOyVRW9lUBXKh5ZVZ
q7XjjIGbMoTqU6GoYLojkSCAL/sXhTP3IT99mJb+HwDCxs/frhKTdffDULqojYai4uw544XaOZQ5
wfxkEl9eYMp1xfRy+772us08/xquw2qOjgKXMo9B+ufseR4iCwp9cMx4F4O1BDCEmZKlMfxGmp0m
F9J52X9czu0vo/spcO4/c0Edv1xfCOySUOhtSBWhmJ+2b0D/odcGtf+qjGPDcEV7NKZfZRT3XrIS
i4DtICwa5VJ/Ukxzzq4FXrU8f6CpDsRDBqKVp5vozGAi6aSUjkgIu/UdfaVqCkhFsBXUxx56Lnrp
GizNgH96WwiyxHxfJFYabGP0Hd6lONbwc2nBMxrSLLH9zbp/t5qjz6lwM31DkgOrlYH1AcsSQ5g/
f7DuO85s/eov22pa7y7bvcou/AvECCyI/jJt2n51zYQu9tqjWiEwMC546byDaFgurXpnfoJiGRG/
rC+yXvHa6/OBJQkcdinrYd1VAL69jqTQM6XydiWwsmO4jG9xqLtq/xQy6MB5n9DyUOv2xj6nkTyt
sAqgZpMgi5JitQc8tJaq0K3CXgylKLgsyxJnAbNJS1qmzbl3J+TytB5knaYxLuhuxnSy/l8JAYx3
XcYYa1PAfUI8xMid+HbsD0YDEyoifwAxbfvdE/b9xkQcMvoIZHWp8VyfW8OJmtOO9hqeEfiGhHMq
eAJoQuzG2jv7+yMmiWax7viIN818OAXmbzy1N0HnLaf4k48+AtO5Up07Plwl26kGuWPxsZYUpC88
GPndvered4Dng4C26PSo1ISvTtCVeHvD2vduwCapQAoQE9T3McuUCn/gG1eRCGU5ozfrYQMRKg6F
fLIgIVVABhRtxm6L0UESa88kA5TEkJ3XBBnN6qb2lzKYaKiHFgFePyC7vYqHd6wk8150duU+7kef
hVHi/0w8ebqR7skwPQjIlpgIrU28c/0pLco15QU+kx+VYKhutRgLj5il4Ot2LmNqCV5eamXukX4t
T0M8dQJpO2LVpnKzq5/vcJRo7ArMJYQb7Aa8tJ2VRkgJTYgL6im38SvRHSYDYqpSDi4QExBtayhA
M24qKrB4LIm7AhrmjZ8WfEstiUVDSZHgn3/V+ED5fswGcRuheRIbC4mxol7wbtcYeti9T0DRxkTy
Wl3pCJSMNSYcuodF6kbI35W4eHGdphKWcDIWn8sqmjbOa5DYg3V2X+txihkFPgRL9llnRZIZ/1UG
kn0uO/wpIRdY5FkvD0v1haPny3x+cFalntINIAWrFxySQ+ZQNFvKfayzZfSXvCHEKE3RDBiS8Oy2
s4AxiIexFNjCx3TUoS++/P20HS0ZpGbD9l724daTXIhcW15PJKA+B+F+l3+RLHJYTwPsHtp4910t
ohB5+4v6pKFrZLOUTBEtaOati14nHDmnhcvFS34BZ+J15ipCIq3cVO1gcPHcOxHIFdvis3c3YXoq
ydxaxsc+9X6oQsj1bqSQZmFyL1+trRV02mplo94cigykePdXhWSCMl30LjVBFZn60w3Ex/pQM3E6
kLibc+7Yr9PnuWN+6dWtOnq5StOL78c+TrAz2JIgRSSPXCjTW6+S3XcnxOyvh/Z9s15hhjpHbY+n
Osn6F0GyBnsUMtHfqzETr/rJuvCZJEyDp63axLVPNJnAbYGEnUEa2ZNhYTniOZyX5hQtYNko4/iG
6M4Wda5lJXoyWv65rlyS6nfKt3/FC7PA3VOIvoI2Q2p6SaS9uEC7w1gKSHRluV62ABkck/jgSxqJ
DU70U4I467SKVdlcdarcS8wujAA2JRW2H1xWFYcaPsgS+1rMouip3c1ZWQvantPS3r7je7m10FT7
nstKHA5U+w==
`pragma protect end_protected
