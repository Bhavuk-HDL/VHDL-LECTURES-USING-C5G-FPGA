// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:39:06 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ZaNf5BWxDGaJso72qIXUHFmTbYn250q+uQ2C7jaMZj6S/RO89h77pqEVDTyTifw1
SV85mYgpK6Bu8D+/gs4L7DiTudXxEnkIhmPya26sg4g9xk/XQPrDsk5P+hMdim8O
2lNSmDIVGFFs3GZqtHzVGClVR3IZclbpVG1ogI8OyRY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 184992)
M3yvwR/je4RV5kE1ukwkZ3vg5WWwXY9hxeem2qY5zZ1hgK0gdNhPIs8NmdjamXzK
3+GdX+YG0rmWQFwrxhSV2H68yotjjjrc6mLdCMD24ck0drfwObYSjYVIcx/KkEyN
GFBn9gUCvA9p96cKjjSecH9T3FMJUWmhVhhjLIUEpARyfm0r6UPBimS/ti2yOtBb
JJjfa9Q3HjdSAwJBdNKcOWieBGHnHg3NV0Hagy02AjMWZa9aye7oP27mCSaakeik
j2Hv4x9UfJ4W5KyrfK8dRrj034G+jijuqUS4aGXRFmB/sNzfaSVkQcbWtRc86cyn
yPww0Xl7899uHpL1h+h58rUXHi+FyK7Y9mbbaX6yOI3cRztKAVD669m2yjGKn5gB
3LZLqxCNJx7ILWJxTFB7+L5fNM+YG3PMeavcQqm461qECthO9Hi28KYoYXKTsB4C
ObiKl2a2AJfiGMUG/qE63HceRn/FCiMTuSMCav1QmP2431LKSC9QPD4UgsBalPI+
L04TW4czy58pLnVWx9+VIvspaMZcdpuNSdgfT0jyODlfTY5N3lUHsFAt6zh30kWc
QVuFUXsMLBBZomEQYtSbJxw3GZUlk/mm2qIKMz4NvvOUCynshnUyBXHZ8pBqzZPN
6CLguX77Uc0Foalnre+5PbU9FQ42N3IJwwXjX2ULF8+8d/dC1gEcEsGYZrb9TlvR
uHB0bUFKrZfv0g/zmMJHxMhg8lZzAGKfbR0Exw4Hp6g73uYpgupP2Q5hjE9ISPbf
KGd/biTnjf7Z/gWfMvgwsPm3gmeCW3WICEGcIlgFgOZ4naOL+f5A8ayCCe8i0d7h
xHIZrcBPl0/q3trJUEz66YIEjX607saQK12VUtfX0u325v8Vtjb7Qw5V0ymt8d/Y
aVqrVa1DLKUJnt8a9D4aVoMI1zj3eV32NAz6kHJ3/lo66bM0+x6/zQ9magJ4F1ER
QNBzU9ARiLfbgZYFLdPcVL2YIKPIjnLUpthyN9yv8T4JjHVCV5nL8pai6IYZujaU
zbUsE8FFjcW/h0nl126/A3AcZDtcsWUm9f9rmYNIDQYd922D8AkqWnz1Vil0Xynb
YY6dYw2/XrpqjCLItJaztIPZnMXPLSAWBuKXHhJI5OXTUbm9ZSt/Q5DfHB2v3vws
W+wdAMjKY2SyIaZDT9Yi65Gzc7iFZV8ZcSMMlFZnkoDP0ea8Fj3rc37gQJZcBgIE
bNXGoDyPn98g9LzFVRGocsxRif6b7n2BNqGWa0jbeP5OA2I67itLPh9WscfX/rfY
4+7JCdwCDrMScKQVBIyyCUpnWjNtwds697Ce+iYi2nT9MviyljiKuX9mJqEDP25j
ZAJ1Q+rFpmxJNzjYEpKIhZy+sg1wxWclZT/1A4oZ25EhNGmeZwv9j875z4Gb1qOa
hJrtIJHTstBmfteXsdwSembgRu0vTOc8M/JNatSMCad6NPro8yEFI1ed4t/gAA2b
GJ9GzSz2oUkiC8J8Y2Dn07niNlq/V3GQP4/ey3ND1JV69R4/UAWmCUv2+Cn62AX+
U3mAVaRXi+1XFwJyOt9TxfPPM1Cw26vvOw2rm4S2v0uzFQvQWuuKyrdMeTuvcD8N
Q7XdVaO7psPlWlz9nYWJFFcddyQK4M2rhCjN6Oi0Lb9ZbFRvvbJ9NBjVvKgsrZ67
qkl6TnfkZcMNcKV7M9bHsKY1oGSl3tlSwiNWNB6/ACnvZZglohui2w0ZH+fdHOFi
eLWMBI8tD4ZuivqSHFnhERZ+SRCEaLxbs092zHKH7r+FAI9dprjhiRiKup/9/Bmz
hjK5zZQfvmw8A+iJ34sMM1Tv/tCfmHzH0N13Nc7JI0G90ckt7gYf5bxZMIFPBi1D
Gov7h6zDmMhWrwcf2hIZdRKt4X8WdI44F3wVjKHyKHOoqVMMvovd0zrT1OlZNnsQ
qtrXC9GQ5HFMeMjQDijkZLPltmkhXVmeKrcqzoy1lJ4l7KXeeO/T974CyOLZvp5N
YfdqirxiG/ideOwJPSYCVdg9J3NuCsoXvZMLVFQyhDz5LrstC6jjZR/WzZgTSFFt
P7izeDbekRf0h2uZ8vdOP4CUd9zcGmLXvgxYFxImMLDxtaSlWPSlfQSM7AEeghYi
tEINhYGliUPpmdgwK2WNkx8lydMBjHTiL49YQGEiX+Az+xhxAgTrgCj5T0+H22mW
8Fq5el3FRU1V+3uAkIFDRt4Xq7Rbh4Xx1uaaPbLvUxHhjmB4l4sruYFHm8D3k/TL
6y7lsZpWmSSZJ80Quu6MoKeuTHO0z44j/iTtFrf+dbs/ErintAJCY4AWXvGXhQTL
YKwlRujh/htO7tebiN01CcMwogunNJVwYjRZJa+KnVwe+tSyl1rYeAsdlA/DhDIA
s6FBkBFZM2QEkezRP/1Mfwa4uy5zjuXZba3ecQJOgW3daJ7aEint6HOU0OvMK+m3
CF/ImsOxrquYc18+6LD48F+gw2AhKDmELEGO1MUDRT7GKZifRr47jUrN9RdRilVR
0e8uucl3zqUuNmFPPwdOEn1jJxZMPEOP/i5dXReZcvWDlaJ/k2f54J6i9I0IxSnm
HD4XadyWkGI1uJrVoKqsTS/AQoM86XKsBkaMF13qKK3+yLhgMvzkckVEX/YO/fMe
9KRnh8a3VQR6vp+WHTkx1QmW8wqAZ3qmGsO+YEgr+ijZMBgEZzEopVzOjK6Cjs8P
GblH2D1OlJMpR6V3qCC42k0cZ9SZzNxTg4ciZm6By+xOCO0GOejo0UmS4MQ27XMS
H/zpGJb7v+XTk5MtIHDAfH5+m1o57wfAtUJ6UuC0Kzv4vW5HO8Jp94rCJr8xvI1h
XOFn+8ae/36H3wYIBFZ317beiNQLxj0SMfMfaXL7siS34boZeRhlA8ThiqbZujhR
34U1RSxDcneShSncb9tZ0N/GiIBAZIUi2DoWkylmgoQKG/715J6/SdsODWSH+s+T
9n2iEYR+5YyV4CPlzY7zIeDdrbbK6fV6KZiBtciuggUvWtHcj2ozmUH+19ZPqqPk
VnHmnX2CwlpEgV71TM1FqIFcpU8z5kbl/wMz60dECdF5RKhgv6Tugyl1VyNSoGwU
yLnPllVVVP48S6aMtQ8VeI6XVoyIIV2eJ4ypsS4Ri428RpLDjsQXcCTr45KO4xwA
3vCQy83Y9kCknbpRi4r/vE7NwYcbipSVgQAAnx8fcYLb+e9iSm/JJnC6uVHjw/B+
Z0LDRDDzACSnSQA0a5kKhdaAkT1VQCEcGylYBVnP/LZmfIX4xGbsqcqVk7i5rKWO
NIIbnaqUNeGJiJk1iENraosbucPnJ78P5+vF0utX/bW6ENKSRHnU1LxrdBAzJb//
NYzB3mhEoHlqrbSrN1hknXx164vHNySsTehlmIgE0BlSEmfBLuRvBbuNmtryWIpi
0QPNMCtmQLFmqDr6ZprH9SD7LStg3yhYYKPbX0SPZCkFxDUt4iqa813dDF51WEEx
mv/2ZM9AJLfNYD7CKL/SnJduA9qn1jMU+cG3JgUyVxGoBuphRI5swCJk/AxysjFF
SWAKL/UFF7jujsZR38eYB9G27EDXxKqEwv3ReezkM1TTsz/hDxjfRxuj+ghJwRsM
3HHUQ4BZjt56C6UDU+hj2GITvCUqEdZgicwTFk9jt80uJftvx76BesJDgfSeFiUd
H6Xyn/9r3fczfdvSiVO1hyPEo+ZrZij0u+7jWbp0O51Kxpwzr6e3hg0vRl559Amo
fd/w3tknzvWqv1WMYLOsh/hJyUAbii6b6LSNwaBsNr1/MRxadlXLfq+qLiq/U+wE
9DTwEVNCsCWJPV2cIviCX9n6DeQVBdBcqqne9zOiQEN31at1ut+F8IlnmvvBussb
Dp7Let3wUZ9T2Oo0s8mTxJu5LMmQrLPgw2gibq0fMc/883PNJbOOfC2s6kr6FzJx
EfjEOtipc6llGFlOecxH8UoOXScVI3Xjx9Kz+oR4AGBToFV1Jrfu4Gffs5tCuG9g
ir5XmEBGN5sq5TJMn01pYmdT+W62n+73TN1cWBRT9cEuoeYBmOn2ui3qvxmzHTYB
EOcpnbW+yZ+o1WD2STrbalhNvPU5S7sFlJpwgWIjZ5koBd/x1rfpSxYrelsELmLN
8gghjHgJ4IT9HZJ+YqSbmNGaKfPHIWv4eYwDZhvvR7B00Tpvqt5o3sShtueGWb83
r2k8JIsWfzhP0Z0uooRi6TJS70cswHUOVM7cjlYZZU7ZkKwsrJyiGMyLD0K5p8Lg
ZEhSgJ08hZFWP8FooZ26XozvSaj1vwx/cBk24wjV4ro5pTni6gBGgg2ZOTN/CcSz
SjHWcPUlXD9j/YsmIc9M47TMbwycC0verowj+DR5Zsgf57F7uZgKyah2zhuV1VmU
ezz0fyoboSKopTO21tssEIvfh00GkcqDmgl2ORJ7d+nklvKJfu9O/bf2WWS6lVMV
laj9Vk311wED5iec8VQs8f+d0ftUQWkLs4yd0rdQanKK8dGLbooA25mEyYJPlIub
83Rwif/zNAKS8Uj7JeCLEMXfKNsxIPeIXUZ/3VtO0vKZ0DXeSw4jmbpYJoGbYthL
pzVl/gEj7rVzTpqe9g+h2TC4nbsWE03Xj0FB99zK/P5BTffuzpHLyyhG8i/tTMYh
gQ1cSmd7QJ1Xqr5ecjHlPQReWB59AWQS5aKXtrVGRvDill40e/9ASUy82pro9c7c
LziFyADGck9pvSuqJ6mrC2qexqHnLCZ3vzfr2ZfpTicXcbgF3vZ4iHcryqLXHPUu
uPHA4uONt81gS0us1MW9yE/2U5aMk8W5JmiSIVDGptng8H2fZ9sqCOOeheyknMn5
+z0qSVy6A7WdFcKo1us36VKprKftxBHMzH53b5XTSUzjpafFk+euFDQ6/tURCXSF
YaRxF48CEgsbhm6fMAadkvhhZG+3tUb3hjU3r0DG9Ihjy4QkksAlmBO56XHEIxZa
byrTmjcNiW9zJIBI4e5Zz/h4qzyaUpepax5muaByvkJUqcrzsuS0S051pztR58lo
dZaaPrp5T2y7s8CD1H5UGC8oUjGo8G0IRRuMcYZMVMsKgCD4itciUQqO5oDyOWw+
7HKYVMBZAFulNvWBWkeCOm9GwmdFlqo1bzNc8/BdXK1fNCpn7INUNGPdG8jrbdyQ
G+99WymJT89ivO55zIq3Gf9/RkC/tiVrdh7tAEbDFnHuQx7ilTucLtZysJRJNdhs
sJppMxb0kEc1nmIDqcELQNDmlGugO7UQ7v57sVPRizlttsNLBZKXgoDfFFWIZmu9
soGYy3ybBbSNKAHsYxVdCYLg5PIxPaYIgxf9erZ7rR+z5LhZGZYAKmoI6p3n3Uq+
8DCusuFb129Ns1PkTZIicU4rcUzrKOSd5KrsBKreEMrKfzbl4bmdx9cR56v1lZdN
1EU+1S1v1DdI62jeZyR31CZP3QP41S7zZRucz7JJyLTutXowuLcXsvDoPhJWh8ra
nY8PC5pyRXVXtCHfuwzuvxR2YQG1tMRq6fkt84BOHGoCnM3ueGxX4NomFTecb7gN
eiTxdlCPrpKeFHtzYvkZWtQKOCWOtyZzW0PSNb3O+zHDv1l/c4ERTC9UH3Vvurmh
1Puo25ghYiLqtphSjV0Cg1H062qN9z3aWpSHd4SENXU8LwkVuOS/yi+2Z/Ttacph
Azn4lYhH6JJUbNTZ5NNswxAK2RQOmyYfA7DBHmwBpwM438Z5TUdOVdOI2vdH7cmb
ARJVUxxOfIMIAnV6gND0dBC/O9Yp8b3Jh+ieHmVM5IBsNyBRZvncqTgaQWssgtNq
mee31Ub1eArWlazKJtwMbyL5ju+DyGjk4H85diH6821TLxWhoHBv98GRAfx2Isfb
oqEpuUrhz1ONjALtCJVGTBqHuKfGn9QXWGDcnzxZY9tKWnJ6JaDhMsUteKBh/89Z
qAZOBVwPY7HIWINxdy6l80tEPACS8NjTlSPTzvxH32gTWOqSxprM7Qq841race/z
LKFHG1depHmvzUs1Dr2NKlm49HKon2lwu0zQYSMiwkK3kzszZCmYG95MyV0EBHkG
07FcfkHYWfmIFBhaZN5jCLuQUh7kE3Li/vLJ+lD4anoC6yEImMLYuc/hubgGwJmK
L30Lweq7zhVRSsmECiKz38FwsygXemoBrhW1Rj9XSTVqc99Kjo6Vo9xID4xuLvUT
/iA/Fz0CTfJ3ZYMPFNFmTfN8Pdn8k75y6QIZwITzCs+YZflKZn7VFVfO6XNiYwXx
f5D4vn29rr7YTAg8Ce/Ki+pT+pNomxJfel/04kyyaQ/PPWQ9JqZj3+cPu1y29HwB
qgn8ZsE0Gn/Z6R0n29n8pAZewWfM/bnjS2ZiTAQ4UbcVUKcHXNDjL4eY6gQTEL+m
gcTFiCiIaqmAlq4Hi9nkKF+WLNxfFYp6p1orj3ju6ubL2cBkk8HM8wq3Dc1XWZMI
2s8B4VLWfHvQZqjdkKwqHfI/huLviLJuOzGYYQdLngdVW6IM1At9wMrEVSlqX6Dr
WMyAhCXVjY/bN3n40z6nDA8EQETC/PVCqqDueU7pambnrOSW3EinYVm2Uz5TdYn0
+r/pNwvYJz/Xc6fWK0PL7+V9iZWq7/rwJrVdrka17h8TbhTNZ/0dsZYoglEqMPJf
bYCSrbFWgWofK73Slv/WSqzk4XK3jprY0pptIMb3zApdb8LrgDgNUD8J8O5efNXN
7+2j5vr41br7WldFLo6ETW0aOD9JbIvOSJXv3vmlYxYvrrbS5gsx5nALmPtWY2hc
Vwj7GnCuK6YyNWh3LJPfrW/ATfcgMaoJLQRsS7ORZod61qUEdaQps0jfTxKJIMSc
7fcZTb+n9HZyHWo5fJ9mLqppCPlUCNGzrdXer11w5N4Rl7Nc1+2p/U/Sd23ZSMOc
E/gYjjI25ZiH9ULbOZOr+FRW1u0IL6VDjQqHX/B+eRVGSylaCeja22S/N2yP+mzm
77uSGcuBY/xT3MUkgHRuOlryPNjO0uYLJPC3JVEZiPgtrLqjH/8tDFGmiMNH5dd9
Uk0yUswywWdm6cbuah7pqIeQh+S6eMvBHCTZ2tViu1jFHhGEfDhQzwQ35+2ohAzK
xnZ2NtAPDX1ku1qydqHk5lUR2MzQ55ztddRbfdY2MMH64CNj9UDrX5ijEheQAUlY
xlbo9AFjjdb5eRqHkC1sGHGIxsK40gnam/y6CKwaw1JsLJajll1jA/YRpowFo9nx
AZXwY/vqJzNrjgStnM1P8ui+WCpf4ua/3zQynqhf2AVp3UjrhFh6yguCKUBLF8Ga
qN9QM7smYt+KYKApBUlaW0v5lRUU/rBpUVdYDHOER5aCl6+1bAtGlCuLt2hun7NW
K1fWdWB8ZTBqQhROis0txfqcO0daLEl01An5670iguE4e89ALUPjjXHPF5/mtleC
TtdC54vGvq3wVYNr3jWi8Mag4PNUexYlMi0Sk1XK3SaZk1vdtNyc2+uh25MQRgpH
6ninAZ8ewTYxjvsV3sXaFMVRMa65w6w8ezHs2ZhtHJQa80p5JH1/0gdYzUMfv5W9
zob4NnTxi9mrNKx3VUjqxqVu67hTVj6r6NPHH+9MAlSo8hcT2KEqFNMxB9+qlasa
+Id6WoHBjegLVtuO4eNj/Jvpabe20f7Nim+I0Tk1dT+rzsYxM0/CabRjJefxg2CT
xQK3cYav8F/3cuAMyc1pWZHLiUsGtzGm5uHe8x3LwL7B4KXhZfR+5jL5C7/dg0YP
qd1o1Svkp/znw852+TknfGNS5WfuInki8Z4dZ0ATC0THnpQJ/ZXSZDJ5dHZtQjq3
Ox8e6PuPDxLYzRmILV7YAQRHBqKdyMv1Nc493bqE0HXsSXxpdHjL9W0VCQb0dQpF
kQKgqJB1nlteM4H71e2vRGFdULHG2dZt8ug5auCeOTCwHQ76Epkfc044gLVdkz/l
+iZeKiX/vgMrWCPcs3KeNo6F8wxG0a9eTdBq2hF3vH1hY841BHZ/DYVfP9IyXR1v
XoqZFTZQ3zZ5/Ru/kvnhBJo54dsr6FxAvg/O9Zt4EjPJr499J3DfOgnX00TnzEvN
fdkFF9IbARPtxD5s+XR6vrfZoJmDTT7r47pO+RMcm4NL4pk561dFKNFle0k3nC9z
kLLutNFhBpq2qgX5mSAxf+yk8NWjNfU4FEFgz5K0i0+5o21N9wIU+JnfBrDzeCSO
eR7oDofPh8k35+Yo4azuQR5pjkrUySy2tc4UTBmO6G2RlDxy6idEfkKMtLYyhRhi
L6AK7tHMuxdpzOBCf15knlUOv9ffwXF7kouiPMHTfHl0vYoRHHieaymTwg+wDQ4x
okiEJ5Sax56mOX+OD59yGsUYd62VO4bKJvCEdcjkNJQ3ifrFm9qAI8hTms4KxYrd
7sjwkKbVi/KvZ/57elPXKzb3qhWtT+tvWXwyr/D17s27hOdElkmKsxH7bcgvdmz1
GunbgHqooh7GzXPSml//6GLmar5xLQYnbwMTrsjk3YjmAZMBPqGaikmtMjKNAp+p
RYHpOXkKR0jX3lRiBmneK6Xb475+AWhsIn4PN/Ly5RQiZu+8PWXJFg2hMpzMr8ks
5ToCYvmetyA4Pa4M6lBjHtgTGMpGFa5jKqRlgg503q2JLIl20RnRc+K6HlSJR9fd
wIJg2POiptQXmkn/9jUql4sGUFZqI6etZwfVJISABrmibRnIGaV8+8RR7JBK5bLh
Z/uekNhUnrvo6hF22UYD8ur8+xC/vaGzbfvi3iM5PJ2++Wd+i66rUuYUq1CC3swC
RtrAeFzqcbS+7Xwhq/etP45QxpNpwGbPHvy4D7PXTWolMZmcROx0VO5Pz8BmUJWg
z6PrcdAZSl56pQHdXfVl0gI9j9QwIat6G42btIsF+2QqcSv+KHp4tc795zxDQ73+
8U2SBdhqCNyKCc6NJ91K37d90J2SdT4RNDJ03srfR/j2yQYxlU15EnI/rzHLgy7b
LyGdG5VBWtkzXs1EWJyDicdAuhe6LqgA+4B+im6AV7WFe5vcWKm9wHREg/AGnFNq
nWxUXzrKgTzz4FmewkhzKsJqBCxJgyOMOX8Uw7blR90mEaiwRKm0wrFzDuHXZQL7
6EKsWTLACjj2v2u3wvD8KGtf6XLDedKFFs3dYVeNEQCtP6oOs2iwZDb6J6ZilW41
JezeK7Ve921CCbcBXK7ng7G8QRDVwp3jkd3I4gYF7IPJbVbhq0Oin0zudcLNjEvq
D+cer/DQnLfl55G9LMwJEktNd+wnjMOo01kvWfHMca0uWqCMObXfELmSsbEjoS6y
djYccOej7CCiZD8PFeTLdc7+PgwlYNp2OW13az9dDhZhJE9IaaS+RD7r9svxWxHJ
fgx2vyyl4UHu1g7lmpjsgty6aYImICGV+tyQbSeI75JOBe9KocE6VrPynum+FhDb
DKVYDE0vUbuPJqh0sprV5fRP5eQvA+KQGg09w3b6Io+5SZQLZ4BPcFZeJAOd9m5l
fC88rZ+QwB4IJoROx5kAzMpVJF6OGJDh4/s9Ku0GM7Y+bwlJ90YlagsSu3kPCYw8
a8h+MAPJn7UJyto80pk8vrVGg73X7/ST1t0vY8PVqC/sVsbd/qTU96ksUtM6koWn
8bb0yjt0q8QRBlCnNULpbUy22s+6p7ti2QMHNkyZdPJVfE36JlB5b/cPeABVYtMT
nc7nl4kKp0z0y+4S+hTblEDg8XbK3lsCT8UYon4KFbmZn5QIA6uuHgNFE1UFfXSn
IMYr3kMbEKQOH/WeU8zeuY5cbKlt6y+2GoNJQ8spVcyz7gvyjmVSm3cLF3NO1yIS
bCTULwufyo3Tu+Ns+rsoE13tUbuKU4d0QggwclAK55AZ23gkQ5Mm0PbCfsCD7bge
xzOO1dboeyYSuQRG4BCjF+a4OWi1G139rpA2tMQq49sih9jwSPB2L3Aetgl0s2Nh
5ZDo3QEVxHaWV1NLCja4A1978W6nVTw1HpFSyFrktTNzzA/O9gtNRd0P7xkPnBwn
aOCtl7wk5i+PA5yOyzpFnn0PIjnD41ZxxOqIReZHrbHGPCqELrxuln5pJHlEbN/T
t6nWUf3NoxJwAPrlhzhD8zjDXZ4H7Wv2Mlg4l+AjqzcMpWwzzfhV5xuOaEm7g9gn
0sj6KtbJO4Qc0B8C9r+r502MG1DDZ2sGlDtLd3ifCdh+8Pb0lKNwbQtgfkRzG4HO
UjRRaUJoqCTbiANTa4mSNSQPcAXdXjYarlo7/2MOWadDzZiPpLrkXyRIUszTpz++
Dx0u/sAj9p37LVLsKIwpfZTMLTvVbS0piYYpdUFP/+sX5P2/fFqzN5LMDqqdPtsN
CDcmgxxNqCuajnWzK/RAALBKfRP/JHtfHkUrNkNGybDdk9cCX9SI5XtZTsWGdaNW
NLagvfHdMA+2Q+k7L7+ownBMohTu08L5QjohMa9UCtvqBQ7Jh052V7QT1Zg6+So4
ggLdJQN93rueLkB+Dh5C/8Swg6PjIXCFBCDZAPyKwt9xz11rfnhaNZtihD0byj2F
kATnkLK0spycKYXb8xCzSAmmMqCAlBTsFjGcsQtOHHrg/gcvj98F8nlq8xJXYkzj
lzU7oDjgYeoxguOtp7xnR+KfHhpEF+MPfyXZjgQjIO+nNVMfIRVjmdoY75uTAYlt
muUYe6OIeeAZ+DEW18EjbOftSUyAE2GW9c2JEcoD82p2Yqbc5snP0kZJ9B7XRTVk
z/YMGwagErXjizlpJauyAg95Eu/kpo50QuJfoJ42z3OrN1ullKfxx8i+PEN6r+Zh
cE/wbjbn04+uTrZw4Xr2X+qlDkRHjkzy4enUxb1OciiEPdU3KxOUNKysO5I0VXGd
vq3/vLog1dBVo3ojuDhZYnEXWvUpQB1ssl3/qZdQvJqCbqFljS1zUD2XW9YXERzG
4iNzXaH1cRqEtk5GvxxGvAuosJjhnLyGerC9JZzKWYAhoPrTx9jHEYDlSf0Q0Ojr
XK782YJlHYYCcESco4z73a/NiuXt+cVJ0TAlfCwQbHShCLO756ywce/KaXY1edZP
nzz/EuSNFjXWVH74Gr2vrI8iZC1/ayfs/eS8o8d5sgLW5jtyy4XyOKw3gVnlGTWM
h1qlyw0HPiNEIG3aHL/nbSJlWwjW4HLgTvXf7IN5QqEO/zm9/wzcgOu6DunRQDof
fCCWUXRvh0pWZKanrcRnF/d8nxbQrzlyBIxfMtqpt8rR8V3GQhWPyi/ZVyGaC5Wf
Ovm67GERTgDT42+jtZNMEfDTN2IaHu8ygKOusFCf0h/FJ2y+IlNOOxOeOaHyDvKD
fEKiq3myVcNki17VBHTjj1uuaTSpmK+9RSZVAfsOO3HrzGGeX83hqp0ZBBW8NPhd
TJQg44x+//MEOrPG3TOJagma4/9JUNRAyJHQ5QaxPffB6C7z88v1AghMcvZzZWAo
b40vXdZkuZhYA9kAI7LKKKkidlxIKzMJKHq0JBhhp+fZJBfRg4qw0YYhqqUT4dXq
1WQ3oZQGlKu0YcYBh+EgpfEcobksGgZhAjlQjJ1XPP8M8NKT+Yh6B679cCY1XrSt
5c4aMMEdGuIgsQ6561i9YNcxdRlxKa93X5WrqyvqSU/5MtwR4Q7yYcsqAuhLIl56
hwy5gyzMGadzWkEqYYnlEh6K4GuNRYRpoDwmtNW5tBC2VZzE+doLOu9bBvKDLmVo
YtvsTP/Hf9C5SgbpA12p8bNGMuq6NKSrWGcrRQsu+OGrudXbAhkFNHVttls8TOID
vicy1tF7mKltUNZ5QvYJ9sddvSIhADmv6WlvQGaehJEA4kFJRVgBCu23BigbYiCS
JJSKhkTlyfRGO2T8oK+804u5NbisbousDXbawgETVjSFkKrlp3nMAkEI+3O1huqS
Th92juONlJwqv9a1ZMPdkJ9ACcijvKV5Ak0xxs1AdZTkLQUb3tTrlNq2kQsxQWix
iWHznjovxBzUDPES1v6yiaJ0QiCg9FgeBHOyQ86fPrtLWra2XFyC0Y5j1vtws6hT
WXW0iHYCg0q54Tl0Kp1fto85fEiicieCXN2T+51YVYJ39zObyxyBIg0uSftefE8+
W0HFnumJ7w0uLSvLh+boT6G4mjNLvwo4V+HGBbi/kMm+9hxQn9NNqn+BZolSgl7C
iRdD1E+GUOr7HOzztPQe6ley/E7dWFZ1s679iubplJxTWkdd2FaYYtESkN1uaOjm
dimE/j0R0KceQITdbjPvWN0aDrG6wSc8hQoHektwffYdi2VuIsxCQYFoe8NS+h0E
j5YoeETYl+ksDUWFWZeDVElosGxdUNHuRXaSV3kM/tlY+ma4SWy5qrxyGiJs1Mwe
KJnt1IVeli8Hn3tkOqBYCrXKJqcPRa+sUmxifUyB8u0bSQAdiM1VWlWirsRiZXRw
RN76XKeFr3F+A7l24WkjbYU7X3SG5WWP+lJvTh2TA5L2HGDleK9U+aoCxBK8Abzd
Qw98s+LWlZ8gEQbOcBU1+AapIg44zE+tIAqrd67dxDB4F13hxIW0aDIFQRHd0kHA
tnXi4Eq5NEGx0tWZiemgawVk3KtaOq9NvTFgIathvOU09s18VfrM0A4+pLJ2UNyk
sJGo9x1iqBsACzxzle0UiEjKayi7wdvkiCk+aEgZWufjnMsSrtBNAzRCPE/WQ2pH
Tt+Q6GJbZ3JORPe2x/OwFm63BmkpMA5luyZHBRnsaB2u8qcUWCgXVF1i4Jz8ydvL
zsSARRXWhoW6vT04RLNbHyFDR0m8F5Uwie2y2jpl5bZ+jhFSqBbNGFYyJAdv9aEA
o0Br1R+5ZhAT3DHyO20UDRRZmd6TqGtwUC2/snIUT34jfP2+rmwONDn+sO1ThMuo
NdHN/2PGWNOHsLEYhoKtN9lb72szmDVmj6D5EQr/eP4ALrTRz6bv7znTHAsFe8/V
9Wg74NR9QgNLRvwFaUH03SXcEJp5lT9gVYMP4z9RxyZW68HTDynhLUVc8QLmcE+j
rkneK6Zixq3bGIe3or2i6c2IVofklw725CQ7FvY18iLB3BooDSzPRm+vLuAgrAdc
4A1+vMM2R85HB8ZPCpPca6imoHUSHMms6BItdC+fReP68IV1fMCaHKcgeiUAjhqp
67vn+h6f/47ycPbPMFyBDSgVzYy9tci6boqBI4XnQPoLt6PhokwmhwHi1OG+FKlK
RWBtmia3bTBI61R/JDICK0patG7Sj+t/fUVmoV/DKC4J6+F30qVlySk/WRwus3u+
duS2U5Vfkza+cg4/SAICiFmITNCoIiZPkom6leERpVK4+t4c2qpaTXZ/tv8QjHPN
nroCig+JBLkQUbje4F3uoHIAx51X4xxMaPY8qnz9IqZyYdqP3R37JY9QsUFubDN3
0vqfI6mSgxrVKiTEREXpak12WbE+hN9UYopyTUHwDTvgd+GEwCxgk/K15ouCkdkt
Efk2FiAlcMKk92hZ5fUfZ3l23P687EBlt4kQqFESrTamL5A9Rz6RGMtJFo6iu75Z
sYWHlACDh1Kt36lDEZ3h6EJlAOaR13edCY2L96797DrcDCesXtjVYHOwP3B2+yEB
PVT1Jj3Y05Xf8eWkRuV3Pa5SKBJrwMQ2cTxrIwUPwpAi/ryOPu5RnCcZMzHwuyIP
PVLkh+0TA6VjB8sqxRM5BlXMadRImL0URpRyRsmoO5Pwc7RbdOOpVj1GNMZbqFS0
h50IU58R2san1KY7RQYD09yfZjN/ZIi1xIOHOiDTKYUMArcbUyh9JJ4dmjV5z3IT
HYbUun9vuCIxhQtsr1ooMhMRMhM9uwNfJr7aWoEPx4jsAIz8G1u6WEbVzrwgzaCE
RRUvEex7WBQWPV0ePImlrdJXq7+X8plwdj/lUYB5ntOwB2xOu6dpFb6pRW/XLlWs
BKLWKuXpiFI39+Mr2fDcsUipJ2vAkeSs9Z3ERN5srRinVDICAOg8dir9nw1fgj+m
JXEZ0uAEMBT4UzgnzuetPMpdas+qg0veiwGicTQNiSs0YEYh88gFZlHAlxtUT7AC
agCVMrWPGfS/WRsOTzG47kzEszXyF/x3NOlGeTSunIw4Kwm3m3KVQipNblJtJM/H
VrSZOit6iSNTDpHcNSDH77JOVQQFH+XVc18KMebqgs9rwiFsJv9FoDysy9njKBm+
4vQZiAWH9+8M7kmQORBmH1OXmghNWAe9Zs702wL7AVhoIK/i+16jLzJ81NL4KN5U
7XOsqMb2ss7n0SH+wDDzPB41gYU+Xn8+uPEx8rVoO3JqT6xIqxqckqgYjgNOwQyF
1OiABhLXhQTTAqUL5b4Kc4N4Jc/bBNoyiaymLPHlI4SRK8aq4OrYdjvNe6H5D+rp
4C/MofBfmPvL5MLRXO6zDVChZLBs9G1qZYQaVVklJdRzGKIarVZMM/JfEdam3xfk
JQW9BsOolu/xMgGYe2oVotaH/JaZwxpzGuem7akwJcbQC9QhOSNa0jR4AYSmq4g/
CAeZk7xdIYfbveZFNCFRagm/NEWIpMrMIleJk7HrLVNExSULeIc4RzdufdSFBYPa
A0DfMgJHI5DqFKfaReGvbVWiXxjdJi2kGJszNWqyc6VsShX+ewEJZXanuMdEgIRL
xnNATGQUvrE1xhdgTl3LuZD+CtB93ykyApSyhmOqdV6wLpUHE5pZSihh5AwtkElL
TJ1TXZv96FpPMgWHWl31kwhUgGggGNu4wu+3z0tIrKVQf+LNgyaDFC/D8xq2XWzm
pA6OQ81pnopwuEqwIR+8UbSHAYb+bnTl7IEBSEPZ6PsKWea2guG2V5nnx2QfKis5
vEIek0ZlyWhWMoO7pbV29VXf1ejt6uMv/zqActaldOTYzBwt4psNEUzJkHNhcxfR
WQPyww/Dx8Aeog8+PFUnQlSocHB5VMOMVpfRfMGknkQzsHVetfAdvDjwU9Hw7pdy
rMgrgZpjZRItyLGeA9Rf/+NwSjKl1DqupfLtXqlpC46MiVoI7QCILpb4FmPfulQ6
rBcmrDj7IwxqFhvVtd43PYMH1dy4rtx69dNQJJfOJJttJ9fd1YmZ1/YARqO2T/Sv
cbaWJvGF8nttHoTb/CtNlsk4p711K5uIXFJ2ZPxC3Nu8QHDJd6qJ+S3ltK1SYh8r
fhcr0gYY+cIhbgSV28ls9iZ1fG9qWyVuLQYoMjh4HiEYB9Vl+olqcynX7Xqpsu+9
gGcdEkBYWzpWZ7fmgSnPZpVjoXl1k112iCW0PSjz92BGrUUmTlgX9EuqzrugtWtW
BFShnjm1nMTvhojUKrUxqn8EC7JBFKBai6+TZRzzLTAj67xKnXjig2Q52X1t9k7s
GY8EeoU4UguO1biELvHfsmZal/DKVnyFe4xWHqSG2ZHoIW5Qzej4KbmhKdslQENE
8a6c+GV3livjRG+MUyMxCfks3Ec5ihMcohxbgwtuGI59sL2/391fqftLkZWa2odb
xRuZkw8z+W0NQ288i3IRFtYs2dmKawcvonimVYLBCiVfjSeVwDbPoP/+KhcJbCpT
I9RCUCcu0aRyiSGey7/Tm7bsqpzUDE3eTraah6FAJbf0VuhSpwWPRypHQk6cUq33
WneGqNYuIeCPxEXzG3jwwd0Vqzx6ZOOSu6ysL+6nfHuVSyGmOLS/R2k3pOhAgBON
5lryvgZvny4oQYX/9WEyZbZ5DNtWgfr586kIiCLUI4C4RoDAbisHXH775+8jKc+W
5d7Tt1sbfdZ+1Qrw2V4K05VriPkXB+UOoTL8WPfIC+WKdzCr813VdMv85Q3HTPAY
XxPBz2AfYwbhSRJExcD1sb2U35TtOdp0G7DWUaZzZBXi1JTxxg9QnDYfQjle/qCT
XBtR1++ISnPWtpHQSgtdHklkonvoH4VQperfgTzqtH5lAO+KLehd8k7VaZZtgvU+
eOWBN6wMEzPgw0KncJi1HetxtQs0MWP6comVY1Q88dsmoYr2UZOLJVCstRtY2kjl
+tjSGGjVUR9u7E/guk7Zqdqp9xqoUeiresd1QN8fWMppgqjcdIcjv4vv5vcrlpfp
cfh6+GcodTFqYm02DkDVznL4eNHZsNBepLzOJ1LO/Yb4g3qFxqxTWGVzYd/aLquK
l6lmSu8EpI+cyxaBHMPjcEm2CJH/yLJfGyIp6Sh+f+lRijk7xUmpMK/oYTuqMWDz
ogGlIDQ3mUL5Zm0vLx/wfUkGMUZDLq3NAcri3ytKaLIUdxTIr7/A4t0Gg141Bua6
oTgQwEdrQyFyL0cMFyDuAR7cHIz31RWJLtZQovimEKsiC/eGBiA9K4xhRCIUgzKU
rS8C2tE+l2igR3Q0BKuUOvGF+igr7symJQevthvF7xtUYEVl+XpESW9OGIZqqIxv
pgCQ8PfTV39ul855e5BWBGDtVzkfwBv6XVLT7cfMhWGWljkqD3KoJYnXPJ7P++f+
rJdXnaP5rwS6sEZZP3ZWPavlStdYsOFdEGo1v8aPljSlnI1YNXDeQuIY9Gdf+dse
1Vwyd7hV65AmXxNX92MBPKrg3f/5SJoQpqWw9k9w0n9uTs3iKSrDTuXBjpzzzFeg
O0UTnqM9+el263RsXRacS626cvawVIoyQu8BOgynmyO+ezSltSQ3vqkW1fQkSaBF
LNjsNTXXyERonGdRbvI3PTD+kcrZUeZ1sIO/DrW8oCvJj77mTIDmJN8gshMVPJbR
tCl+sQHHssRWX+2mDncrpCz2CU4IxJQ+EN1erjQfyhCKZ5AUWbVbI9anfcjwLo5o
mL2qd4efsYdXWNKsVh9lNxtbCfRZqwu/X1zPoWluI0bQErr/GD9twmvBbGTjzZ6Y
9PdQhjsC2mYGJ4yeD+9sC8eGqE8tcdjvJ0c+YFxPLm2nXTtkUK1bXYFWkRo7FZS6
0yeZIT1uFsdkf6jF2BU9iXNthMxdOhzk9A7VSZTuXNybEHsy5xtxQU1fBRdLzjjK
mC1ngn8Zsquwq/4pF+8EkKOW1WfPiq4kjxJ0en6l/gf7LoSPlyRjQJrVfr3M+z3m
1yQdTKpa8Li4Xz/SI8vrvdPhaLJv/3p6Pnk4DnrOAZM7UCmMxtdZde7aI9zKkpeV
2VOsk9W0/oipTczH0KagCjMAh+pavDcPWxqsLCT+YYFw3i2fN4zr4baKGynCPUaT
3/J2J9y05U0MOp8ZFyn7av0OfHtPi7/28jcUB1ZO/U+lVtJulGzREmU8qjL5CGLj
xa5pg7JDl71mk+tWie4eKe0Um4nE4xfhI9wq2FclV3/TWu8iuJZ/bVQtutL3FFTe
L3Aq91jx9kgQYET/ZiibwF7tyM77MUWswrNZdmnm63meo6UmhapA45kp6oESrmaz
DiheJZEzsC41r6nE4eESahozzZoxWBh4U5pABaSOxyfQwZG/9DAZaHtFOaDlxUwG
sRpt9tdiKCJowbSa0yvUZ6Pz/NesLQb+RqaPFyidSaeHN/9f96HPQbCuPop2EN65
TM8LSx83LQn6xHk3dxDHmfgE2nDHddRgA3pKZPi4WIyX6PhkoPlY+RndBV7xLjzm
1QVEU7IjEI8tlfwzCBjWpSOHT4AuL+GxNhJFzDbDikeiIqfh2Ej635W8j9l56vd9
dVWlpHAMMa4LpImXlEifAXlFeHtAJeaP3exjFqvNnW0Zy0itH27aR7uPmL5Z/84R
AiIKwvgLk4y/O6HTPbq6E4WuCFgRn4A5+FWXkxhawE4diILubRCql6Tqg7oVNp9x
4nfpuzyUPXC20EUYHJ2ww7Os/Kb7Bi1aWhWYgEq8RBasI8qLd4ttr/VcvKtkk9dG
Yd6We9Hsz3Hs+2pXoTWrLHtXfh05C39zVnVT1YQjACSRd+yrnJ6AlkdzQKHtR41b
/YmeTiIquqgJ4RXkqoxrnLnJWAgDKI/rkNGwjThzP34tSqaYCJgSTGcNN/kd/Bs7
sEKUipBSHaaSNjMeNt5REG6GAZH4RU7DcM7XVkteQX2DVWAs+TFxwswFMlSe9CaI
nFk0JO2dnbJv6AgiQX1fmsi2oaCCo72tRGe9LzoNqRdY9PW14ZjmyqMo0GihynAq
9jCahBxsSXuXIdZ3hOXPp7bimW+oUjEAddh71WdK9+dL742xH08vZbyvPvoP5byQ
wA5m2lyWqIwZg/v7v/dj1Mls0zRus4y22EbpqsmFLIqV8pVgk1IKa5gafZhF01+8
i0gMYwFcPpVAr4v2BEOMBENxVv0m71eK/Chr5yyAk1SCxIQ0H4Mo/1Hp9UjVgR90
X/OweOzLlhmSBw3kr3ZoOqPgbuCuTrmIT0BGBYXjXzSdok6hdn+mx49YBKTL8uC7
M1IIE13ys2AfmyRbibw8d+oZKIfPUXlQyljH3CU+XJkHzyEfh+r1TqbRBsKVOlmb
U5qn/SrNV7jVyZmu7EEbOpPsmVRo3tVmIvhY0q0+vTy6h7njhwOYT3pJi4EkXY4M
+oHUVFKurR0xYHD/6S378IT/QSB5w8E8IjTbB1t5zgJ5zxety/tdTwkmGgm1k02c
pFNGZiKNCrGWa3umR1OvY7MUyQlwxNvCgGMg1wYsVc7On5NWJgOMnLNJfNlcum3L
qNeGuP2LK7T4+TG6Dl8z4sMDduF7sDY2QOgdQHU9eJTlsMa/n/9tn6lhui2VUVaH
W5kTiPz5gTFXCgGwobPbqyEHIsKWFFWKCAkDuinkpoR2twtRDJFT21HHhLdbLtj7
QDuePFqXZYApI91XGlk8ylJ7lSHs+s0nNohwjfAU7mfQBhPVSdEtZmMN1BQ5lQzV
od3BvIKhEYFBTaDOkVmDZ8n0MzKTZ91f64IpMjy8MI+SKHBWUPoIsj3Nga89nMML
rMo7/2apgQg67W+gu7WV1dhAgtqVWcjrd2Yv5HA5sqOzj1J60PFq4sX9c+7XmKNx
JaQoNcWe3TBjUUDnFJd+QfwmwYltI8gjaWwmFQ4ezu2v0/8N9mIu8LlAMrQrCnaa
exjE5F0rHmB2CdTFH2D1UmXSvDicQCZzQX9DtNdXuGm+PSzXLR2JBOtieN4pHWUJ
+YO8G0v8fyD31dJU11Qo70125A4fn2zoErjBZ4YdmD1sWJHMN3lDfGiV7ihH8Gtp
Z/2HGOhsywRJCNxaCd1gtMJ83TAJkVxCdbwOFhi3tNxC0bsraJkPZciI9CERAU2i
MqUiNCb6kfPrnIYFrO2SkE6Dqt6v+rtVvIyXjRS1OIOMrCas69CzBpdjC0cNDxem
6gIwXSism7cEZwvgab1BI1HbNHnb8uvyDSb7P+7zsgqne4FaJA30mce+LMOPSBHU
Nrlk4mZsax5nvCE8KTojN+oxVAvLx3sCuujIJrtFRP2Fzl/XcFex39Qcz2V8f37g
uMc3vQh98NJovjTg+JGA4+sHQ2pFS59jqm1yQakH6I5gZYcOU0g4qWCAzGI9h0rh
mFXMITlfV6QCh9d+9wyiQIr9lAwIM3LYMXJ9Rup+tARTiINWObotKfKYn4cuBAu6
znUL7Ua7HiCSk/6hzP4KFHLGlhKQVVySmFkBA4x0mGvQbL3tm5VEp/4fO4kCZag6
ixcYDGxX3H9UL5G1e94ro48GFNRAd4eju3UKdnZUwWJjl4zqiDo4yqoQk7UFB0+W
vkCfaMKVClsgNmtPCY2n4KQ+0Z4ADpJhKj/Hi9CmR0PjkS1wGafTf284qlgPZaTp
EpHFwAEKi6t6gp6krVmsHkCLJIxBShybvmvkXks5Lym5OjUsRYXHjQONtFKZOIdi
znjNip/WagrYvp3Azeuob/CHO3PFoeJZBsysXDynIv+W9jwWBQ6cSwY+nH+EHv0i
D2idCJfe57t7UPJXXcVeflhKqYT1SXfDr0KzybsBE1/gO+DEd9QSTZKuChqwstpx
dxm1+MhVrtY0xHVf+Xa57heccol4l0X/Mb+vhVWS+qvyuO0RXPJ1cakW5la/C8H+
5zDe/y+lp1NdewFfA86TAcxxCKuN+y4PkZYn9UKJZ0L7+7LxT5BFPgXh4cuMF/0A
RhER96EBI8gxWh58jaYqyltLGIUXl15K4fGbhW0ztmdCQHdJ9jBRe4p0OuGPxFBn
ieIHL880TTANmvMBZc6wHOKAoQ8xEw1/kK9BwEL8vB3liBXrhYEGDfHWYiFxItKn
ZUJ9Th3jq3ji9mjRPDQd9f8Xlvv6GqgJX5Zhzv+4QYEuyCqCXiCW55sigpzajhoa
baaVutR26tredfobdkGf/HJpWSnZtkZg/BWo7rGeWvV0k2Mwm/pRcriiX/XCvZqP
3K1eeLF1uINig1T/+2+XF/gjODzswcvMYLwtVRRSFJ7IB6LU32JpHW4gf4fM9JUr
aTAjSuoFSsIOoqjKi2dkLZ4Lb8t3LEbmxa+sgO+ZEJg8OzNAQOkqnNVG70l/HiJ0
9ZMlolD3R86nxjp4DJnae4YOR0hPm4+WjdfMhyY8iardumTauVeVk2KwY+TB0Thd
CawxY4VQks5pTn6O0q8sFA4TGLsS0Rscap7HN5NYLzIurO02raC9cs2sj6tJJkua
3q2R41bUhCMMifErov90RQ8X4U7UB84qh73HQ80EWInQtGs8XIwlJ02MaMbel+Dh
7I5ILL3DdFG4GqgsMpiRoEWvV4nJ99VCmQ3kvDzQQ4C6QiJ/MsNM3l8AYdgay2S+
bx0GA+XAO40gOROS2lXAZq+/8mLcCmTvGUDU6DI1FqMj1vOApdN2qYyvVsns2z2D
9w9MiK0xS7u/UjNOUDVASzibUKd0rVAX8qp9jRQpJF49A1XeU303PK1Cewi+vQhv
yzGkDy7tXR2kqFp0Ky7CgQwvMwhlI5hLHk8GEBAOuI3JhwVAAg1AOGLn32X/YMFr
710By8N+KdUZ0k2RtVmzrym6W2Fxog5P+vLeMFD+1e50T7EtCD3OsBSs3CPWXgXO
PyX9HblPK7pYXeH1a0qJc46HzcHxqrE6VD3fQ8J3spsKATYK0OqxWrcwd23aBSiJ
y4ueBFt6+i9s4vMhlGrugWd162N1ktzzzBR4VQmxNp6qFEejJkdBsLXtB/H6Zg9G
UglyWrZpV3s6Ge2RTVSIyWTh2sBzp5Fg0JCVwHnLiV0CeDYb8MSr+Rh9LXe56VqO
AXBOevYKplT/LqBIVX3Yu/N+2G37o28oSk43uPghdd43/NI6U5XSaouqzr71Fuyz
rsm+ltEhOtDdxkJirwCZtMVdRZkrXMKB4KtLeOAoxZjFL1hx4iJlez3X2D/Hgv66
twukQUc5jWC8tPciCUh3/B+/AniFMNiHNqaCUjhP5v2CxwMBhFfoLpqyNfF37m04
GpGz/UsejGTi4vk3lIe267yTbo5AsFuNKH7ECPJLX7yF6ZvYJJtUvupWAz0VijGh
EnxORIG310I9zGeu/iKbRxBRkQ55H/VfBZolQnPxmfrfupEqBpOQxe3nqMZ4vmg6
I6X5hGi6ld1jEske5RObPnMi3i8+wy6GanGfjzO3wF/b0jim/TcIk12IJNgu+EER
WbNODtnYZ9wSkxvzfTbe4RQCZrnas8wckbM9mynx+diuZaPkO0EUWTytk7YxPsdw
MOIxazqe9h8ozbz9fUx1lABqJ7yHduqV2yuVLNlAEqe1J98pykyyI9Jddx9RDA9r
eFxclmM+gC29RaTE7XT5SMuyj8cSqcPCW7VZxcMUcdzLn6nj4+SHopYk13QYmODX
eKkUflVkQ2DviXjtADkOKw1vjBa9TbEgOLd2GH9WXP2ieimHqN/++QN7wnDEUqjD
qVSieIHeEWlAv2Q1xuP+YRIENywVeoDfo5s2jOeDm5U8AdfjyrmhaPSVQijMGU+r
81umTKQAeMdUosDixT7SbR7yK6kyYvWce321VRRxhLF0PtLjRIV+BOk/m7Cmg2By
Z8CTE0TPtHChnSOXBEOSpm1l2MTLrbCw9LsGgV+3GrKva8WslLve0FR0f6+vVQ9T
qy42VMSr5z7BDGFMMHbVAcPdl7pvoASEGuHe/NsS9jdhn2qtOOXOnjKJPvGsKl/+
z0w20S/irmq7XJ9rSLjRXdCJvI3NUcW4v+FfsEoKu16ABGTpaMb5Ws3KOdoM3s4A
uqZMOp4NdfN/Awm+bmCNjZv35hTcjssgrELVj62pL6hAcGyWcaROYndKO4GQ561t
hWJbee/hQpxNmBw1gVFywYOOhUlIS0GaKusn6uvhaGMKXeS1dDaep5Haq8lXx5lP
D+Skvshr0WWSC2lTbgi2xwujMeyqWHR8QSFhBqZKBWvc31PQdlA09Ny2ZTd/elCe
N580fBsFYxUJOf7yzraDnMb4e0e9Dz1v5pR+AHDpAJLC8HFThX6TmlFebL8MDC3s
iH51qOfIpsSRtecGMBHrpC6mTcLScYDVrTbZT5rnEM6MxARv1zKRvUWlLLUq6NyZ
EHDO/o7M+iOnCjgKWUrO0XwRC+iRMxZcSz+QOLpz5JqbeCGZODQX6pfMPvRZlPrm
1fJM1rFc/UEg1YPoi3D4AmIhMH6MzXHFmZ/4Lh55SXJQIOr+OxqKu13Yf5xw/MBp
NqDNtvjRfYfrVE/kdf28bF907qjgPJ1j2hIX4Em6PDtyuc20EjVHnevuyvZMt1D/
RbCxRy4LFpRIGnmUKMG1SZHHYT43W40nOasRa0B2tXdCN9QwQ/dcHxZL65ab67El
W6KRErZ3TMcGDp5vANPrka0iZpmXAwIqwGuuaRBKF6JMwXTOmlfWQM0NHUf4hAfY
ON9BwC2eIHnj4NPoEjaYbmjXjPWl9XmlKFILqxvsEYZVeG5m+TrPMATRpDv746Eq
MRUAOkO0SgTWcQi4Q5fJhbUERTtIL9JAaMd7L37IVY01TB80fN9AQWjkdQF53Let
CkiCUoLylu6yrBhPesCfc0O/Jiisved6Ts6dpF43ILA7ZMxvSmASh0M2rwjmnPLO
6xKsNHbFDwHm1q5FkPg5t5h89+WS6ei2YkR4suYAZ5VYxRpDtRYiLdnMomQgNzXz
UqWUETlgDX7bMrhZ2EKH878072yMHWRVIDM1G5u5X3w0jYHFOI/m5YHX8FA49y/S
lJkJsouRTaNDJWFb4eFqG7fKOKAYBxL85lt5rf1+gZ7j0WPLDDwmdu1wq1fgKkhS
WfL3zHGUOfXXmQOsptL+Lf+WxB8mMeF9SOMf5kpsuZnZYyynfpfICrOivuM1YqWJ
43jjhICRpIB/xlGYk1SDYH0dsTBiPvvQUKCOjdbgOGKE6Td7Tjx7n00RvK3pDT8a
LUim3JA7j4/PvbXxpa+ohNjTJkY6Ih7AkFtvALvebbm4bLQd7sO/sCBrmkzD3g99
oWlUCJtUOx67rQjBi38ltqOM5MeNqDkZrV45Qe8f05AVG5pO7+6FkF+uVzZVMVyk
AO79UjQvOo/ndiGTF7xU8oZ5PmwYioA07D2EbvOw6CUuA/cqpvXAotcvghTbNO/R
Ekp5dSpKN3ytACiZNcvJSXS9czqO/XzLgKFD/6y5aUOhTDpjxXJLzCKSgQz2e0x5
xr57qjZ5NmtMMFVtRUg8i/+oJL99AHeZHo4BZX8Y9oKICsV8U2ulcD7u9UhVq073
tibR99J1jkfXcHaIxQXINS7gae16i9O7xqUfk0auSUD8T7Yooad36FcJaH7GM8Iv
Fhp9i/pvT1p1yTndIp1/hNmW/Ow/Jog6nSrorVkXvNj9W0I/vNnBohbNYEnfgeAp
k/LIu4gnFSP5l2PxfR/JmO+5xLzr94sJi/3OYLMBurXSWvvB7E6Gk0FIhO0a6Wof
U/IuTjp8JWnvX/0RJUrXRtJEDar8yWE41npbD8ROuYlGnF62temhyqNYgpzFEerB
oRXBvco6rXPexVk9kfWnJfG2yr8HVVNW035DfayFeoRmcHaBoP7hTO1npNM1v/II
WzI2KAQa5nNc8cICUONUv4bECj9kMPatTneKJo3KPw+kqFLPOccrdYSDP0O6DFBg
94iArGJTLOp9n8FRzCf51RHfnTpD3q8IzeeBjWrd2+VuvUWinNnWOZy29+NRWC9e
CwXZPYasH/aOc0xDBK9GHvJVMVwH0A0+jiMtTqjqoQTP+c23uxP/51FiXhTbUtHh
TiedWsljDoMlhZ5sezgMXOPUf561VjviFiLp7ztPDJ148gxKR0AAfujGx3IHXFkt
G5pcxR47yZBmCmEQvEEtncFqG9pwGstdB/63zHiWfJs174aenVBtNbFKEXD/9c/A
a7kqTVas4G8ebnpzkFh0GlfwT/vCAJEZGTrXd79/lvvxGZezf3Oa/2mR8aFLY3Ua
To3pQyzPsJa8bFaEWRiX4ZvnWgBdTH8AXzpzlvNBIw/akg2cEawlBitAYx0o1uLt
E7I1WalGbLIZi8yRAR2aPJ1Coxy+0yftpX2sNVciPJAVy3gq/v4aSR8BBYxr+/D7
YpkljtAHXSdswOlNp54SpAvfnEo2JqQGixi5cRLkpP8ahk33XPQWryKGkWrcrtRY
Hi0lFW9kLow/oGCym5NcGNmKUUfMa6N2ISVcZBLU9CJejMicNIczK5li+pTVNNik
ZY1UWGKb/+pWBBGIZqdTh256dvmS3pPmur5pD7U59cFHHPuirBWAm0NJi0+3SQy0
LaDNjYxmWGgZebyeyMmDQwRa52So6mBr1+avmwO9IQ5YmzswCOb8LpDsK4U5/R8Y
TYWxn4wjEbgBLu8EwRQCCry5kPwIohtwqdp41lESJKix2WPizR6aWUbXVpgfG4s/
mGyip2Ke058edFkqwSjG3tTMxl9lYyklXdR3lULOAoAfhULCyaZjMyaUq8MvMwj5
txcOrP1pR55QMX2NuXHxEnKW7TSaqfO2WVlP9ybyjZBBy7G5776TMHLBHAsSvDUv
6slC4H2/LAjdsume80xQp5hn+mo13r8nBwWB6ewOTOJ2AppKJmZeqHtujtjkWlld
JPWBRAIIOcIqxEZBYxKn1v63YSWdXf7pvArRBQo+z02NovshaqkQ1QCY/TleaQhL
K4NYxnv5YFsJc9ojwgjujd0B4lQOQw3HxZMleOJeorQ/YjkKQAY+YAUyuChoJB3o
9ykqLR6BsDu6LQ3w+JjWuY/oIIln5G3h2yOjYMYu9edRSvWN7QtkgBFkFXatdD5y
ZzEfenzclm7M7AhloYw/ONhMpzfCkB8uX330LjdjjArh3TAHIZSzWRyaZ3zSPjtN
SpfQpKNs/q8rL29pobNSjJtOwHrnHXNZOdjuAbdB9cw104TZcurMO5IrNXyRdHFv
F1Ut1roJQHoP1qSasO7ShPVevzmfdRtFuYUkXKGDCPw6nGG60f40uZIN4Q1MmxL1
mNRQJDQo7SmN1BBkV+HsqWXNbuU2fUh89X5B/BkcArqIrWlLblMZx8MKqLwFZpFs
DZRNuaK97o/GnkMJM1vxfY1VB7qx0H1+otbfAT1ArjUhJShVPh+22bkeHsK7yfeG
OnDajv/c+qB4LY9e1TGHdI5GMZAo3hbVDe0uNo//JbvQ+T6dfgV55ldjxryBh/KH
/pDjkUen92rKfKvpQSdl+3sQCcB/sqSULnQEvrLO9Mx3adWQKSJGHP6dcYyq0P2y
troLHtwjuDUWTicXEZPEaLCFYuh1ivbllLKQzlt+JB7D4HJRCM3luQPHOyN9WitG
Nu0wViE08oSd3U41A1E+K1gdAX2xu+UCA/erh5XMCigIJ82jYTt1n7wfeIVwiwSN
1PCADcUcYaRlZY0ck42aIgA3yMhPu4dvvCy6BhF7KtD1xPcgKQXff1a1Jo5bInAZ
1e+O9BCZSnD5Dh8h8B/d0Ou22M+X/sVOFTzHpMunjRhVAs6m6yWUtsplhnZq7JLo
r5/XlP56klBo7LPdWS+s6jYJrpjLGfoZuNoq0vNBGQfzxFAbk/5wyO8mWOHWrU/u
AckuhOu6KqAFb3Wbir1IPmoOmu8w4AQC4fRy1CHMdeJYBAzdecqqzvbGFs3Xm42d
z6347K2NqTCbsK2SiYeNmMUV85ure4kVCjU5z3wG+IdgUHlrsAPzy+ljo5Ni+IBp
IgOcOseuABofxjpO1rZ0Zl04gXEmY4VmonfCq+WGf0AWLw3qvTeMpo7auGIm2QuT
BVCOyI94ko9cASMUh9W6/eMcUhqGJ42qPzK/HVKlz/5npJAvjqFZCr8IzXSOIKeH
uSGIn6B4tCGSDYe/9/gsnW3VtLxp61CIbHsRIhbGJd8WWsmQmWC4oTa0uANwdkR3
qxyvTd22gVQa/kF1q+4sjxRQiBtQAUqsYkKUXW1QWszByn5cPmqFxOlmLmIGu4zb
iFdSdp8K78DUUI257q7boCqC2GXFqMwUQc5yhl/yhKOeqvCn0skXjRPqy2x8MrV6
8SaCNNkp4jkgzkZ5EDakhjBL+K7UTw0BdcLs+G9iGKdjxuRAk8FqhO92KVIKWEUv
jVhwIzGDCgon5CVw/WACD8xiDmvtueX/3iTcySdupBwlycQc6AlZEPN+g/KFlr5Z
YEpU8K2p+fd2lP+KMkOmA/peASKU/CyPZiRqJ7/sVTBXMrs48l+BRKvQZ7Te7TRj
4JGPFf/HzNdXQjFojAZgFifNwJH7nuTYL5NPyQ+PpytaCyOtPRKqj6G2NqZ4XA2v
toToM1GVe4YwKaTVXQA6kLLwh02PCZo+DULGp3xdIpqXLjY4QltBNUVBZFgey/XG
2ywUkAffdyCsOSsnweYxXkNp8ex1dMPz85Nb9JUSu+oOINS7H3GGHepGZypUDhvt
FSy85THcE5Je3QFCgiImjU4zcij2IZ2wawtSnpPQwnRiJmwmJ8T06SyNDL3bjNWP
HijYdOzDxKgz9CxvLVv+OUNFqB75Yt6rmORonIdfgHtpLahGfJcMEbkgKUWi0Ayq
7MPqJU7Ad72QTemzsCjf7UU5h4W76sLM9UiwdyBwed0hTiXIsko32cqgUUPVrKRj
58mTFFE/5g1pzdY4m7cQuGWk6kiMLNq3C+oW2XchLjsFEQnHtTt2vyGalLO4mSbE
wSVMQDgsJuyiI++vgtknzXWViM8P28FYdskQaPYncLymhUGp7mRGm7EI9RCNR6oP
4s0cCElxH7P0l8sMUBU32GvTFUUzgQi9vRulJl9KQ8pJCaTVlPnMW+8ctyOaByaB
IUHutuc+2t7rPicdRmx3rmbL9yp7kpLmoFY+5Mz8XtzT+LgLfgI2oTqTqtv1ao7J
rDZyRl5IHtDU52/6m22MmjCSn/yDmVZohk2WADPQV+6PcsSDKtisZYmvin2FB7an
FtprGCL6nDHSXxd43b4WXobn8a7qmy3zsDPbLMucxj7QFK4q5LX7AsDuOw8hdS2z
8KBoEd3FwbH/wTiCshCF/eJ9vJDzMJ8d9+EoJEVI4lfpZ5Zvkifr/st4TFQstV2b
DScxJZGF64OTjcXALS/k9s1hDEh2kr1rkkJaz/W+QXMHGV216W7Yn9eDuBI5vCPu
MbjsiqJ5B3Khbne+un50Q/nzVBDBiJ0CTSF3e6KwkH6sjakRUIAwdOfdghrDCfcU
H9Zp+xR+GlwPUyGxypiQNU3Ra831FTSA2SKGojMQx6cMMB2VeBZnNTcbf0l86g8G
mRXFWaGrjFvNw8fTe91r3Y1qhMgAq2ujpedSoiCvUyCD8DYNCVcM/Tj7TU9r9b3m
FWJy92ah5ZMzOmIdIWE76p1kc93dsatQ7O5sYQvSOUw05OvGB1FWBwOnQc8q2HVV
tCPS6YZHCclfSLCz2bdtnUQGYft4QhoLXelhdZUTyNfiQxZpDzbahIcHtRcMqPgi
nsdhcdOdoHROu0qjJo7FAC7+S5OmfJ11gfZiouahwx6iXjuUutHwW7W0HCGig7dg
wZrJGX59i/XMlpkQd7aJC2qjL9A/h92K3yjJeep1ix9l1ZiNJXTgqLSSfoH8r+BQ
60stcAWCFWWzUSQXUb4JwI9jcyrKlKbeF9t2fxFm9EHTLUGXjaTvFLSMPD7UXb24
4/z12IfIzL6ZWVovz48eZ61ooD4VisPiajVYUeWsf2dUBUPqipN7kxyr5HS9Aa8w
ZJnAvZVOmhDG1hdClkHU3LFSQL4wcOsTy6dkebmlYnqaJ9bNaWZ+wFUg62OYMzZI
4+DtWjm5b2sMm8mXPo+8nYs2P7q2mat3k7lU555aMjbk4gkkC1Z0hQ04/rpScZRP
YnWRSUUHUFfG/rq/hZWDGNrWohZCoTIjmXAiyamYjrh5oycColhGOau9TSGGTsu5
q5eeJRrPxzRcyVpAc3Byfz8EWo9AZ6jqNdIVjfcFiTQSj/Ckr8Jo6n7NKkV5HwP9
Lo0cYX0fri5JgTPWwRgVNX1ii1lKhw2iwmIsCLeTqRqRNZQTFVo9sLzhLxxF/Gx5
/4zhfi8NeqPeZzb06Glh96Aw8m83841nQTBpmuSkEGZ3Q6aZWv3tGCOcApoEYmHr
BcyomUpk2SoYzFLZGDX40rSQB060RQ5LrilKkJcZBU4ebjEArcqklswmz4Vnhnnh
/4uHaSBrrxPmjwo/MKIswgEoQ+BvItJukjEPUj2Arh+5s/CuvO+awwftYzT6mX/6
meRBE3/Uou+DuAtUKk1sre5zeJwS+kCW/7Lr9XNmWvEls2u1H8s+03WQo3WAuBhw
rgv8eR8AvXd3bbGN8B8Zfnmfkbltuq4IwzuHhxywGrTJ4HBCrOix/25iFZLSm7Ng
/6HUKJaJq5ra21oGhgMmq927r0bpYsOGGXRGwOFZMyZSZCwxL4C+YtafFkYyccMl
M4k/Y2u3wYfchnrp0ZhyRhkMMWd8xPP7OjtbHQqElSk/zBHnHtXHMGB2SPhS8GQ3
1m/S0fhKJ1X8jTGzM0RO/j77LxNFWT26JCfB0Mjk2L3SnxKLbkjM5efhIQ6DBDKT
onTEH+oogfO9MxfIBW/Dr6HvBF2TA45+hsu9+l3zvPN4LG1vjkxizSiIPfYCyurj
nOyN3nUOm+aharSOEVLpXs3o3x867aa/PVV5yc9TgzTjj7SAkxTRYdvWnhKCtdhm
XTJtHSzGydQW1GA1kOsTvsPxYu5/zuy8eg+MNkRXJk/8RY0IY/D4JHaba55VD/b5
PWhWfQ+SqU1EZZNU98iZu1ZmAICCRqep6DdmuU75diszfNwwzmnTPSTsqBADfE9v
cgYYxhxWaMAYJJ7BOmL6xf9glvtWtUw9s8ypUHj0u5OFztGqXi288fuPTgs73Fdu
ZBZ7lMS3L9cXCOUr4/o3vQYWIRzUFDGRZc65AnIBtE/IShM4aRL+oJTDRCcwPft8
7B6fuTmzqXBPV3N/0pVKKzhQOUm7UDVVa1S3LSO5kpFAYOw2IzMMQcYpM9ETfZc+
AODnwl61k+JiG0DE6+Kc8NhFLHTgiZraYN8zcIEua3BLXuFi+to7ByxdI3Lhf9OY
NU1Z5cLC9XkLYXn04p3MOf58tZRDMxHpHeVRUofBEB9cnK8E+uLMqo0FYV0taQn6
NTkuc7c0lEEM0jLyShdBgC5Kw78U+njqsUADYGMdqKzJz2vJ1SfM3vwvC0nQUbpk
bM6vsHMfmbF0FeG7nu5jbBNzoARMA+71wNBUNN5J7wIvMEapsuCJcziQlDVtkrDe
v2tkJFNAjd7UIkNwYvLCQE18/N8Pk/4tfI2dTCHQ63rfaW6Y0darpoAz23Cl6GU7
GlAXrdJNSmqEwIu0vu5LKwNwvo6+/QMURDFv9ws/xKMCdbeL7efaTI+WBCT2OfzP
Jym55hhu6RijJV1Y01l9C5JBrVIsce1P1L91UYWMVGvWVA62xACbDctt37APukwm
bUCZ/mm33W3Iufd1creMxRzC1Sil212dsthyTi4ADXvW7k+l8fptJ2LssyPHmgIM
SgW8A+wWEESKptm00TZ7oxXmhERj5P6QC5ukSF5+se3u78ampqctJLiVvDDx+eA9
DINwQnJn0wQ+J1PPu9Ioq6OAI4ewUHdInd3i6z5kFcqUo7Wsa8cWVl1L7vU8gKdM
kppN5yy4H7ieF5vKDysSvgLRjKo83hlgy97/KCMHC0x7HV+vzHsD0O/0XdZf9P4A
/3drrJ9oFybdjhUDZVqQA0CHgps/7cddEDsXs4Go+UCzHV9yRMpzBfaN6urT6sHj
5cJIbZMoF+s5JTzwtsW6dcB1V4QaorocWzttQ3dRwUwxzDMPJQkTzj+ipfemco9t
k9g/UbUSP1WnPOvyK8Kb56KsHeJcU74mBTDcfVEiF97mfNJ6y9jl+i4bBLzpzwU7
Oc1XhMLBQLn7UnI+Mks8SHOMp2Vb4Lrp3VPoJN26Va+LB4bl4FaN/KIk4VJYBvwq
ylGA7lKW+axHEOEx0KhZqG5ryEjqx1QiQrNDWl4TzkBJ0WrfIqa+U5iBnQI94E2G
dEe494iFFmFReglf3iqA195emthBacPy/wopaUMCCDB4tFod/PsnmWb/b0na4m5u
321/98dfAl9v8jhSO2hb054n1s0ezTziQw6lxJyngwKb0nFNwLmedg5fO8U6bnqI
l8lLX5630OHG7OPmss2ZG08IfA9lwxvpD3X5JPOp1BWUZrATH4RATw8CezdX1LJB
ZE23kT7jnq6KTbb5wsCR6BO86zzKWqWTI7riIPXeeStPssMFiH+jE93j0cXnsDQ+
LpmJt3rLBH2vCWisNZsSK9Gx3X0ppxh+8e8RW0dLYDfqME32dTyF+1ZNURLaetE3
zJ8zmKMvELuYl7b8Ynr5AeM2FLb2tC8SJJZ5dUKBw2AqR/sHgGB6cFM7Q+eUTQF9
fR0OSnP+cmjCKSS+By8jmWeFDGVYXdgqNJOsy7OZSePJSLhhFPfZ44RzS3Em2Td3
OvqE3fHyb6OPzLwEQbxR8Y8B7acsM1fKmsVOmt8U5xoiPbUpXzhsijbGfIAoAJ8O
+NTQeXS9aoYwf1j4HUydfDCADX0rsHUSaaorKJuLYZVq4EyouEK2il1Mnm05Nn59
MFTYDFAbHhI3lehLIwt+rRBcQMz8XhtOkmuHhi9hmzI3nYU7SQW82bp2uk+iH/kA
FViW5ivixZ7a9831VIQweA359DIx6OHG0ce1uoIpnbKUkXrQU7ygDgWR0koElgJQ
Dvbgz2dCPrY1fM2tl5RrIzqag+/0LFy0W905guUFz6slP5Y1tzUk1J0TWROxjojA
a8SDIrd7yE9UnoQ3vX97O32voOTdvRWc/hnaWHeTUSudyml3Dj8dWrZZyjMmKwuu
nZGCy/awPz632NfPDvSWprWUpz6od0QsbzUIigG/GBHzXQJ41oWcVr8Y4RNVveva
1BqEchxVTJAyNHEyZUJvn18EDWnUcDq38MRRWaJlTVS/IG8QxzZ5edRpqBlVzXlF
/RpDUUBRoseDJey/44zHGV1ZPXL6TTecFey2EbiLffZbPy2z54O/zIGbYB1UQV8M
sWrLHXqRVwcLaRogMu1NYhPVk6v1jM6vnJ6UMmwuUK7aZforM/cG1BMVYZ46uIER
GquQurGmPKoWwGRmTLGnSQtmcXWOkUTSIqlSrOgZUhLabZc7QUprAlC2UduLKDd1
FxRCc83L4VUk/H4436MGL1s72lnM+E6rVzZ4KWB61I2SldGSuWtmp6/vQq7bcRFl
YmQTvIVRCtpTJ2YG3kHdHt93t/Dh1DhwiBS/D3nPXvj19+gbBcRUdp5HnWBbGBTr
2hJb3jC5k/HXp7AY6xCZrH5E7FM+X8scQQq96C8q9axBAzt11MhhX4upjnXUv1+t
L2u7DSyAmUbVGCjixMzIG/b77fC5K47aV3/st8mFBva/SSZuf9UT2pF/m85N7IjQ
2SH2WpObKoLYMJT4ZUZV/xXWrqmo4AxrnkDviZbChO9EYhGeLoRLQ7btZvEsxSl8
TY1QtyEvAbRJlMokTjOfDIWByQpohGZLM3ErF7AjZ1X1vVlOwaIl/dYtOh5D8zBJ
EO2XJsHvxLmCMiTxMd/uT82aPY/9XqN7GyYJkI0qbH+XXWNbOR2MFLkg2BuvU5Tv
iihp/pYY1Ty201Ht1ECtfJaOnzE+uXucPCGKY/EgAUEDBjarGTQRkzpe7GGwxfxg
16bkDqqpOXsFseyRPWrzD44RJeZHslR0/gcGyyAqc7kMWCo05U9O/HQJCk4b2DF3
mwbcXlptlTI4Y/ikOj/3h1ftV+h9r/XKAnvnFsVlU5CQFUV47Ca0uvsKCFjxY7iz
3uSjndg8lEbrkJGSq5mkLjP7KWnAO16QedO3XqWi5wooygBGazUstuSqDcthyEyv
xpenam2mZE91sFaoZQrr4oV7ySjGCV1D2mHl6hcjgxRa/giGohoHiYL4m4VUemMo
Gma9by92OV058QfawPXgn4qScgFAY4XWsoEL7LfiuxV0CDuC5oXGELUOo7dlgUbr
om117UFJYxC6NwrTtJ4bt3Olk/oBlngec1sdky1HgYZLAhIMvZ6VO2Z8YaB+wBCZ
klojy88IjJLqZMgsQFU1i2OcVa46qkjko3FyWACf6HLi1C2an21ANWaxojAo9jzs
fp9ZhEhVFv2+4T+yTbVEK5LDno5tury6Y4S4Y80/gwOKd14Z/tNAH3VYR9q8Go/U
LSnE9C6tyS/b0w0kqBhgiZHYpFwKqNJZv++vwwvdp4dVc0KPJ3LcPLPvdWv1uLFH
ayymvcz/2dUlwWpmu0dKixqQL7Uqug0CGvudpCnu0PM8ewkM8gXxXl2152Czzdnu
WMDOKPmT7FT4BQsCXOyl6WCWiOQxruaPVECiOTXLxbIg4vtbVHLS+3llh0V6qeIk
TtVq6OlCHnSlFL7khGSFbufVRCUF3hQkENtdmXhjog85s4xser6uXHZpk7CP8yXB
lvDk7RZJeHZrdKVswHjIOS46kMtb1sX69wD+EPL6QbLAbRL3M4E3pDQ6EP5q8VFc
J9C8wRVL0EoqL9n71Lm4jKWvEu7q34eXcmB5rXxPcDdOnNcvFHgqHNN7/t1xYzNx
RJkY0dUDvjZtV3dRkYDJNtQeGbB2l3Wt62teiGEbJ9GF9hKd0uWQVv617gq2meel
aFE/9a2H2ECS6ZQszbvKKmNGBlesmCw7US5oUQVvtqkw86YprGQcsBS2d3cORipF
3wFjTdBK6NPPZiX4/4XPx4MBtKprIBwfWQHcs/lSCxkeEhTNt7ylz76qBrmqBJr8
1hzRvlQVkm1O/8KrKIrf0ZJLlrlGgYyXSEDK2tzVsBVOPdfbi/FYwfCTeUguoSgj
XGyZyl7gN2QPDUMYCHlz84cRRZDCF3qZbu2PNnK4Qd/IeYfj2QOkqw+MQFqRvke9
vK55w2sabzmQU6mAHh8DUiR6SCcmjB9UchrKAxX/lqxTbewt0AOEV98w/iIYtMUb
4Ce6Y9FInpQ0/BmM8m4gtEyGxjZxrm/CTnvmaFxSQ7a33Qpuox3f05p8l+shDl7r
PFxHCGY9RFnJpS2yiEQUoN8uOe36tUucwutmiUkQ/QC3d8E9H0D4A8Jvrb7hQf2L
8GP2KfqA/g6xkoAl6JZ+IrcGghL5/th2icrHuZT4jIlaE/6PshejMkAqeXKlsMC/
2Gyr+DEzsCE7LYiCqqrBN93xs7KNffAWBznifs0VhMMeGRfVwLdwHpomt5SRQDug
fT0Ph4INVd1e+yjz3U5eUg8SGlWx/2ANSRtqFrhzJlW7G0TBNAs3S8U9QsWdI8Ug
COU0s/pTU7S+1olILy5SCTHxzFPzAzod1sPwoAMcL+4jBRhs/lLzmfb7JoIUsp/N
QrtrsDEFoIh/eAZiDENs7yimEPtsKCeKy4PWBvDBH6MffWzR5uo4XLfj6Xi+w9NI
RvMTfWLhHDxddKVukSGWhNwIOpocgGe0gscLnD9zOBPJI7D69Xl9Oka/AaFjZm8/
MXwHJHp9hALSNMkR8pk1J7V3edHwVbzPAielwzhUXlpCj0oTJ2FdCPrNiCs8TEx2
SmvJtGRFlPvUbiwetQ8xc3J5YoZyQ5ocZasBMgtanrEk6PDJpP0Wq8Kj5Mm1GPJf
Q34IcLWF81aTXdeHQxNJtm6ja1Z3FKHRtXbUUFijBjMKI0xPxcRtbRPzAMrtwQz6
63CdzGRKiv8ZcDWs7uKCHnTiB5qjs5FeyreaZaxe2nKZUTpoNjQaN5lo8kbtpYkL
neFb4EiQ0wzW1056qd/lBpNHeOjjLGHBq1XQ594leSR3SW1SgCh1qjzCEvKdVEYy
8k12cSSq/3xX8STW1lHUCcbOMLxZGh45ePjFzafokMW784qmT/ec4h6n/N/j4Mbs
NNHftnaEmo4OhNxXK9rZ5r7uwSEjNzsjCfWYgSVS2sCoHj9GIPH7kL7vpTDrnRZT
0zH8VSyauwvWSl9naRCjqp7UJVfGxbdoU8XWHH4aL7HqvBGK2clUxoyGKRQV5XJI
ZyTDx3PA7QiLHTqxXVY5WJYMpbp1jBU7JVCYXiTywDGXX4O+/Euz+pPhKQDG3jxk
ZwriP+smuwosFBgZCyvFg1GNFGlPAHWvoVeChBaT6EY4J0eLw8KlS3IcKHONCWpd
erKRfJoBAucwstvgkHB8Z3xc5bdUqsCGqvo5hlx+3TdiwCIfol97IbyscA8YF+lz
yX/J1110u/yigT7WNEwZSa7txJa+0OGRNPPrtT05P/+gmAkCvj7uFGpissB33E/f
VSRfo9aK4mL3sWsTlK0lqpyiFoIzDWGgDVA10XUtnN9OunQVyk9A8XYfhtF3tSVA
3E9p2BkwRuGlaSscd5HkOsW+SgtPAxn7lAZ8wSY5OTQvLISiLG6u0zjRJYEUrTjh
St5ZqsgM1oteKwOmIH42yvv8c85/LsF8IFmunHJeGeXBxzCqlafN0xDh23pNWlUr
ui8epqkxR8wqdlc+oABug6JFeea5F1Pz/H7MC1pfmzju1fZBC4aywVZ6KQVy/Atw
tSYN/NQ5vkiVvCC5LRu16IcIJkmXijv2QBzh3nZqzOwRfd6Mc82zT3bGH5Tkv6jn
y39aq8Zeh2RfYPcEqZN4MEWpbd01kEIFcWMl80fLWA729A3M8W+2nDMvd4W995gt
T51MjlPpVT8cFdJsXAmzWJSW7F0DTccHem2UlQ/7Le7MGxGWmwpw81hZxi0J/HZf
8jFXFkA4bR2SvHCqAubahnWmoLXmJydifsAeyQvaf0djrYmWEm3ohoMQ0Yu2Fsv+
nTtIVP/UmXSVFkebqnzPrgv4YqdVp3xVTAymOaNy4/jiXGgX/GSPPPFoU9CtcR/e
u4CPYJWhvHiqKHtJhZzeCg6pBXd9/jh9Ti6TAd3wTK09SMzy8Tc+RVpLTN5klqoo
LbHhTUSw5uON6YkT38SN038MK1NcwsTJPJ06fl/qK8/OIstv6JHA8rSI3LhNXJ96
+R8Xd1Tvxl9cCd9+HOHAq7hEkJtnySs+A+HQRO8AGPCmgd8/iry4LCz1jiVC8qlY
H+IbiPdXEa7IMWfBzI8geIpSWQmzEw/4qTkzbI6IHhYADRHd35sE7PBomOq5ygHL
eR9Sby+kqs6V3pqeSQw/fUN/8COZ/7PiXXlkH5BB7/BeniWAzTUj4Gkk60ZWDB2m
NB8bT3i2AODklIgEF1yEAcziJxYLJ50rw2HKBEZzgOQtEyfp2xoaYoeALivo0cDK
165t5q9mjWOmsIsdfShsCFajTTn56nmkQicDFIzvH0oHdxUaVDDvl7XOEkJtIAWF
CgM9kcQBZxMqdf6qMzsGHUIylTnNWcIbXf6CV+mI9XwTiiHcFEeIAEzv8o5NrNrk
ay6PaAypYJv1iVr/TjA+E/oNnquejsmviKCZdd2Fy52pQcEkgVtFHHYNygENDnqP
ssIUNMm4jV/+xVTeZlTmnogDOS2dDggyM88EtOWYrB45Bv83SULLhcM/g4O/38EP
8xZYW7jLW+fxKEBHHo2aU3rWeLEYy1Q8Ysu2XtqC43BMZn9Zy5BhQWc8DPYmwgMP
WTW6Eq9hgDNVozRltDquP+0WOVXE30pJtHPFC9IQ8I6R0TNviSQUP4mlsWBP7iJW
XUksZVqbUPjA9Ew9SBM4gU/dTwMniYdbRiHve6hQnN/2JpZxe/2Y9eX53kH6O5Sb
pq78aKZrOQLwDQtF+C1GQO+2R+wRvNnVwdBSh0c8wb0amf7I79drocAVYhMmDZh0
n/nuju1MWQ3Xi6OtfAGQ2AxPyTJLAK0OV/04SKJZg9xyVMfANcoqIsM93+K6e1PX
WG/XSSIRtGtC0wMR69VVwlWsiU6gcpOPKm6ypUtLRyRRFaIgmhMrimkycvm2hJMA
G67/leCjVL0+Razt66HMEi74X+pctWg6mD+kOaV5XLbIWWLq8KBhyKXi0k7EDolk
MHxXVrgKsbAm1Fnf4ihEe82XjLjBCdhMC4a+LNyehC1iahfAQ9qAYgjm/kF3bohP
mrv/McUhRRT/oG2nRQN2J8VM+JJXZl0UmHx/sFi5cd6DmTx+ELTunbXt9eVRWlIF
iaJk8LDD3TzzL8Yz9YsIm9xybTtlDuzYe2GCwmkG5mnXgK7OIAIpJ7NSkT4OuN2v
XK9baa5/f2GXLKB9nGAfW0S5KlCDtd84wb9ZuHKOKgqInTJuU/t080/9DKpW/IF5
U1dlwj62xJBDc/3oyIS9IoTCTAqjEQChvefe3lMgo37NeicnBk4kQrONXpzE7DYd
RjbP6YDFMihCbc7bx07T5zfUaw3i1tu9Q+ZfB+YQBn7HDHenJIvTi7c3w5gw5AVN
wT0OuhLF1F/L9riqIibwJgPwRUbVqBo9w6oXchOTpmgX87FOUjKESzR9MrCI6Fg9
1M5xqsvS54hJdsHrFeuh5xrsi+HGnCrIkU9sXvj5QxqU8N7Z5JxcwLXbj/2Ib2Rw
Miro07Y4qY/yQ1gbZATQ88TaprJPhVLh06CL68aR6crbl3Wb2OJxuS95E7fWnlwp
nWbFO2i8TyRmtBO3QRtTz9mKwMBL7grh46yGwsOYV8XKxc8S9ip1Fr0M5G3NmICS
q4Uybm9cLAcG+wG/azeSoNTbqCrz90Vo3rgKrkKJb73wC90KhW99L1Dcn7Yg4HlT
NPASWN7Y9PHiLRfhQaNhK6TkFvIF0Ki9e7tczyutE4xwzvqd9BeofS+2C3dUYP6o
2u/URUyh6pHKVX7K2SLH6I0OQgZn/nYUEcqHDUGKRDvRofTSXleLFoXVMYxHIXpR
6BImGsROG3FhxZt7sM7RYHXehxYx0UDGbHsGur0jzexfuNSfab5fBnaDX6YLjjbf
yQbeGr0TIl/eSsosh4pFUv8oGVaV+N7tJlpbltP0DGqrCcezknb4wwXRpS2bMHfp
TukTgOUaKRrBjl0pRaq9UPHKRS9qWStBSlskJIgMNOARhKXBQT0+RAJiXzDSyCeE
OBgKXw3K9JchBU42vrj/tE+D0oQwDYIXAM7sT3ZHjTSqH/owBx3wo3353qeW/GF3
RktVIcE9ghTvY7lhiCrYobehtyvdTGjZ/6Hhi/5t+a0hYfRLgb1AKPmOHv0IrWVr
l23y2t8rxSzpVZbxP2LgjkJ9V1fcQ5bf0Hfm1svOrsGHwGlH/HXPI34SITIfVnYb
2A1b515zotngRjl7cdExVYHcxrFlav2smjaHYlfVeh5BtfvfY7HgBAh1d+TbLUAo
jcP09UWOr9H/jBM3niW8K28GjPHNEHP3g5Z5neddf3Lgv+cZdwoEX3D6n5C5zoeU
Wn4mvPML9pKKS8idauBtFRQYx6w9kbkktPG8PXtiMg3gn2Be7CT0fAXTmmX79p4C
mxgRaDJa9KJ2rGnm+RMa+clDIoeM6ILtsMvWs+Mp3Rfqj/44FoM39HNQHDUKq64b
ZQbr7Iiwc7gUief1AZs5g02wWttxjUafxnMQkkPxWO08Zy7T8o2eoUgPIEEtWiIx
GwmprwDeIlcS7csZt9F2mc8NeA0GykQ8eiMTIbO2+xdecdWjnjMCMIIgAaZmcVjj
ZWx05jFmsQgoKrCV9f1s+1pLbxBCUe3tF879p8GbfFNiq2eWBzdmBTMLfbzYSCG5
04OefRwbLlDk4EzavPVxmCVS5/gnbTiNgPNEmVeWQivDlxnLyos28IrYWccyq48u
NVIpcycIpHVWZcQSmxSxSxBFCE2z8eFMPTZ9H5a8tiz3FB8gwMXW74WjEFE6hZ9K
815ZwOjxbRsZ1hE/MRmQsowXDnMkVr3PErGtd7lJ2wysSgyng4XzPxtzrUOO2Xlu
HcohGrJ8GPoX0iiJU3r8/UVZcdnhOnSXzDkDXN7w5Sn0If4oKY9jav2zvLnleM0U
PdyghEsBduf452cfgHqQn5p+zYCqWobk+lpVJdrYik09GZSVQ09xV4pEBuUizcG7
SWrG6TYAvor5H59W9iH/Um6XBHb8i/0OxePWgmj9lAcTz8rf5CKAV5gN6SwwM3q/
ofzXLChx7ESizncP08Fdsjcjr5HUYmmMtjx0/83MjDw+ea1FWgw5W0R6g2BWPiiP
trLYHH+D+CCmKkO/kZGmeHAwiGxwZIp9lq87OXdVCkr1xVyKNOlhPcmlZddFg+AK
VLmuXziGn3QpTNnKShU5Sb6DF93DgufJZhFy1qkB4Q+rxFq7081niY4RtWxCumt/
eB6mkBT0uDxm7Amxcln1lctOEiaX5fCoNFdSwFuuOU9hnF0fuPULs+VRSdgHLfD4
9GX2TBIBpUenWSXc+85BOiluxof3jNCx4DMTGbY/YBZFYEE+k/JesE/vMV+iAYSA
Hr0BvfhoMfxDB5dLiCvGVqA812RcRURSs7aAxlRw2QMgxkPq7MCn7Rm2VEGChqBB
eyMoDtOPXnbtPVod5xQhLwOqEtiyOJ4x8fCOYtm6kSwKRrWx2LpyGmRxX+4Bxd5B
2AiLUUmukQ7vMbroIVt92Xj76kWaMr2z5H1wKd/poghX589gXfIkaC1e+Q6EKRDQ
JcuA55PbSeIpTmKzmUKkamNbPYsiczsz6T2NCBWaMEj2R2rxIUwQExtfpIgO/dCZ
Ml42x6ToPh6yl4WOn2k/jLrRYEikzBKHpfyByDuRq1PqAvil2u760T2Aji7lDHG1
bW52uGx4OlhXgjwjlpg+Xq5HzEJX5BJS5kKp5P4CCQQRvYWkZ8POeMBrcGOG27l3
8/C1BwdZ/ORMhCACIM0QGSz0oXB+x7qGco+CMZoyeHRCF8oWEp7U2nJr/mQkmelC
HiQiYvyCV0hY+aBxMIbC7b2YEwQItKlgrqbGzcqiIJOo2z7Ilma/DPtnTv2Bw3mq
2K0K2HXZ5eKwDZafDjv3CE0PHpG8c8Crn/pGsheletzG8ew2917fKcPuCYmCsdt9
4EC5Q+juacHn4De0oSl8sTq/XSzeu1MWgPbBsiOO8RWq/OkSJdFVouJk7HWYyj4w
8TUNwMBUtjj8ZxbwNaHkDt6/BIYrzQPzfxk8VBppOQM6FRWjJyGf71yDLsPvyG1F
OLtR+U7cAvpbxmg2CHaC1/tpynriHoSWQGemqVOMPIXaSLQTK7unlJKil3jLOpzt
OQGicAMajfzj+cygcCY+TeBQ09uXGeh8VSw7LvefCPR93FyrlN4HR1iKu939B/0N
/Ns2j7tgTtKA9KBEz1y7ZaYCk69jpCjIkZa5fmos+qs83SZ1K4GcojIlOAuI41Fe
3R8gP+BePgV+XjJIv6oQcg/M4+4MOcI+zIDAif+L54z4msWqtZd4msEQjuU2/Bph
7Huc452xk9JgPzvMGj5Ov6IkPjwE+qGeP1fnIsXNOC2UHO6reBGD4xLZzDLPKCnN
dr8wf117HvzlbkmMdu093kNVnDka581NurLMS/fG0PVHw3iKyK6Q1rlzQL70ybkd
WJTcpd9V/mBvhtExRitbW69Zg/y4j0e0EcxHsu1Uh0zav9C5mZhfQ44RvO0aj0ny
dc0hg5cvJyN1YtvCBBL2yWHAxEh6nH7okmBJ36W8EksvYmuqXqSHDCXchErZfgyS
dnlePP71NdzGOISD0yE6Czk6KJYWWe/wkIoDtN8KbyP3D/KEQshY9p12c+VMEGHm
ZJJRkuX0pfQKWw6eJf9BqDJXlcyOrzkfHWq1XlcQFDeKO+DmTzYJynAJqN6vkyO1
dA8h2BZCnlKuobjb4wTxrDiGPhtBfJ5NVC1/+jMeyZMx2yhCAcyL5Kcdb7nPn39g
LtVzHU1mtxCnTreUmL1dQRvawGvNKgoZxlr6wV8P9XoYMlpDor1xy7n3TnOgvwnz
SnEIeRoFLE3hFbSZSB11jdpKcXqdwObcADzcLMBstZpWaealowour7ZQHBaw1MMp
JH7R84n17cUZpN46NQXSPzk6oKzmnI4SMU2WuH09yG4SsOCz03vsIrZZPV6LVXcy
HIzWEdBEYalJQoKVYQQBCPBx92s+Z+OMo0YnUt7EftmusJEWigVgTPGvg/oplpSI
YGLD+Jpmx0NOSp8FX2VUbqc+cGAZQMO/sqerk6XqSF7D2ZFVI+B9xvJPvZV3757X
BNojyfSNA9BdKQefz+p3gv/zkPKXpJzBk638FRdkbFvIQEpKyqJ1XPSwdSiip28v
giUW8xd8MhMFA6y9NpD+o1ANtdVVLZK53P1VcSfkyADJOzyehDDVRWyz0dQkXARV
uL32hiAoq+uy4DTwlAgtzz7VUeUdI1Exdo+xwOP5pvaR0VQh4ToCfd9J0NRHkk5+
zzXJPLMzAklQAVhpadzAI7Iv+TVern5IkSnm8Atn6ttWe+OPFDIkRhEEZIpAQfib
Dw0N0AeXv4jiDcGvZANEd1sXKM05AkZPqz+i5ySyO9sr2fLaJpC4xPjq2cMc7jS+
aloCxYn5IU6QgVJJx/RTASRuaMjv6fpEJBQQ5C/dLJ8RD+GPfFAxE0bCImaCyn+l
VzBEjUAEiqQS7AIRPwl/UAlMN5J4sXmOapC/htksRA/Y1hv5Aqh9cfKvRkGcSclS
SXmO6DgmE7TtoXy7nbZWKkks9s9O0VlboQnhdJ1ibq9ZE+A4uYdbMdaZ6eH4ZZAX
wcRFAKx2mW8ACQJFJpY55fX3d9e1c8p0YXnnwLmM+ExtlmO0JczJ2mSzM1NkHR0b
E3HWzbjcRdjvnCH+G69dVpQx7RdtTA4+kKG4YyjpSn/M3X2c+4klLKGwjvrTyjHv
Yd1L1UQWwplyZTdfURhI+gqRZu340zkDXmOm7fuc7sMadkAgkfzvAvzmUlygIJu3
F0MTy0qCNtj5xfaUHYSCLzR5w8Ey7oNIWRwJlTejiIAE+i9jszdOUMlAxcRM+Bc3
s//BZvbtizt/S33xiytmU70HNgCNsFf2mzmAFqzeQfMZVrr5jFLYUllHKL4emKVz
FXhX9Q/M4irwV+xi8AEMd9NK9pz8BLamM4xw3JFIpQDoj1cQhZCPhV0arK5543Bj
45W9/WaiPYhIviUAlDkntw4eHFchbOVUiB4KtQkUdz8kwwsNqvLyvP79UcwWFrDz
4nUh9iZxdtwbboBBP/E7JcodOtO1UzWqLOj2vWfwPP3ridGsaqc5syARn0+58Ot3
JNrSuGnRDmdmhz/B4AW2kAzzbmaIXJ4H9Is8kTq/pc9PtqjYGUe96S3ryM4f0GeZ
UcT2EoarIuBk0G4uShuMjwtc1vv9P9A92trNZLZhhUEUd2Tv6g/tD5bLu3mfqC9A
IstEGuPK+rJ4F9xWxAE27fu3BDSEjTPcaatWqlSkrU1cOUBcw2L4SPyFc21K+aTT
tURCRgSeZR1uNu+VW313sGds5q2dwMz+3ZreiaGgDOd4U4P/lkKVztTVwjCsoBqb
R56pWD6pZ0KJU9h+TWWlx84B4J8pFSCYuXkz/+XQ4NRS9G64QgRPSzP63tpc4TQJ
ivCkpGTLhWuji87UjIbZxtHBC74HRZVst+9A56Vam9/ThoIargYZWCen05U/X8CV
rbZCnwY592wkEICW1F2mjNdHYK+9r4Oi0da/AAq9ropqONMwTT9eXVTBFzmUpFzu
UZHMkOfhMJQRenHt7/2TmAdISnA3X4VnmHZkebiadOH5j/Knx2lbL85CJt9kl2pz
+1prnCbP+M+qCjukRTr3XWQwsQvgMDC3xWSDzncFFceDfKB/g5WUcTbLCVPD3qp8
sxUMEHxnQORH5ZOGHq6mrtpjloVoirs4k31IGFxx3AWb3U+aMXcKL3LpH4OLIh60
s/dYhmYGKJWDGhIw+dIn90XT27P0N5nz4TnIswXxBKqNmessQ4Rj0Dy3bFlLrlrZ
dADra4Q8Nd6VBaZXh71FhJzBlPwo64fKo1vTa0izxUNoAuADw1hWioYELMo6Ca6Z
00wijyUT3pQ1effzw0H+ScpF0cB5q7HJHKLMCHPUglDr9nFzgXYmDUyYcBR+j3yz
g/CS/3OJdDA7sEAkn8Up9G4QCC0b74RHIgV3F3+5FtlPILsaTvQeAlUL7ORKGecl
74Kwq7wKr0GRTRONhpFhiRLoyzdfo2xlPh+Rj+BCrX4jx0eECWNhNKXJ9BWTWLGN
RD7TrJHkU66p1Zr0eIfh7dWJEFgAvK0NzR4ugIAWpP3WxVJr+D4EpjsZKHAu/4Jy
P+tCFb+ktd+rbhH/Rnez0JTXblQFvbV73RcGVQvf4JBcBWzmCGJ9rnb9TICOCP8q
c3hU/43KE4wMTvaNzza63EDNbxnkyx24dj0XJM9XkEfPiYNsvUPsZS1GRZzhrY+0
e3KAQZdJbXBug99oR0aFcdrcJPYFRgOu8pEg6GvUO+lcCr+2LGMzF64tQo3uK1eX
Nmkij5qHMlb/dHbV+EoI+FnWAhksVC3e1WRFEvjzwCo3jEY1VmOw7xh9s85hfBEY
7lVf/RxQ92Pg2yFNRCYUFUzw/1HtITG/0+aXdmoCJS8XkFLr/CwDuEv5TGOW8pd9
idxp8uHenkrbEIdPL5Eq1WFHLF4rL+Oet+YuGdiMu22ERpaH5ze3O1RQc5/WQn9a
H1SLedvYaNmQ4Mwc795DnjE11BuargxCqPdTocf7Xo61P1jX5Yd2PTl8WtrE810y
ewGv1whnO8Mx/MaHgIgqzR1LL+6AkNeyiUV3ZXZd3QJybsi+0xTErgdA6n5KBUCi
EiOT0JjcJE6cDGqDI5vpSxS0uKgfQMhpdOSjTi134CjfZ4s5IBlNCtnIVk4ozLfp
+Bz4hrlk5SEzc9EFmilLsYXLEzmaipGzAuF8HqBcZMCBYpVQyZz2VIVFUDy+hQ6n
dvJnX9bnpa2UI8dwsnmWoEa5pcR/oxl7D1vT2dCADrVxT97PyZx3k89UjDAfsSMx
AN6fWPvvlGPFoLtbvBdh5TRJFtK8msN3akmO8u0PpvGeRH1DFxSirNpNUZ8wqurg
7R/IDNVdrll9B5Blu4+xJgqz4VKv/Rsyc8SIYRJqPsPxFhj7sj9t6o5cZI3Yc7j8
cDbZCEagon3FoFoAHG3dFrorbBOHM8UhoWJXjo0sX96C+UDtD/AF+y0px7Yj+xDA
B5mttdn2G0Jk4t4U7IhggUTNUEwsv3Ma8SjxSXKqFWqZq4JGZyRD2UjHhZU/ikDJ
/emhBcwh2pBwqcuRQMxvUxt/Ug7rRBARFFc23/0LcfBrMGd1SNJc6LsWuPF7omY9
Gzi8Ksa7k/nqrGTHrXpGKgOwPieeAj+CdVF4ICbWVgnSpHcpkK6uk0habhY2nHBW
+cOP+biCMxkUjzMqy2p8kLoAHA164k49+rvUfeifYv0hZ5JcSr+gqvP8dbnicDjW
sfMC4ZXkRT86SXdQ93IkXRv1ypgY6NFvCB2GFv+JLAPE6dKuylYVXljRifUcCi8m
eXIx90UtGVj+hRR38OBJm1wxYqtSQGGHwVIZMOHxQDgxjewmRgQD44vA1XeJP+vj
Cbe4VBTxMP066RnnTIIa1yYAKfXY6LcV6Mqoh9TLF2gRQtOAdvhqGPV1RTky1ae5
fWAfSTI9Dlf0mmLZ04ulPUBAi2qa8UBumB8lBdoWo7eLvaGzSzaYNiuG6fcU8vrP
8W3mzzPlbd/PRAANF/Szbr5Fa/TPEOYFG8Jcwqv7nPG+89LOLqMun4CzzgD+Et9t
OAcogMfNfqkHGUKhbqWGEMVx9/S3JkfDXmX2vi94gXsB/UV8XKiATzW6Or1dANwV
2GZDAL+GqJWBP6gSXxamvHODl99v6LZJZlRoBz8PJlXwML/IoQaW6WLnbciIPkmO
58MuxEDGq3cq64aEAQDoPkCnWcLIBpIflE0y826GQfsDzgYXko+yTulb0w/EiuQb
FDpFkU1/ObEL4RR7JKqsAflvdrHcnhesTqrsnPwlvaTi9VI+8S27PHIjZ+ixp2gG
RcgKr2qPkzroc6M9zcs2KlNdo+xnHXMsd713zjgen1QmBYjFkEYpyQjgq0doZ847
/HCxwufcvHXlk+9DdcCV33e/0xB4ddBmvtLkhsFlO9beSenfIM5R2GlXL1Q1zqlb
bOX+CJl56AxE8uMpp+X2R3DOE2HhpMzefLpi/UPCuomYbj5/PT5R0nZSXixES/sv
O8h4ly0ZR3LiOrIsTttR3NmWMwc7afJF8iyPauLJa8h2E4VZQUlHvhOzDHyyzWfO
RseUorUDNiqS0qlQOQdplcsMQcx7riE2kr8iZMcOyZ1/vO9fSE5Fpzz3tN5tIonc
MIo+LwfXXpL+TZPUPR13X0RBKTQJKBPM1D3cWTovrOKkMagWdUYfdHLD4VMiM68E
LjJUoIy8X+PEsVFDsq8i6uQ60U7eTaaZof6vlRFP8dw0qGvXRB1mqfkWler8Wre+
ro4zn+xQTCWSGZAg2gkv9ToSMQYScnAG1LK+LfbJs0gnE10mxxk0g6A3zWMQerR3
rIeTfv/TfWYIJqhANVSwksGW6sDGbr83JrL5z2ro4jBY48MhhswFciEtnTdvs6Iq
u6z7Okh+tHXomB2xIHPUAi5XnkE/bvxQBVDOU5sYLGeG1vUG3quottHE7TrvAWqY
5w2+UZCC75MaZ40J5AZrgVKaYKOkRWfiGsDZq2aszRYadFbYhUofiR7seBbmiZvi
bfueuh/9KDZn4e7qe4+q0juk9OG1qaHxLL0A9pZs0jc3qpJt9tzuyvhoQINRvDwV
qjFYOx3bS4DqvzAfwMaY+EBc+i3AmIdD/b1eEooV1U2/PR9/J3O6+Sr8zRMYtpH0
HUncUxSITiwI7shWDetvqTWC9u7vgODDFKPFKv/y/sCs2svI6rP5fBh/6GHeSdPy
EDBaa5bDTCMQKFoz0vJ8yxrszO1dbx+8wLaOyIirT3WsWHwGt9+8dJszQFr+YW9E
4djnZrWhB11KnfnJT51comR3PUDxaA74dH3dZPwng4agQf84xjTOog96iu08zlf3
yQrbh+GU8zl7iKnlIiqtk3spIRRHiAVWAqg20lAMz4MUx50hbspuRU2KXIDXe0Dv
g8LQQZDlYqoJgAgch5iiWAJIlERa453SJ0/7lchJoek51l1vkYLE6yaTxY1KYoIs
rpN715URgqVP6+kFyjzRBFrKEwfI1FD2YLJMLtFs8p664zOfTbCN/i910bT3v4kC
GliOEb/Fr+mjjlfAzYYlHKaD22SbJVHsT5zaXz0FB6qR2dvStu8tuUBiviPZVezz
tZSpFfYSVSh7mHk+NVEq8dGn15HsqWsQZR/p5/Qa0gfz4WuneQIR8JtzhDxybDmC
YIWBKaUF+0P7cx5Q5vajKTvBi/6P1MKbscPpKyrZN6v3a2ZfGnSAPrS+rXrz909Q
Bpa1Xr3hzB+gpVRSpD1ljn73j8p7TQ0nxgimjmNs7Zvoz5d/DvqQn09i0bqIgOsM
lSeT4jxf8bqWGimsFU7Iwb+eFGhwINpW536jE2KdkNawS6Xsn+5ekWEwuan/yxCn
fDyCaNhlRTijEhSb5Lp0AIMk1UkowEZeYta4RnfFlvVyjHYw2pirB/LGQPbWDHgM
hBvw7jk57PbQo91EI5+UdEwOwAUbte78snC1ENoNWatMUDR1AqwstfmFmlDHmrpc
HZTgRP4pJ1qhIGltpb0py45+LsBeLC2l7ge7g7C0VigXT7I6vcLBsB+0LAugL/vs
XGU8/su3LDgPitY1fSQ6Lcw708nbAlgLocg7bQ1tikdw4bSKUfxr9U2MFrkaXeaV
KTfub1Vy4f2xyX2iQ4Ms1LE2jGOKVw53CG2oeP4U8+yOObKd9RztDSS1vF3rXQ9Q
kJ43BuoyCLPTelhJwYI+IOfbHOZXnvYc84/706vDDtoLkI5rMw6ByuKQBwyLq0eS
idzCAxxIb9J2nlotvgN/atV72798BJXxGFnxVxGTLN+yNyTFSqj3v1V7KYsY5Loa
u32uzLlJKyIE8JYRMjZrE8W7FUWx9b/+lYPcS9ms26NAXvijqO2IZmuFI7Zfo9SM
ZrcQjrxLUgcJQci39drAQpSmzFSd2RQ6WuR0Lnroi4TYCsyWLTVHCB/9Ed+ErqYw
rXufqB86H5sXf45DxWTqOM57m3hYQsEODAICky5XNY+kspxLjCuoVGlv31XOt5R3
uJ4cWuT/Vx9GQJ4GonRJNO2a9x1WtUK7nfM14gQv4aHaeC059/eznlSNroyjeQA+
J9tdBqWqbc2sgU3oz6iBt/totJ3idbhQAzqm86BIB2tAvlpCQkXFkvAu3tUUaIdg
3n21h6MxquvVju9kvvhB2sLiu1CmIOtuOEFOQ+LBsPbcQX1/EcMgUOHnCFeonrjA
MIrmNHcMT6BlX3I9VAn8vljuiCoXWlxuYsZnTDKjRyE56oXVKrm6a8vsX7EqX2J2
9rlf0dtq3AtNhQ5MVGLHG6H3vngVsBo1KLI/2uiO5xJXcih5p5oh0nJ3D+kCRIZ5
JZ8ZshxBY8lAqPaXv6oUUyub8BuxSQQU10pjkC98X3CTPvouKLI1WU5SvXrfAbxp
F/XYx9nopxTvANNHFn+PwbjDbDE1OzjIKOO/5Mfz2wE1ErXPgYA1jv2Mg1ooqEpM
1OlMe3i0NnjFy2M/zzI1UviqvlJKlyd7vkGxYcJs96wi/fMRm4rJs40nCUHoRXov
EvtKP0br9q88fx6AgLnfeRs//7L678JMYPACFhIm64m4w8Br+QCnpxPojr9UISeJ
XRNBt8JDaB/1GsKsov7MbLBpDwfQKQO4qD6b+AsvM6yPwD9SzlTPppDAVs4zaSHE
VcR4xGkSHCUVk+LW3ZQ+nJzGI0FW+bThv57wm5mVU5kkzatiHlz+b2XPjntSWS8F
nihRZ35nxrv3LicI6JCVsmPXPLascw9mXuxNk3lE9QHNK1Abwgp4kywJEstCEikq
kS6tARIdoAZAow/NIxjhJg8ycVMxts+5i5nBwIxbpV97x/99htnIaH44mWLWKEnR
FPkp3jze8z5m0Joad9csMrbcNtuIUUYM9r7/DaLE+P9w29XGM25bFJ3TO0WQdLuE
zCdh8xI9g7ErcsaC+vGbTkCrjnmCZk2YI5Q8oDqN4EAXy5xQf5h+Gw+lE08hywwL
D1hsfb5Pb+UW/UtbE4XF4wbRtQ7pImE5fTmn2xr+8oi+2anS5OgDJP39flGdKjSk
d347OocrW8YVd6j5Dr9wq/Lj1FPDWDTDufOUR9igTvwXbiimjvaYxpn0qGeL4cjI
2Pb1NHExIl9vJggTz+xB4caXNsJRbvCGI5xRQd9TL7v+AqWptOaGIyCFYQO26ClN
YweFJMbMUW8LiMJmXyv21oDT6Xk9azZW+Oxu/UVqCJ/Ijs5WZ56ye33rcg+DCsaO
YCIIS2uxb+34JiVZFPolLmPfk3zsMq9yQTUcP820ZP8ni+5cBRypdQ1jHYqnttAA
ZtqkhLI9p69dq2zmEiyay0SQYY8A+YxTjktiKm1vSBRyrnE2qDm1T3YPIlCo1kTK
+SmrDIPzGmgnfTld5loByGcdAXrvDKqNTtlzzzLeD0L9q0xR3T2QjxJmw0doR9Lc
iNDlFH+y5NExp2S8b1A/Rc+4sEdzGwVucgZHtoBMc2hCBEjtGDCsagcsEGitwxbq
ABJ9tpZ3fEcpVxZKeJtOCzG6AOJhT4BOhO3uPbmcOlXnJuQGFNBltmxXCwDxvhU+
6kv0N3fF7Tnqf2Zk1NpGXhuLieNcqSjnCXlb9lXoXpaQSSd8TtLHjTy20CsNuuW3
37n37itsjuaGDYC9N7qG9b7WXSxAIjfgotUAAIFenT77UJetD3g3zCh+9TZ4eB8R
M4dOiDFt31I4fnSk9VimT73yn+AO4wClwV/A45nfazoP6FTHqLOcXGQSm1hkilwF
lOjvD9VCIo8E8bwR1Jg2tugaigaBoD0+13lYWDri6vCh1cl1Bu+weYojaYPaeFVn
hBk/MYtU/kfe7c02k+wN0yh0RKteA56R4YSpfpo0lvZTA2ZEyZL7iri8mey9xLrw
zuISYBAMjeaRrDwHbo4Y+TXgdR3H/AjHA8t8aBCMT2odbRGjvEBDeoqJ85EEmo7S
APXY6sh6NQ/jII7lSgTk50Hmz5yICZZeahKXpgez7b41VeDU3VL3nfOXzKjpDO9F
JoOKuqVVE5XCaZWNCEIOAtkpQDprImKB/uC4eXqJkTgE8zSFDKozqkCeoYe7EO2L
EYJqbPZlCaxGGJb51+l14vwA10csnhHhobkJfpo8wFbJxiwG3sHyqWu14jhPujg+
8qv5y8MOFk/wSy5lCcUXtzq4dlshVs5i4hhvnzDyvcIo27cvchYqWcDcSdkGc55T
Ia2WMxCJX8kG1Sp74VVS0GHKg8iS2axNGG8qXCmZNlOL9CtE9V2YaJEo8i4BDiY5
IcJ/2RIeHWJ/+ZX8Cs4zL5RFMQI0J6LKIRoQ0GtVHiXrQrv3YaM6v4a744nhVmqI
U0kX0twOkvWYUije+ZMaRZfQaohN0NgaMAbpIoqh+++8Yl0FnYwJsTol9Mw+WG45
yMtS/2xJz1fMZjbncas3ceYFii4yDaEV9J1PFAvcwvCev6HD1UARojquiOD2HrKi
/tP9p7kh/ZmdPkEnSRcbqhzZHQPKEDxXiMCLomD5kVu7Y3NOwshLKSEt8xv2Y4rf
x9z62BpjYKXB2bcgxjZXyETCy/YHGpgJsOo9Bjsp5B2HzIHS6MBXE4fpcQk/d8Rp
bEetbDoyjuS6bcpi4JLWIx4w2TYfqq3sA+bFvby29EHXBIBCWNppnpJG6hspw8EK
L+X0r+SEcFV+FyEmq6KpQn21ezybhVjp3FbcGLv1Q7oAmfOOo3Bcxm6uSlAto0kC
Ly7f6hYa0MIv8dxU67Vi3ycNxjcuznt0bpSvatte6sGFe5l6+uBB0vhEUgSmtNqh
jUExU2SxsKC0Of/PH1mqZrlQSmvMbHqCrXxHsCTv5hGlAjxzI9WoRSlUQNBnwA+6
NfZw3mp7LXFezFk8BBqVjUtV0PLd00sRZchkc6VLZJn9xZuqES38ty7Kl5i9bSQl
eaKGTEd0z2XhE6XxYb1fLmetEBnchV1/52+Oq8g87om8LjU2jjbZMwc4RzhPyKYX
+xzA1f2baWva9Ft2I/mgFHSYB0ATWeCvWA5WZA/q7yZmk16/0MGUQXxiADrlpzkZ
5uQFQSiGR+rCJ5H8h7k7sfrpWnuNfKb0kscAKB7FFi8DpCRzpn4hK0d4tHZCm1fm
jdFhclWHNj0foaWlt9YMQFB+Cg3073+mrvhn3Bu8XU1aUvpTzoiPs4mFZjCAMObe
zz5UvTITDBEyuizL5T7SloWDMg083DLJI4ml+IvewXTe+cxiSYHTWVot1p3l4cuH
TA7wmLrWe0K2/oR5yLjDiKoEVoMdkeu3T401IbNIN/C/mkPGIUafzso8xAA7RDWx
XdDX/cPMb6wRQ+tjM7ada/aMoVpqF0Uo9Do3yYXLPpMv6A3MS6/XGanW3j6My330
pALksMjOzrqNx5ZBLjYccGZGIAVWIZ0a8SqqFoclC+vyH9aHUHt+QT1MH05d7juD
uwhA7+XPD8CghbOq9K7SeZUI8G/cdoqrUy14AadmlkTqg29Y0ExoozjC4MsovWsd
eIal86IYxEVANDJJMR6CjQnaMmqUuEx4a3BLg8gU4hp3P77c23OaLfPpDc+XOC7t
3NdnIg+TgjnXyYKzsXiB/pDl4Q8LNPeg7ekrPvKOuZPzJz/ifBPvsYY5xmsqy65c
d4tQnRw/djoz+OVOqcSZnuPSDaU5fC2FS4R004Urh8kv9Mrw/OuGcGCoX0r2ZRHi
TelFfRSz0Abkp0+eiZxvuxVUIIWUz+ITGKvNTbDGHRM19DLMMt+DlLypEiEVmrHK
J+qmojFxEjanNqLGVhr+4QJ7x9ysoWJeDjN5yyX+phSslyAYDJqHbcq/NNLDDDiV
MiDNJa0VCNgb1+2ai50NiYQjnnwAp1FFuAVQkHR2G2Yd6eR2W8lk80+W4ffyse9z
6iq9WQG8Db7UB+DySbqZPrg2185UEpKWwCBb9JenvNIzYXVa0OWSkqVyrrtjCW+8
VCpQp5+K1oDOY8e7ZsBpQYXUzFM5YSBNA6H/X+cpHhxK8WkcywPo7zh1nMtBl7yK
8WlnQ8mIIKVogt0ispOoIxrn5XrB4INj07S+KHJbrugFcRZYCx3JCG6KchcpZM8y
VIQYAFqxB5FrEJAAtfnryXLY7/2kbsMWQeymdus/hspD/ujmxGWc0xiWt/0eh8/+
LTq82UPg3DNUbFUNYhSNM3vA2Hms5zhr3cGalbMlvd25Gf0QYQtHgi6RmCI2m0oq
XfV8j2Bo8KZlLNn95W0oSqK0gWKUmprD7cnvB44NIXDWwXGZTBIuTO/iOMHJeD0/
YY/TOsKmmkGx+IpUR1R3wkOtbUggfxRIxFkoQ7VqizzesYthXQAF6VV1/y/B1pik
jH77ECn3h0EMkKreMARvUKEof5gdA1IBzEHmywmTpZA+JyBrqRfEpK3ufeeyea4T
gZb8JszsvoegAvntUIU19bWhzLy6HvKSLebroUmHJakHM8kwzyBsK2ma1Rv6MXWl
CwPchl/r4VsKXcJn1tMe/HiVLRAzx7K6fApMwU+2fE8c6ZfTpre6CSKzU52G2W7f
NdeYO1JfiSZJe+kvXJy+8z8+v7gRgR+jAI4bvtoIQEsIGC8Hpz/7SdWD3vfFKxF4
zj1+nwyTKyx5O2NHXKWe2ViHk6MjuzsZKXaHQmz+UIXu4CQbceK9YQZD3nC05rqa
xeUhAQSrmYCNHkNgvR8rUAH4hkLtdVjBUtsHdBXHioWc4EgqK1ElnWKDzgCKk6W0
K2X9jp077KbW539tshmiX4zVAk+ZpUADpKI5BHI6tYTIjPbQkUyqxFWfixz2qYQ+
cOj1jc8+6wZz+pm/4vh1zGOpHP25g/NlwWxOXXkAf2RWNZJRANUJ9I8wXpAunwTG
1NMBYo18VBlu6vHT57LZu9mE8WfG00tQOQaFhXMVQ8sS+5K4b1ciZQVIQpjHMFnR
rG0vZ+6BIsgR5/MfV8Sgm/N0kxw28kbepGzW2HQV/KUQEiDNTmgTH4LvNyT61gbM
J3pbV12686eAxEmnUwm1BI3tqKP0ZC/f6ScqR0xPee04Y9f6xF8cgMorWDFpCn+P
IDDCIHTzRi2sI/bTkE4m7zAnjX1NgYLBYbwW/baNgrU7iN0b7WLwHbyTg8JRTKHb
0lZKng+8BJNu4tfx1bopwGw6tO6hfwImKkApRHXFwbPjwL2QxF2V1ZRaftWi3tSX
EAhPepiWbggaZTZQuMub55Ll3usD9ZD44F4Cqh3/5P3e1Ahl+lQiSwvEuICur9vY
j8p+31VgSfROVDmRtUVAf6mpg5s5XpU95PRM+hesEbc2LyYzwhyf5NpiZ8AHp7jY
zYgZIyYq5NW66eoTTNFMynSHOAWM3SL0+OZrs//KUA0xElZdoNtdCRn+JmbWSYKP
kwgLjvFWDr7nYcHKh0ycm14u3a2zvIwN0lt9AHAUR0tro+VwN8iCwyUc/NXJ6LeG
mPr/B5CCo89tPhlRxrwmPUKUSuIw1zfcR7SDkVT1yxeKU3x4c2TSPsqDzLPUKTSY
U67ufsCsDY0ZlQ9gp5szmLYn2ws+Rk8EvtbH2QWFTi8jWgmPJfvo+i7mUZPByAOJ
bnwIJ3r6Vwt8cKec4dYysAjFqy72wnI1dSFJg3TwxsIsCgWaEEmL2qN+wNq9kUpU
fXGmL4wqO50rm+2P9tsYd3xMKXSl8mGSyORpgIiv46B3D6s9rdCpM9cyiT+be7nJ
DsR5YUEMcth5KB+LeiU7eRWd9p4bVXORWw4Oh7LpORz1AvOE22zsTT+XU8t0s+BO
1yalgi0UTTpXUbPVukU/mYiGuGgj5L412wMv+nPyy+rI6+xCZcVJ0mB2EACPKBSm
ea+vbu3ES5keI9xyz2M3bwudyeo4FTNc23pNifugx4ttZblFgp4YALlDy1eA3hTi
ppDSXOBncCQQ6du+JcoU292hUucROI56L8pOR09dGXSmtWfIVqXRPI8YXeVlphLo
H23SdmtVcdGnJdN3EaX5ruB7IngSVaIOqvIw1nJfkBR2SABOywTkJe6iZVSIXqsc
acZGUQxBkewZS6JO/9iwlkQdl9f0PU/boNfyU2OauQtkpSAYGXYFdCH/NvF7g0XC
tzGNEsUAHjC38GSAs+iAwpkVPIXclKvSXP3LvFyXQLetsNVY/RR+MU7ShNxMSugG
MkEEt9BnBKoWVHN2fwa1Miug6g+C7eXluCz9cuWB9XSMyQpkaqpS6ol91srxUKUm
BFNu/p5KMTfm9atkJn3dwUZKiI1Qk2LHZANri/9v4Y4yeF3hK2z8K9HTe50cUxzU
WjzaPE8uAeEyf2MI021Qvwh84bazqNcqVAZiUQaD/bEvtxLtWx0v3BjFjeFn0mxC
bpOGRuc1kvmMY6shqZ2AmFSSmC7sSm3O8PaCmeM4fWnFLitA+z+HhqaZ2uDdWdZK
0WHICPTNQO3TSjHHNYI1jhykAzP9LDFkFSRbpjHTJwiUah/QrClmbVui4MRMY8et
VS4RHsO93NKQD7Thj6H89Kjpq28Qw6XLcWbzQwFVlJb5EKiBnYrZogCPwGmZ+++o
OWbR22K0fC7gyXno0tssThosxSjDU2qmUCKdlM7iOPlfDlSqxJvlekaHhPFkOCkp
kF0Q7wEufb3I5Y3uAEPUtKoJ4RftLhUNLC9rnmjT6yVMGlkLjArrMMIqVtaDwfHY
d6sRwdJupXyKOWj5fuNQyz7zde8YNO/J8IR3seoy53LLcat+e6rUg64Zdq1pjwUi
d67za/bCTZWUJQeajbOKjYDMxpQOZuinbSj0zNUApQYK59qXo4nZHF72yj3s9gtH
ia/eOnIMALM/oJchpYGLfD8OX7dj/bGAO0fWU8YiAU8gcpeOb21khOclyWhK7p+M
gBrRfKs01wVO3aBn7twOdsclh2YTRPpNr0c+4psgsvfXDEn1YKSz9ddYX3L+Z3Ed
HZhjGMO/noAuWlin/zEU6/n6EjRYoh8wrPGRUY7t4iLfh6h04pm6SOOL4l4WjLfu
VSGZ4KuPl1PLCdtd8Da1a+EjcbE1elaCItlyJTGF4hVVt0Y/ZZnm84KPWRfewZQC
Z0T4Izl7ouU8OLcNWoX4Qwi3BBoZalYEWpSymRwZUSJDDj0N7aRXWaYxDzzRD6qR
mofvQhFQAT1shF0oB34STtOeq6e6s6QMSMf+baB6dc0jFjwypzYQYl5kbdmTqLFf
CIpHpUTWgg7GzHF/vLpKwXUTCVPoVzvjJVR+lpQ979oAl5QrmP4U0dzSm3n7moIn
8uhVL5BMja+qbw6QCV8hXcaDl9mApNIaON2WX6Lvqp1NvOpJyXMXR6RV/1AvdATI
dqf4OqWDsdK4We+1kaTWsqw73UdkOsSnmSmy/+c8U7y0kV07wF2fp1/Sc56f3kBP
H6/mvCK4W6Bb1b9kXIEssk9tPaaXVsa5jHv5rTDVo0Jm2t7ARsOmwcp6rRg0vuul
WqzAfZYfzJBMyirCeLZwX9GiZPdpwI59YRS9//NZtBOD8uXcEU3a5HvPFuv/aayo
k8qegDXayFpkd64I+Adh4/CxOwsJtz7rXU/AMe0esFCTTTTRm0tpcdCLyAVspPe6
aZRoFIHiI5XNEu8n34dS9P4LUSXR96MmdyuLrA7WzBsHNoGCk5VwHakZWUsTe4q2
aGgcTsLsFZBwYnocFP+gGitJKg21JPAcNT66rxqFIit19Qw/h7pHgxv5YdZ6/ih1
fpvNy4YKWZLGX8eWckghzwtfCRkNcD9P84eR6YW8KZEMqlZsTnPlS2ziqJYzeGWO
ymmB5VJx+f3QBMaKDTSde+E5Sp17odWNQl3QiYNTDfIaoKbux3KRv4Rmm0Lk9NIB
11FLHYPavBQmrIm0DhG/kToFeoy+KaJ3jCCAQfffQxyPiau0vyRAXT8si/xvfGzN
n5tRiCKwHaZBgi4nvdkzFth7FnwdlYjbfPjYF0ODZzGuQ2Jg+kMKCrbiTZ0ycEVu
N3Gp/4x4oupCYZSWFw8p0T8hvic37qXs3diVp6HjdPgA8rgZkweGOvHzYhRbkzIz
3H3b9oz452bKCecY58qLGI9g39yIlb4Hm75P/Jb0vJXynTHAQUwL74Ld0HbnLOFn
TFi+NJs6H7Rj/NVwptNbkLqTRIdTgbbs9k3uOipxx5fd1wNuBxo5P+Viu61QG0C+
vEGVU2cNDtnOZraiGGzZWAHeUqsvEwlTGREtepYfA6AzAM7YFJPLADvNzOWj3Iji
+Dc9nFs3w8lZ2NuwhbH4wzq2oByXJbIXTc2EvIkxOIi2ZfWs+Hnnl8suR/YsFonK
vBJkDoadDEt8yz5OkFKSTXtJUjmjBx7ihWZVEqFVJpCu5ZOkW1j0L80lP07U9JnY
HaEa2hXAOiWKtSxGZyA/Yn3bnBqciNPFU8EPtokn3lY5pmZRtMD/HY4fDp2BB++K
ogonefqVrKEPqISaK0PXgeTSmRTDhc1GAbFRgQAIkdHxhW7Ivq3gV92CO4k7q+UK
4kT/S0VDsjCdK6pJuA8NmlMbjp0eRyAJ3XhTTlohzALK2XDlKM+jiFdvdh2Lu5sW
WiNk9OzoEDvyCc/P1p3RsDQ+lWI8ht8Y1/hVbdHTu9Ot+70GFzwgo0IF3JktueY+
1xcl5g1QVZ4ITeYzk6mFA/JP2cQZ1vIibeMVW/BRk8NX6DsAOS3U1i+w3pKVwbOV
2HLjFKK5Bx5+B5xXhFPR5Er3LVkDrKR/ZjylfW9He4LSQ5XdwFNFpTPMRCE6ulkm
Kcyf0xOGVS5PKmoanUtOEwxMUIjUR40i1ce+chC5VwIE4KAJaaigrT6dVINWLRaU
3cF7FOAPbYxEbsZB4mCdB3pQBVAJdKvNTRbBWLlgbetfF/XfoFBFph2Un0FnNBD0
SbD9A3zK5oQovIjqTA7MWOBZP8l7p5ecrWl4vkD1W9rwNSFxUd/MwcaXrDiTBr8w
Awdv9gJTcnSlDOOuzOc74C21KhpuU59aksC5+0OunRTXmSD46gHClDKXQ3ZpDRha
pgj5AZTXFc7rsT/UU4FQ2XeWyfUHhPI03+iW4Gn2ddbeFPimMX8MGa3k8o+3lTDD
3ZtItEE8EjBD1iOQq5VKpjLQ+cAn3tL3FY+akE/AXLxgS9bUjKMdD7uuiualjB+q
l5PVv7TfqL4WgZ7l8OSHNv+8F9BV3F2vP2lhqiQxi/7irN/kRAuVTj38mYOGfa2B
6qXqn//NMLSM07KyPSa2EnN4KVZnbmPyIr7wyJRGDf8cQjZFCCZjCdZ7hydeS/75
H6+W3iqcQCTYRWB5fWAOwvBtcdgbZLZ52Qpp6nLQ8skLKv6bQxVyWRlMZdGHkSsY
2T7elICCEjwB/cHx3KkXf4kK6wxr7eEFXPH1hLfPsdaeb0T4J1xwHw9/VKnr+IXz
ctL2/eAgaBIayqxcxblelEdOSuQS+HxieBL6LT4FGJab3EO/VhXU/yokM7uQ8fms
ydVVYbZx+nU9RJwAZbTRdYlMtHpNb0z0tOtDa06M+N04F+g6+5mZF3IvQfR+diwu
jWwiFPhEhKmUmqitbfT0r8ze4piiTHBErYqE4/ZFfHsX4FD5VfgzFyI1TplitS5g
YWws9hPN0OeH5a30RW3zLQvxeFrm5ihmp2CcXAaB7RdR8lKYUWUd7tFX0tKDBYvb
gCBwrcgkb7gFpi3lrMW2Q2UZXx8YjaOP403lP90W7A+wF3dnLJQFoG3lbfsPbRIK
JluV2lpjCBIgMlfeDDyEp50HWHq/DHI3PR3GFcPd77DA62rYI55/UmA85CmRDl2P
1bWvhH/2E3SlpeVrw5bw89x1fy9EHOJb2VvGeevzRzV0T8sr62wjgSMMvsaRJD0C
m6g1xL0RimHfmiA2tKbDwv1/zHm3QCONOAAg5A1tI7RNL9djivdpZUuDnKh6UBn7
G/7vkJRNtur5nBAmTVwq5ewMx4yZisCtAl44xJZ708bTWKcXAngAxcMcu7R+2s9T
1JDJq3+lFEYLKEzmzpMK9XylWsItZEkCLKDVybVRUAXj22BVyh+NfPWZ0Up2aNkr
IwhYUzSQD+Z3VcaUzQdwi9DBxywmLHEcCTM60BoHc24QrrzquSS/+91FNi+FOcOi
5dBo77g1ikFHUQCxpSQIuASla0WDUwY5G0X9jk77RpF2aYhvPjY1DFE1KMPi3W2v
Fk048CJJnlGNVehc14gkjxq2JRlIY1vTQI47Ym2FYHXGfCuSfNQuULSoYHLPFq76
yUOOZEGajyE5hBFXQPrJeOhqzQnUxfy7OhwxUoeYIU0FsSA3ZxZ3x0o83py3/sFY
aj4lZvFNg9PKyZOdI2/LsGANlw31cw8fEq9Q4ltYZ86E2LbW0fafNmpoucxclwZS
9XkDptMdL0BFy+sMcy3BaAYe5zRDeCHQpYqRiXH5sKwVT2pJru39GyascxhvEzUB
5p3MPUtHccKInvATBQNr0CdXusoMfFMO2U3X8WuzdNKz8DXgkNjFryNizgdnoG9m
AzCcTShCcA/Z/lsA4ll7+1AQjELo5KpU7zgYabbn6fuhxTTfBf3aCE9RizTQi/QJ
BIu9rKVoZN7kxbSnnTG3ILEFfI6UIY2fz8tYfKTS3NS8S04PKYimhu8J+ggVHKsV
kpRlA2BR0FJZHe5FlExs8Smkly4OYLKZxo1bTxCs14C1k/xDF/oZxFpvldYmCn10
0vJoJBE8OjGHBlWVjysntnktmaolWsfaYBFrakUU1ihnDkulRG/zy4JKiAdFfi1a
hKSsCiBecnk6liMt1PE969k1zpcyJrkBMjfnAomTLhbaB6uK9K51rPtF/n+Nq0Km
0FMoQf8IfH6/LBX2rxyBOoSqLhwxi0ZO9t6yL8uLyX0Me1h0TFtlmwYR6hqwy7NM
1ujL3IM+r4FoFb2+iRw6Qt2X+uEws634t9GQqHA435adzfytYywez3ouQKFI+5zs
cA3hUCM/5fM/cXtqDHNz4TwQ4aM9hY4RvulprdU4agl+w3bKH5xYvcORbgF+KWee
GdUczO3ZZp1sAEsh71z+wiEPBSM/7Dmsw3LLFsrGeFpoYUkIhljE1xGcb9psKXC9
P+7o5I9KIRD68xg/AN1nZTPVQedQztwI4hcbJFvaRjL6sUgefBygsY88hYEh2lrp
EfK1LLtleLfJhR5RyT+xM3Qun91ukqKgjyxsfcJudxfMj67sZyNF2pB+SdEdhxpv
1uj1BBqHYggoTmhaYWwin79BEKAxEMEZv/0c7doTz46LGG0Hp5RU1TVIrVjQhh/1
CnqAwYW4m+gkbxHXZTphEirqhgfSn2i+5Ynktwoeu1+ec+DEh6gtvOnpGPo4zkdv
rzZnM3c42S10AGnYR335P+0YOhJvjtMWP10eVqPj3H5Ovl3pjFlv87p974y2k/EW
7KB0diPZ4Xx4iNSsVH/j/+U3y6CVDd+32VH69p+8aFC3t4Wu5HZUEwa/3UKBI1X/
w4rX7GN1cCp9H/Vk90T1QvYMt9NscMAqQ+GnNVMPb8cC/0azKkF+rpG+wkbTfNgj
GkbRYI+h4X56dT7xzzELkWZYu8LgWqnJEw5LASWLyFAFMrn/mHitq6MM2tkZr31A
FTCVHqTFgUKGheaQv7PtV+RmBueGhG0yzeF+lhDD6CKpkpbTSVDY+ShdBfcJsFdp
0f85gbkHtmKAq0nsc+A0935zfkLjNukspB8XssdWQM9UyAWScCQybA8NARsci+I8
bEX3vBtYWsAYaTPLHPySC9JWksnsP+ALjGJOd69edzorXo7Yq1GWnLqao93gyj0c
FszhAilur0VezeV+Kx9KXdmdBB6Og7SIOn62lyN5bIvHGt6v9ZfUMBIy19CYZvRk
+FvwS9WhURi5smP7LUhvCXZPyKUVKppbqwQJKktEBgMvKRNKUi+D0cLxKhQgfIcp
HEXNzhvlK3gzez6HL/pngt59qfWYrgk4E0pjvIXgcAQED7ja8ei64DSTGvCS1q3m
97wzn1omUa0FA7JB4TBmmNxnv4CjzkHVDZgoxoZGTu8HKjUcWVVzDHy0+5lpVQO+
No4vPJ5nTKAgMTM7DwCYlaZimTUxWqdAzs9WqFiCdisgKwmV1em9oelQNCc/JScm
94WIuW2kauw9l6uorcYeoz//AJuwYAQjhj5og7sHQLFRDx3mSs+LZ1cPHfiIMvgF
CqtjL3cvBcTY+XCQa0vkIw60sKe7XcWSWsUod9vuym9AydZwBe6zaeG6AEK/1uFm
4UNIKOx94Mlk7e1d+bGzIb3lc5a68RdtHNEeif3zLw8bqKakliFy60+wkHwuGUZP
8INdTiunISR6YPX8Ejez7j0Ca0pdHUTqnzASdWJUu3lOGU6eIoIsnUSvLX+AYOWf
JLqxZDuuuLrFPXX80EcYpv26W4T2vgr7TxvGfNC1xMgDVmY/37dx+IgJ81S979E1
1BQmtJwZELX61Mps3+b/gTEjZoQlfBtnDyMcEHxEVTEsyTDuFyqZM/dBhScJq3Re
A5s/tkRv4qgfsYXhzadoXlmLxJfyhSMqHC37zR+jwXvyB0oBTnZblDjkPDw3Czli
8a3xklW9/seP4WtO7/Qu/rq367IV55WXzJziEFeFRkTjFn/2RQAIUaNCZWwM/LTt
c9ZbtOpTrMrjrPh7q3+tRulfQtnqWdgW6B9solK5Wkhdh4aUPiimlqOi9E0csldj
PZnt92/o/q1lO9/3QFTEvwp++nfnBpzIqwbj/Zacs/CyV2FVBC1fmup9rW0UQOiH
et66n+EOBPM/X+jni+WNUOtt+ucsqZhdgZOdeiJa1Z6p4ftIhvc0bXEQDKFU4ESN
LEkNGFNhwPbK1FGO6sFafLvn1S+IJUkCWq3BaLSpJbL68S/XNPm96Zaky6XmnWbK
PEOv9ew2SdhyM6XQxZZBZWA8MFC+181JXww2JZXhM6J4nbj8XFTw65xFZlZz3ZMA
cK0D4bWtSdnP6/fBq1evrPoe/81RzhDEip81JP4dqAeKdKrqVTgyNzVLptJOJ7b4
e6bCTewozz81JPdCDIb6RbHCHhtP+NoA/SEO1pvppPp4/OkWgKN38M/hWGv35fN+
5pppXEdeQ4GFhukJGZXZEKI/ijfEIAvvcb/TdmohxI1yXIYQhHM6mjU3ReUQxGWR
RmPZvYd4v3p8svWmdJYz4r25FsDZf7WY7z0MuR6XtB6PZ09NWl7zvk6GWOGWAa4p
cv0TDs/jtjmWUrp+M+iF+FYtTbBbOt5BASZnpQfdWWQqgwnqq/1Ob9kcCDgekQEV
TIqzcL0k2B2rY1gsd9NmbFtddir6mWoyVLI2lvlugG6H6IVXpuD9BRjYaukyj/dg
H1CXEfjHLsibxNW37GUslDUvgL7lcnED0AvbURoENnwWB2iGj+HI4HPZqvgxCV75
dzqIEREBnKZNfM32BivZxT/kEH5bwCGbnNc8IQL1LZcL3QkcQ5XN185Jc4+AC2/I
bDzIzVdyz8aeiyIAklHWu0eR6QcQPap6qHC6AY7CIUNaQb3+py6/EjOILwmdFojS
c95ZczlGCU4qtVFzBnEYZNZnc5tRXg4scnCIEFQ0lArU0SV/zRScXaRnTNmnInXK
18zaS7aSepvY6/xnepHRJZi4Rxupl6Ddp7shLtHz6z1kfMtl6fd505ZvN1xB5Asv
y1vha/FAypXM2AgJAOu0VDYIyRcaTyvhzDHhmt0N/eNZ71FXSoqReOJxpVIo0Xnk
9u60/joHE/BtqEjaQpGNMFFyZGNrpj+MuKtVTcE2WEWxocB4PpG/JComIdpxGrb7
X5hx93wXOHDABlRuDO8nE/368/PjDVV5HIYLduOUNoNvVwByFKLL7Rp4HkLHGDrY
+HAt2haRYMtpmdmUrvviTzMKxIfg0+ew7oHRM4hN2kLRc1dn3gqg+3OaG7KdIB7z
tUL04b07NhhAfYuAL1aIGVwFUen65q16a7Pus5AirdRtGeS9lv39vjh9g1sESVSr
vq1LwXBggT9jqCE1NBLONv8ilnzkg6ABIlbDkitPdCwDc56k4PyhmcXeTMLuZHkY
LqrzQTL8H6Bx4GI9r2toK1c8FPgikl3V9W36OKLSlTJjdst1I4PJL9ssla4mM+6x
JzMu1utSN8mqYEaVtARGABXXV6vrG6oq8g2Yr2ThWJPIy3/wQGWO+PyTNJcSRm85
4jmpMoI7aduf3zjW7tmOY6ABOFOhd1h1ikgLlW3tUgtlbBtVYdUoSeVQZbpqLcKU
xcV0C8nsOOSEW1WswSY0Rnq/F0Z9ESm5hoWHhE6TDphcLGoa5W2QH0UT1xKT0L3z
PXHVt5Xi5IETWFGaoJsxUfJe8PUXrXCmSQ45ONR/YouyDI8uYbWxhDkY0N6W0+eq
hJQx8hZXQPs6Sy9kpu5BvR4S2wUYPQkvmB7NHOCh1Pq25GrvsUIZ2DxSXRjJGyek
V8OMWrbPs3cB0jmBFA/ue2zjtAnTqJmUUPka9y0xoFGxILiF8uxaEo6NfNbWF0ci
q4sHJbbotlUonOQEP17c6sPyhkrS9OBAPvVZE6B+FmjluX3W7Lrark7DKRVrpqs0
DUXIRrUBs/idaSCCsYo28fuj371/L24UWr26PN5AP2zDQB5c8vIfN4NKvFNn30DT
8rpezavsanq9gZDlzdeN4r1MzvX1jZhsgUQh4ttv89jJ/vqaqIH+2ARAygXmcB0R
L+doYUuWzhUptBC5VhUVhm62odyWJXVrknvftH4UhtATHSXt+bhG4Tvl8AoQo5FG
WxK7TF4HqkWise2/Odtjmwfn02XCAn9vn6rYpHPKeoPqhwWADwHig6Uph3Pqusl/
trebYqm+1plKZx6CmfOP4Othzn6WJJJIFZwOtvvZ+EwOwDnNC7jnu3uS9z4Qgf7u
vrIwgKs8zIKA2E5tRQW4IMMF2Gj4SGvXBeEBusB+BG/GHH8WOTZRjNvNao6HFnvE
t8NneV6X6Nn4Pb4SCqcOEn6LwXg9t8BFiSxwps1e/aBX/tsXolZjjqGsXJ1Qsufv
Q0Xh1/vEK/QI48pcqub71YeXL6Twt8WhT8PS7pUSSKlw+IPRZU8TVobkMJf6lvMn
DFCTZ5Q7gtIfQTjYmrtsuPsurw2MArlhqZpaAf2KUfaqyzx+50KYEOL9Nvm2G12F
hzcGisEQJ1ODPK/wAAEhf5LwAN4Df3c7FTGsvVPoocqtCcGv1FmJ5AiDu5+tuoGX
6a0vJatLwQvm/s5AUCBnezXykDz93YYPTohJ2J7GizAG4yzJ8aI2SqjuDMyP1fUg
5nsp4yEbWUrJKyjk4Goc/Tm/MOZXOnVBfDjEzlhomTU/OzYoZhKDxnTyF46E7sLi
aU2OWwZ4PNpRwGfPjw02N0ziQ8beV9j22Z+K/ECFh2bvV39zLpvu4TIDdNVE1O/n
Phh5x9aKHOh3TTiDdqcmhxaBgwotvsk1e39U9sOXrMnD/BIeqrkpp85c3hqSmnU9
ZhIwROsK8WE8krzNuCOcM81GCNBwVUf43TBi6dNj0T1xR/pOfs6a1Zd/YBs0CO6L
EsGWVjD9Mn1/7UFmIP/s39NRe6DMmIpOzgUYjpXjd9KHk6XHzoywv+aq7bCQI+lr
Q9Dlk8wLL6qzzQPXexqiCn66MYpaSgzwaJHuwObpl+hQg8dVlBfnwRXXQ4o929Bk
UvTSl5bmTNEAPtOEMXXnKch+qVEAEHW1ejjIVXzT22KPmERmAZtASsI0n/nWzv62
X8w/zzIAURZD/eHdugA1niAtS1YJqHp+0cNOFNTQubUUcS8xiXDUsHOJcyZMVVLV
uF04r5kHxAQOSOUAipjkQMoioHGXKC+wgIv6v17/kjVS36xeXJhjLoSt+J2r67S4
Ry1syuaBH9DQLH4s9IMPyz0J/QTfO/r+jBskTXLGHT+sSp740VFN1vV9Zv+0S9gb
VJAteIUQhpbfdBfVw8F9zT7KE8fIZ4HU3LDxPZJHO4JqQaEUJDciEpY6iYbm0dSb
2W7Dw/Ph66iVNRgsh0JsWtg7YcVsmPubxX1q6wNi/TSA2qF2zilrqW7L0oiEza9m
5SpUNbv9A3Zq5IFNiPmX8opXEeXbL6Cji5UXRTVbV6cKseEeCWf2lQ5drAxInQLu
7M+BAhFs2+rljSr2Zi7GTqlHsXL4q4Z6EXh+TEzy9z3W0tyRJ7D+P2awZj25lbEm
93cPrnEDFDlDG/93cau79wcKCfIVEr4qpW9vO2UzymcQPg1HIjuIyE29SN6Pm7WS
rsAh+Em2qkUPLExULjgxr4Udbl/0rYi5uL2D1RhJ+ulR2MP1oMjgoKM+e0U57k0X
9mlw6ivZyjDhzhDrJT0r0ihFAqeuaPfj2/8els1ieyE2RXkYZjY8Uo2u2tfYJvAD
yTldEk8jxWpKXiVRXL9f1aZZ3I8X7S9/9xMpkPqOc3KtM9mf+4xMIPrXgBY0Lzb+
zhiyVPV7PxPT9lgJbxpsNtJY2dwi7xtgvx9wiRL8IH3Gjwx3+suZTzhWGJpvv0TS
7qWh2012akXk4ChCwTm1929TeuLo9nUkRpndVYAvJI+Um1CJzPSq+HMLrQH3505r
G5NIX2jigJ42qNKAfhO6GXsMwD7ppRhl9IVVSSiUfh6Jl+91r1k9gCb3CTAVpUus
/HmuUuqSFM3KKMU14Y0VOwQdpXBNnR7U+Tm2YTWfcT3DjEghDnlpV7fKEsjIJFmW
+Etp5hiuD7YKP3NNpWlQcTVGYbSrOJU6GaAZ/q1zdRD9BazxJqPGgRgpKkFt2Wty
2TtPNIPxh/z6ZAkMGhxkhiAl2/pwwIMpPyuap2L75cnfVNFF2uboELcjHIPxrrL6
WwhBRfQmm6NVTeAZDQ2fIW574k9isesBWzD1ba/OlQea9EKgmFqFR/Gf8IDSZpRK
uU23H0fi13sfjZgyqPbDXI1gN+r9jLygLa6wqDrtw6vUqHAP/6nwQaQ943pLK2k2
iYInIPCCoCZd8pmVAhkT3uvhvpk7EyXhP3NOIZLIG1TAOThvpC6h4jjiuRpLt7/v
btfnfV+CSYkv4zwAQszWEH4CGWxOfZlKAuHqh0cfn8ywXosKy7QAgV8VYvaUR+Mk
AloAzGTTpKYE+4hqM6p5JOqHA+qlpNGXqiP/KkCywLjFMw9Vz5YyoSVLFnlgpI0x
KHGOfn7BWewaOpBDnj/bt38rVTYNDKIVbUauG7f2kL8wZyAspa70lv4crLIaRgeH
io/XP46axBxqrVPrB3x0Vu8ddAVx6+4PvRjh7cA2E0RkwazHH5FCi8pwEebjHwCd
rYcSRiReTics3ZpZhYoM7J8G+beoMK9PqHO3fw0guCfeH1ZTemvFZeHxil1u78B6
7XAD83AzvsMVvSXs+db71OInoFZGFU4Aky8UXIrUj7YvL2AMdZVvTAFRTvJmzQnM
wdgTORlApXbFOfFo5hlBcvSU3JiLdapMVKPi1A1GpgOSEZiXbl5vsB2K0R3+gSs5
hkZtQzAANGZiMERIqKQWb1EJa03sqsZO3UKjSI2n8OvJbneRA91ejSeFuM8nYYuI
oNGR7ZQiaEADE6CpvvZjmkJEsGDL91NW5nk0KSdGZPyzR0RAjbjeJ+k6ce08by45
aJ61sDZQnIKdAP7GQIHNJXY2Kzypp8bwXOqvYE4qyFzY+KBHG8atp43VtKTrT4gp
G+vVqVNSu9t9e0v0bYvqudlQ6Odz4b2umxBrOAeOcNIRv7xPe81YINKQ0Pkk+a6z
sjyuYtvT1AsMdr+dPcAgZjTO6m2D7Gg7KAhn/zZKD58lc6+dSL6gHBHJHzt1+Bon
AcE3E4HUMJ2G30NW9dVP6I7aQcaWf/VjMib3pR5oIm1Kf3e6eqXLCAk3GADSwyOD
nZAj0a/D3AnYXn9tG+C7/blMQpa779SGTloDdRHT8Vb22SSkEZwOrFTghklGuTDF
qiaFvfgXMjvdXKok5PYBQ/MK8JVBdBuQveuk277l2bgl7HMZHmoO53hJ0Eg/GHCw
D5f4ugeiW2PQNYOz5UYxgO0ohPmlxs+ihp26X4nSNHn2RvlHKb1zsH1VjZQqlSkG
ZHIRaV+akXxDxzqEQU7kLECIzDt9n+YukKr27uqL5zF3bXeRcQZ30xxfqyvDc7eV
ua15NNvNFEPd1m59Aas9caesZNDiZsJMg3k9605En3PfZu3W3V1k1gPU8OTXhjcW
PhRftyiOB0R2t7XjaCLczYHF0LXGTLMqI8bOwH5GAtDryrQVpWeJmAoFujh19Rl2
+y+XVcsPd3N7TLTM9BOLmiBcOCT2UvZrSKaS9rMtlWDdDgcoRP2fZ7U6z3Ojmrwz
ntY0tJnagM8euyW348JwoSB+XqKfG5aJlkvr0tBTBk4CcZlDSPk+otnvv2a1VNzk
wbVd6+eSfXPziNPyztmq9gX2kDwJCWL8k1mOlc2Xfk0oeWNsfcPBcN5FxUikKjVn
eMX1wukInywrcbhx98WskVQ9jQpQL4ZwjKBLFLdaknCjN4zZvzRlVQt3HZAz+KPo
l+5AsUJ2xnqVP31ERedzhM+egxeQIQHGWBdEwkDhuLHgKNV1Y1gpjhhxzilvzYYp
kjVJuPUupDibDYGVKIHnHa0R+PX0otfGYNeVkoe9jtjsIa+ZbsjhcM/ksASemHtF
1qLPcil2/1vpKT5dvFYprPWBOgzvgJhF7d1ZSOVDY2FnvjuONneSYzh0IQb2Up4H
cV/exloiEtqFYZKHMTjvv4KLomKQGMqG+umLqo+Uok6XVlBM+7rpo+fDZezKCBKQ
3H8DrMA/kE/UcxIM4/DhIM0+3y0SGcrW7yydM0+MayLNXrV4E1vTcLfSCVbg95gh
fSZnfR8N7s1TtR4D7VXZBlJ8kTgKhLaO7udHQuO13vz6K69nJF3opdA8oTk10aJg
HYHtPPZbyDhAOoNGFbcMq8Q8vI7hT+NDzfld9GTaA4iMHg2BhvtGIUazXbBcDkav
7CvCB4cUguy903S+s4NuBOexbOwlSeOnIH0LxAsSK2TO7ra4C4n2luz66YzUGo4Z
efzjr0544rGSFULnEQbWqN5s9Blnl3ONGqDBBEEoYvdG5kPmmcXCCrDM5FUigj/K
LjKX4AwsDLdStmK4TECVuwLaK6KaVJgeIpjVSiW1cWqpmChJQ24DqC9K2T6+7Ir3
XhgINjdd3LHaImu34GIW5ThE91ckQ7A6oAYMT/jZe3hmORWVdFyr9oY3awsYpBMJ
ngFW5URNAxGNHUkW/fSBFDaMg2uAXn0hDMJuPBzr9FUiuKhU282b7lqam0GmJJ7j
8/f2omCltVoTFyDfLtvtsBECLZzdto2ccIvsGfAh2l6DKTumlOP3Qg5rlt5LHq0z
InhufgpoH/wxBcK6oL9hW9BXlDzox5Ai/kRZCkkfrv4M3uxrk42ZK4mhUm3qB8JN
YhlU6CPRmYlM0mpe3tc1C3DHPqO1cbLkTvgfOHtwn9HXibCASlVOWG4zOuuaUFK+
KmrI2LKqs3kInCrMfS3tSCwmMAjwMqeC5O+mFPqw8fWopxPxbL4Cs7XfZ+mOYwWK
fOHj365/y3q8XUzNKteBNSYnUzqda2nu2Ig9Q8Rvi745UuakBGeZr2XimWsJgpAk
0ioo5n7Pehq7BUJOKjf0X7WKhP80jeylPp4CVtEQEhYGNcx83BiH2v0CQsE0drOk
/EoDrmHXLUnw2i3falo1NW5vHdyp/58hGyxxexkQv9Cv+oG0z1HlsS+5G5lrrsPT
B5D4LI+vvkShoDykgZYcOSvK4us5/ooHB/JZZVNFx8ybmzjdJPQH2GYWSe3unIGJ
NxgcbeBWINzK2mzqcLVX30TO0t3dNUFs7unx3+5jV1kY2/08hMUDH8JnenbdpSlG
REkB0Ofwvz/5MJ0S6XkOOBhbpFMzNkJe6T3GKuNrArkKpQV17zcYOSB1v6bhULd8
XG4+I+6AmYa3bJ9qrdmZxkEyeOqwnm94CHl3symBk/zylD8mj30KtYLLbx6CVl1m
adL8T5S3E/rOaSRwYxXMW5oORI11DYxOxOQxgNn+omi0Iwq1SDUe9i1js8zq9Z9P
M32NPM0U9NTZv7r5ZRhTMHKnsVwxJBJ8kQLGEHl3E43c9929ADSPDSBOP7L8WAGa
gQKKmZeqSD0ArC8qpEywaNNK0XWoe0VdhDBvOhJW8T6K1YvX/v8YUcnsCqQs4ggR
iqyonU+IxCQECYV6B90VM46BnFpsHSWqMEPTZmYA8YKG58OZ05g4sXfYNl1NhZyD
44Mvz4a2ACO2o9Zdtwl8+US6OoJKlE0K7nCtScdr60MbHiSgwhSQxPm4HF2MAZSc
O7oeyAp6FSW4+Ctjp8tyLnfvw1y3ZCsQ1vuqdFiLW/EiGJ6RgqgOKrs2cYMeeOod
0inct7REjSie/EVMYaqQlzmrjkTaqghdxlcR7JHyONqaDlgyDdQyqWj4ItMX4Xr6
GnnXdXpQjBBk17YZSQL5zIGi4HhU2yh+/sFVR5NPiil6io06DA3FMptkZVsXvLyG
DvPufcVwmgRVBBJhbLBS0DOcekgbybtrJN2VSq546cnWM5eIOOJ6GiPVnSBu0HyN
TDTmt5ZoitOiNuCpjMV3zoNDBQIAFHtmw9LuYmpwgbup9OmdaWx7FpPTnINdol9A
hkPbdj+C7ZTXTpAZ+RsY52Afox9q2xi+SEe2xWSwvGpgl5SGESC85YbD6ZjNXfLy
gg6GXVjrEGCAvNHK+xp52APL6BzvnWErfQyGTDzXVTlD47nOjTiwjZAGdZHGGJxE
ItBFV+WWPs2fn6WUi9enDeG84VVy+s3TPFLhn0ThUTveavepJ6jhgHt8LTEJs0fl
yXtjdQHNBiNePCIWgSAJ8R26brf5jqVlzwR9XITGPBvxzzVdojx3HiXkfO+dO6Mk
HZ+qEHArSdrEBZHUm/LjkBSCM72B3LNLnkyRWe0bgUMlSPEhXPxEmDPM7HlMyo+d
RIpHpAG5Hk34ITdY7dc8SvO/I73ED7qmePHQLPKwdFIzpBtOXcgV2zm/uE98p7iA
bbMZsAbFh7WZvZMi0+JdrCCkQwSb60zJnRuXdU97DQX+07EdQlULQQtuKo2zkl8V
kYs+BLTXYYMsTl4ZnipCw9VSh4X+UF73bQFdY0ufBGqkduJ4nMNXMrqfLzp7rrt4
kL/AC7FoAaV+V+EEJuExNQ+f0BX0aSXqHzryIpvOWZSCLFgbIWfSNObbo4MvPDVo
1J1R02m8gb600k+yiFb81NecN8oUrBm2IToUZara+JqPoAZptfEyB0CoKGfgK7Oy
1AnT0M7+EEk+1GYpVteeKtOvQfrJd4HUesFGTPX/KU/AZ7xsgxoUmVHTf8PcuiST
UlyNioxIBACAXkayFUa1+Piwc1KVOwQHWtXnHxtV9bOFq33DFq8dDxAzpiFfNyuk
onKkHwbb/AmSTO/i/CFo8LJ2NCgvy6uCpRa39a5wJ5jBTPeShq80Kaj8gVyVE0Js
epl5RZpBzDaWSVjl9Zp3hBJnqg5vq/mQ9x8hfhL3Ix2oN4RSYgsXQzQuk45uVz85
U5LayFzoJGkNjmdBsN2viGZA/JjeZRauZa63WMpPRpp7mgFlxWxnIeLXVDpyLcbc
y9/KBeqfoh6UYnpv50mCTvaeyN1vYKxXSQQE+wpjB/1zJD2/pBuNa35iedYldd88
saK5OJAueumC5dzAkH3ml9r2lTCmuuG0bHOdUiWTYFvDjWZQnDZ79V06KCf7UoYt
SxTdtqi6mUGEkW6pv4PQTCU5jFvnTOS7XHSKpBv2TOO+cvxBxPNJ9vUI4Y06DCdX
IXE1fnnzgFzPCO/hDE/k5j9gpO4JqV3QCjNvkF/Vaj88Fu1sCecbZizVwJ5VaSDr
NDzZLtMsMKV9qAUpBdVgZF2U9PrevGKBPrEuEr7JDtM5frGbcAtGj2uuDbIGSXgA
bquDR7d8plLBOxwQZbH02W9yvqNDgoyaCRf8eXKCKDEPPNvPxN22ZW0ffGaEsw0C
AUhKhRuzDvLL76ej7GcaVk7oNTfOG6cU1ko+GILIowQ/aejGmi3awXAAfej1piMd
vcrY4jgK+14LDKKFW5PPdQw8ajiglTGbx9xk5WSTXq6cmF/7Y2EH3CES9ngiNpXP
LUR2MmB5sUHMechmFsyqT/1kRFDQ4dfArDtAssMSzi2WIgta7z+og7om3BMZ0eO7
AVqDQp3tYVGz4roolNgLKyDs11SNpbFPaiAlfkP+9kO+w+Xlkhg/8nARYNsJvudc
ObsgWk/1Ydld/HpUE1tA7M9rMXvkNrlJ+aqldeCJ/zVPHGECxOSs0Dc7++l5cGbu
RQHcwUitWZoWt/xBUtXXPhdaqjNEZ5ZDB4QUKKC9GF3i0J2KTKKi4mFTUJkq1hrS
l77HuC9mraSw8BQs+3dOjRqS9eEJEuO/VbiPc6vO2Hj8kMM/g99NMkNs1S0AD9KX
i1LK6f/58/8vHZg+43Y9E3KytVMmugFCy0d8eZdRA+IpRT2MNDUCBgsHa95UgxWZ
E6li7a6cSkg/fGqBaYY+uXCpEI7wofykrav/Vb+suL/jiZ43WEVWECzWYvMw7Gmh
iFKQmfVsyXM862QNRbW6myDAa88h82cMsZQ2oV8msC5O8QKX/XGPFF5O2gUrLDK+
Yocbdr45LbRQX0Pcnuh/LjsdSne4pX7U61t195+JBav+vDRSzKM9TekOvNSH7x0F
E7gpsXknNp8py1y0mYFhyG1ioaG5KvfiDwlMf8DAj55tP81LuCmoXz1wViFup6Hm
ikToS6K7sYtiF6Fvg076zXCe4GzxysN7hC7XsL/80JteuVKS2CCGl2UqBG08jXYT
DSDSqkLD2cd41p8NBrX0xCZqFSiCXLLUVPAw6316g0mwvGN7uaLnmVW5OyO0LoaD
7OzW+gMrSBkVgcMfUBDy2JQGVEoYXw58D8inauevPu+bOiPH3gPYKYmi7NtJDlGM
judFhAvfvf4Ro/PmFg/9uI6YBGGvM/Ec5ERDgKYd8nHNr66iogHPTSfOfwHan1wf
eSPLQHADXz5rJvwBy424eMvIUqJbNRypEOLOpcRvEReB1brVyc17KXm+/4GoUrP+
FNbD4leip2nEuFA7sOJn/CAeIqlfTIQ16pEYP0V1yU/fI35bBdRSXm2oQ06PYpFv
w/if4aluLuHwkXENsiBrfG7CgwnBrAkSNv0qaPiRnmx9mO8KqEvlDIWMTm34Wwzx
xlcERArRwaxQ1kJk2aNKwU/UbPa8GsVtE0RJE+YT+uH8OTGpcr5vmw+UYbR7Imlm
honFSMGuscc8np7+PVmScFhQ3yjecE9QVC1sN3MtSh1Cz0AWHayTN9aqF+4f+aeR
PrcrqF5AFfzaMkah2w82MM9HRK9uKTYEhWMDRkSpsMyPj+lwZbyAKyR0iR55jYf8
DLp+KYNCLIV0RUMfG8f5SHQOKlF7af1LAWW/PW0fVmlYooP11D6H1aI7a4TgTSV0
a6ZcnvEpyHY5tNcWsLTvfOYXbkQEJIEbhx+eKJN5GLBpsawZJ1yHWE5P8NVxEZRX
BeyHHGynXB/G/SOE1audflZRfgmoAjIlzi02fdb/nsKIr/7X+XwRm1uej4orD9lD
v9Nph+Glyl7vIBf8KnI2dZQO39MurNOpXMaEs8fzxLADcSss3gN3j/2oor6W6oRv
7XP2f6d4CP6ez0+yHMuYPshZcSRr0mfQ0ADjhgsDi9A1HMgpG9Y0H3LpHADxleq/
KzwBQuLS/4NucDiicQmBolDwRyT3/c+fNSlrUdG+dMam2wav0BgMgH7Rmza3UPzX
F8AJ3e5CFI7U8ZhfbQUDopRuYvL72xVdZtc5zUhADWEHYSBYHJz8Ji++k4sR0ZMZ
LeI1bUjhYztAG5NGHTxvNbV5hX6mF+Zcsq5/iqXo3XnplTOeA4ys5YzJWFaDQvYD
QbHSZyTD6KR7sf5BMWV04kq6izPNao5yL7A9a8U39BfwCyybDT5EMn5IG6OV6NA/
R4mDWMUK660sNsuYwXBGGNWOCrdQTPXfftQkoOfzCTC14TDl/O7CWhJNxSVuOSAW
wlRi+HILoWO8r/YY8yiloniyC2DRykWw1jPCpL1puaCXTVbAB4OxL3n9rvLiM3xb
vKRgrS7ysd2vUidjWo57pHJwfyp4qQ9vzkYxAir/obtb4fhTPrl2eMOcY6ud7siF
pTdb1jrX1FoNloeC4afo3+kgAVtjyiFXmXgYmHkg71CuZYBoOVOLhI0gSuL5E1M6
JdwsqiKYex/+TpKT7ZUpcXQS8kqy4gkAXvSyVhar2//qHZuZa27HrWmRLMXis92M
809AURCgco8L2UwiN9s5RCQWets357uDp4Pvn7Dzxq0/DlQqrgnXFARKkF0O0Tb9
NeDp23+yLvCwFB58xn2OtypSZ3NIPg07G4qF6pUW9LwlC4BIA1y3xp3Rk9z/b/d0
Nfi6n9FGrwPK9TxHm/4/AexZPGfRJxlj6Xq+avbl+XaAOmBNQ6p4lPP2FRogNF2R
zoT3nF1k23leNZRndrbQqQ/4U+KuvEUbvzzjA4tPUEgKYxTBx4CCZDaCGJZcZDAB
VRDcU7DKfBJ125XMsISwmKgiYkNVL68P3h7BNRv9Ahq4wihOBh61+tkdNXlp260a
p6Y8gnaHBEQQowKJZ7igQdYm+ycZ99jFVeejT+6kOK3BgJ//1I8xjeIY3+1kBS1n
yelK9JiziXAgF5UuN6GVzNaKRLZQo16lq6SxzXFBXSuT/bkygyeL9uoELONG2qs+
8a05o94mGnF6mA68opWcVzzOlTo1Zo+PRv26jGVmckQLi3JYgDAvZBBPOLAhjruQ
/Y+5hJLdmyUlbuCTIZPhxbpdf0JBXfMvspdPggt0aJACQa1C2SXGtdy2AEGnPnXP
P9EUl5gVWqmb0pbCOkG1SEpbWNm23yU5cqijVySQxI1wuDCN0IH/164Sg94KzqO5
1d7UhTrU+Dd0GKHIy6nR6LJJCU5w+omKnVb2NivETkZAihg2duK71IhJhopQCvGL
yZTvaB7ACLLWpG+h8TV2wlZfP5n2q2lX4KLZsMhhkRreq14Rs6PIomRDzfxA56mD
gJcXipsVnqiUNwKyCuE7dvMwSaDa7916ZumzxrQCMMF2PtTeZ0a4b4/xZsAwOuE5
MgZqDO40NakNIeNdI7FHyA3xLy5ApcaVi0IMF99tPzp06DjoMKhvcOLMnAYfuF3D
z2dmJfepxwJyIqtXHeUvFifdIJ7m6aJuWyycT1XRVVanfSfaUk3p0I2eVwpcRHyG
V1+57HzMRh2hMkU7jbV8Hhj4j1KELyuAeKobRMfzcpblu4i4kR5Nj5zJngLYuxlz
RD4piQ0X1snYmiN/HZW62DzmN7Mw9VQN5k2LfxmKPNf7K9Urssv1OFuFZC6b3dUX
Ylzlkm+5kLIWme8jMsaqdAsKmFdUokQ3tjHo319K2f7fUYhPW86MsyOKdXSzrN05
edM8Sw1UIfrbEtajOKj+0WZ2YRxoIL7y6AJgddyLlimhCK7DFUb4n9aPY4+cTU14
et9G18ataEdW9CWWi2WQgFDPooaRVI91h+Xw7jF26J9KzV+Ggbb58tsWG6eDTDNq
Ujl8bwF4sdzcKlW5O78lRre0M3D6eSW0LiAZIKI0LTN7RreMxz9Uk4CLdCWm9Ygg
e4f+eVc1ea4RjGUXfA497LkVih053nKhu3UFWJx+PIwsbJP3doJpzNySEKchRGsa
mgZv3h52qq6aFMBbNscfvYds/BYit2Gn8MrzGYm0Up6cWmpgicAULJ/n1rQP0cb8
8lDzc+79005EH2q+13bMRVaKCgi6S24t4mc1dQhS8NddaMeki4QO1McNySvFygCZ
rTJ3Vt7TnWqH++Hva+Iynv5Uoq7HzR8qT46gHr7VUYJEcu9mOfC7LUusVHVshmam
qaWOFUdJB2mHpKwgiv5NBJTuMILD3oBEV3vkjUCyQINi7q4c5y3tWDPu62eR+seG
RhZw04lguly2ZI9SAOvV3zap5DkUQuR/3Sm6nsbPl9TjgxG/LaWqyvyyeeGhvjVT
ChsEHTZlVlPgtWtrmEFhm/McyKKtESdaMB6yxSlMh8CNiCCrMo1x8kgsrdgMfk3g
2eAtPMO4vJNt1UZEDeui41DBCPFhnxiU+prhyVFflQVhjxpPot5vSHeNwHFeKAoX
yKDcHxWtCuKphoKnFvfJ0qYRJ4e16GPyn2I0aZpAEvR4LGvX3hfkna7vwi9IXAvp
Ptunhq9KCMaM6s6kX0ZoXNG4Nt90mVAZnOvgUa9z1v5rHLTpEljprcEX8fU9Ilse
e9heVwvy0Xv301A0FiERL0Q+6nic4lF6PRItON462DQrUYWZdXga7C5bIhdQYNjg
qzaCxuxV0fHzCTy+7SAz3tt/1Vm/nECh/aDQpr1+JH6zZkB+d6Ic7U5HzSSD3dMu
oL8FbGUsI+ginCo7GxpIy8tOO3enkDg1VCI9P5O4EK3beM4zUJ5PT01LqEEroNaZ
EBGkwhh0j8EK61U9h+bcY1tBqLfSwlNbF/LmeNs8zDKWSdYE8D/cqZKpAAGVvbSe
pboo2djACfUWh7HJWQvSUXd+AWvmdcZ72AnJeQHKPDsU4cgpSzx2GpGaJ8lH76+n
hXcSYXXlQIXHXeJ/ngIPO5hEAtc7KnhM4rSBzzHETnrgl7KWL0IHsgoz6XqoKqgx
cWXRAMcCff2IRLXHIcx8sNFCUpIpcuOYxYiJ/JIT6lMKRz4w0K6WpZBFu5c2m//f
PTqMOTz6TlIddg4gFJxp3sprn04MgpdcYv/2Ivdyk/r3t5b9UKHqoHiqMcaTHK2Z
zxx1PH3r1n698bMv7arf1WuBWZwB27CosQgr/RufZj0ou/qv9LRcFwUVsH+ROYey
rbFImU4UqLw9GbBgCLdZUvQzoUmW++a9swpJ+SdhQVg8/qB6UvMRZytmfveWFcmv
pKFADZi/mFcGWUNCIZ+sGKwYJsaXQiBAFxpXWto40og1TTumgqqcaNlbMr1cRMGl
Wjj308GGNF515BjtmQ+yKXu4jtGN+1vthZ7R4eWGWZ6CSAC689E7w7yoWK5Xh4J/
AVhbZ3yv6yYMEG8mUAuBUW/zCSusAlYXvNArur7ETP17chwU28/13IKW4jujLmv9
0r/kvnA4IJh7Wd/Qxu8sMj+GxYdggNcuCp2YKKO4euEoM3jfcgovYOAOVFCijryy
KvkiPCW5HV5KmJdFStILEnD/ZfZKsMbMJd/lKBjcXFgJEAV+tFpc5flNKL1fpFPN
/kWRE4velf2QBjQi/jyZJL2fUIyjkdKgbBkB1UpdmryJRaMCPiT8dlujhlQ1qneB
Cc6GekKgqcl5Z9yLN4D6hkhk72ArvwpCwms9W0P1cBd+qrlizFN/uUx5ME001kFl
YKkKEdkIBCiBCQ/biZBXMoI9H4c9zo9x53x69VEspZY6s1FKLysZ90lEwHgx6VZ9
JPmrLUB9Mc7dFpNf/H9xWQyQYdE/1e3z0aU4Bf95ocP3v98C0aFmv7T4fmZI4k/W
mwrqGu+ScUZjSOsGrsmXj0kzugvrT3YT0BYEfKroOOzzVRXU9ahF2ledlV5RNvck
a8k2PxXUfvRGcKaHTdM6NWG5VIF4Uva/M6jgWMQnPCp28YFz8dIM3P0Ns6pwK3o8
XCakrswjqgR8lj5Eb55lmg+KwH0gc28dac6bb4DHSVmgUTFQ57P8i3YN56G/kAYr
BTozCHBnXRvFKGXFiqx+4EqMoeLCXRECrcuQigljrhDgS8zV53NET5vkvy3BUOqi
LO4jh79yjQdmgheu2xdv2ycMHKljCdNL3PIm9YJLvYF0j8yYTYEY1YdJZqMKgdve
rOXvFo8CGml4PGRL1VTD4sC4q2+Rm7VAlM4PGZhPmu6xqfbq6e05IESnSIfCZ/ZW
VguG6KzqH6RIf0H4A/gwmndn7ErfTDIkhHPE33uY/agYMr3ubTnN/hp4+f2YZd0L
jGaAKLzjRcinhoJahV+QPLL1DmRg9sKwVUwAhYcdnVC66IaPBQ6cD6fhGjFnSJVZ
89eUxuq1heAjqtFKKhdSZ1LI1owi9tsLR40U+d2x/D0XKcbFFVNY7pJ/C/Gp726b
blZKViA+phgiri/0jpUwFoidmicsXjDCRk8mlQdqrI2emD84+thacr1UdVHjSyxP
XhPWyga8pKztzURq5bZnpqvx2kIDYr6wpn9uAn/dJlQDevDFNDV4HYhr7mGaO4Jn
xsqlSDwm9PleOT8hM6wUR9TL4kv8ohQYGV9EWs8EIxMobyL7YJtibcnD1Ke/hZpl
zfyGyDRN1Klt8ofDChCaVri4t5Ij452xc4ScdltKGPLXt0fauKV3gVXRZx2RkWa6
sMSIyhWyxk4XPreAtY1qNC5KPrno2bVZUA50RAK8vuSZxueKsE5CMVPSrG2g1ZY2
2nf4icr43VE7gCO/ZpSwZpGNXXoWcHyqmysjifYWDOc+URE/aHneEZLSKmogZF8T
eEUZJMIN+t+vM4Qc+g2nSHRWuB++RfzPexfFQQTDeTIuBdRwCtKYT1+J/VzCup9c
Tne2gE0u3sGkEvQA8URYiobE97F5L/AERpq6b0wpLiCu0Ne8UPm88h7R+r1JPcdw
zu6ZSbKtC1LysHdm97ZBOiGuSadNaT+q1c8xDAZH43wjeRPtB0NM+PfHcit8w6JS
LPpWT2MkS3bxB4IE5AeM+4/WZ6C+wMzuatvOUWXZ7AcVoe9NbpmriO4iHHS77jJX
+0ilzD6T2LTatLTKoIZ70+VDq14hnGnZH0t3jVUFuPJlDp7yU0cMwydIi6CRY5PC
uD48lurD/eNh/KOej1Fpycs1gEgNyRxzUFDKx/p8v/BZPzV3ubNN4caUdwrjnu8d
5k5pNbTxAYg25bCQ1kIZjZ0uDzrbd6tS34Sj7K9uEGqaN5RyBGt4xZnEP11D0hE/
ZEX9P8YEIiy7AyYK4SxeftFcaARNq9NxZePtAsWuM8qsE4qYOrPPF5cSy89RJf9C
O/j49QrloIS9j2YTQ0BeYYkD+s5vMj7aqFJ3iIMYFc1CjXOUo5xw+XWUq63Y3Lym
QM4CFcFxzYTcZX34hgl2SSXIm+VHFAW+RIS6qArGDVlR3TSivQPEdbU3hpD8tw3y
WHPIk8ks9qibwrOqAOefofJEszsIO4pZKNKLuMPKChb059avCJiU0J1XngedBqw/
N/HAClAHv7A3CBBdd9O9vGGWVmeiS0RxYZSr0arQjOOnqueclLnEGcX1f/oGAbz0
NehL9FqvT8XvGZNMZswliNh4FebkfGlcTWdX/isKarjbImdB3Fu+/FqcoHDeg7cs
SEccnPydK/jkTEo4wVsQBSard8EDqaxOjHYO1mVwEZty4PUyo0zmDGwqX1V7YCQ8
gCiJLP1S/JoVMbmTsUaKbm0KLNtTj6oN3/xDuOxBh3noogdJToJNGS71mXCBqekV
zkcNhP0VHUNNXruP74WkO2TlemmcbuUK4xeJwCKLheMrFw8OU1jAtLVXZ/JQP/VV
+Ij7XddeDbRgpJfr9J1WBeHTUgQ16U9w5nnwBXeDVlWdoaX71iVfnN82j58/D3Mb
EkiN05fFASNYrqvjQC8mw/qARkwkmjJDDQHQrDa1YbgBIRdCo4BcyIpRpR7KIzpj
AC+XceI5lA1ouLTGbShRDRgSDNN9cfrTQMIM4v0TPTAphX0VEnuJU6BSOsKbWn3c
PER9c7sNhKmAxzmLhK955y43gT3v77RC3bwo+pW+/febztvAjb7YXSbpWG5F0ouK
99im2hOm3uZh08BX9eYzNx7jiEb8IWf4zN9uchGRV671Csr3yXKpgYYY6QbQXayY
2hoz1hE9UWnqcP3RLOqIlLraZSqt2nWH37dpCqS690G90c/NiIzcXeOgus9q3vDD
IlL2Pk4Lnt18yq/rmryJD2ySe5qCkLoi2H30GnrZZPC8K+gGe7+SeYZZ2hHgd3rz
5FWX9YwUOFirQeWJoXiYgtG3CuvxbnvLjd/aaK5vPPegCsNgZVL5uC0I3NXVHR1w
rd/CtCOx7e04L3XwgYAp2QEy7FsxxA3Pep98/FSpuyyWu7phv6Y+s35i7Z5izY36
MFQkyhv/qIeSHFGM6bWhPzjhfE46HbfPCDGgip9wZ8LihLXWe65xi4vGpcNM66mj
+rErW4LnYQtssKUeM2YMwUrC8a1D0oQLbJpxKnpbfCLAgUHtsLRpHykzPFZXzRiL
+EXXRO6q/9xgyCwEIDthYuKLavT4G+ewxUtNpk2LrpqVuEkVwL+4mPYJG+/C2hNC
+PPP7cmtmYfmTNvc643+D73+6Bs50UTmEbuIu1iZUrwAsbTD6RKK6Z/C3Oob2MN5
lx+uIA8mAl2bUIdaJhCo70uhWpmJTNYrAfluccCuzO4rRTLm9Twe+8MfrtPfWO0s
PkVf7rqifWB2tjyAXUoAUEbNzrGTGvq/CTWjtoYfkGmQYXVZGKI9yyDO/LpiGFJB
/qtG97DK10HRD70FvwvRROGGSedXm/ZsLLQEMW2aIxB4Rc7RoveYjP6oauGbvypn
1lX6e/g/eZSyC78+ZVcMQQYmcF/8HhZK2vrm3m7VLgJsTaZnjFH/JaaBryJKCJU8
kXzd8IzLm2t5tePEgNMGGMqNye2YJ1RLeO/OhTUWrO6PAZFowrNpa8bFGpGCRHTH
oogmrmRB8px4MlRjOIvahI36eTmXenIUsfFJqE4CkOzgZPZ4ZxPX3BrzcA0g7MXS
z8zn5aQ4T5fFbylARdkjELBOn0hH10RMlz0uBVgaxxpKe130Gn7A6nn0fttnqTH/
MoNzykRzj7tFYyV82vXRJ05I4CoLTXXacoKNjq9D15j5cgoFZm4i+N1a91rEkv6A
LtwLkMjXooLVEbI+XFmzKw08SsK4e/mfoegaNH1iWRZcPju+ocC7zQ95oZ4HvuF5
qQo2dY4fvSQZ7pJFj6nAPD2D8gaBRyjnfYwJjs5b1fqK6CuRZT0Bjxanv08CxSBY
l6wQnmT/BpknP69K7FyOOJW/QeivsKw8pBf6UO8Kc9R9ihJiBFlZOHcbpkd2IbQp
abII24HWJ6tOa6/poRDl3QlkHNep26fE5VccF57llYVy7/NSckuTJV6sK8PbRdbB
gGk3QWu3coxTUHbVqdK0iVW7w9yXAmddFOsaKE6JbAXS62dvGS2t+DZSOfGeEgPj
kxosoIK9QHElY57yjqs3/dAkreRsvXwGLToSEqtUHJjduWWXiEYVr0BYYZlDOU4N
FbjOUhsfr2FzahzsraxPdsWI1pJ2cnfXU+AroSpC58kD/J+6nkY1OWP8yR9wQkVh
bL8EjcSGXGQroauUi5ZKVzGVbLAxGabScuPWSflkzhwhv8d4qxTGDcV0g/9lPesu
3yJccMIO9OfE/h4te5M/YfxX0nxXJEEaUJ50UHoY5RCFYpexByw+eiDz82uuyd1+
B+JoqpvJSy0oij7VS6PUOtdBULjOAFexfmvwK8Zt4oOc8njsREWlPg+7DAfoLjYW
hCQPp6bKNryFF31tpzkdkMI4KNZr5YBRKZ0nB0QJFfcFKz7frcDiVsP45+Mq4Y6x
lx9kTY2yxqABjMNzhR42h0eCb7TCjtIaFG7S8G10jEuKcnXQQvwrctQ542RfeOfT
DjpyugTLwIFd9AxZPq+3xNUbsWGVOHbQ5NEZVRBPpWXeiotwXwur4+Nhr6EaH8zd
okA79vHdppvG5zDJgB6UvF6HwDyuvHB+Id2KQLPZYFR/4p3I58CyQT4/KL/7wbrt
/sCuqTiCR9+9YSzG/vQzddxa5Xrgd5Wqs/2RaFF+pF55NIabzt6VCJeo082KEzxj
4WL/DYIXqPI1UhoNDwQJ7qUI5jXLgyCBAh/21FFaQu94R74ehsKwmy9OVwloNO9M
oY6+GxbCDEi5RGEkSD6dKiIKl6Lz2F6p6RuEiHw/xPef9a/wJBL7aZfmjGarAf/Y
EgFsOztapeKwj0R15vBPP/ItOn8OLpWkRWu8lYDVyhrnHcqg5Hnb/8CAJ0YgX3Hp
/M1gblEeRTA2/dfvui+MD5IMO+Fy18vL75fKR/X1uUniR27sBqzmT+p0/gyH9iBd
zKPAXIpTdQplFi/qODSgWLEFDPRZ+eaibEe1y+TEY8lbHHKYTUsxFlk8kR9JZUyG
dBPARL7yhc0FFxGp22itKiryQ4YNkkt68HXWbxrTE8YABADC/nJFD4D5ztNSmnQj
XjnfPdBUDqThukUccW30rpQ9+gRVYrI3tcJamwCklNwydwMO8PLFQPuNG9vKEsXo
lXiCqNb4EQJP347XGjhaqv6YHWm0GJa79P7WWsjs7qSNk6GNr5Vh1NjBS0S/3Ecn
gJssZ8hIA1i61xHNJxY4Mn35mvHpLuiV1tsNvgOTfDxmdN+JUe25NRdeLNZy44rh
7jeQL/EkUEsNW0Fa0Zg1R8JItYy2ttDTbbjb2oV8ZZyUQLFu1MXlCJjXaW7bdvi+
r+6a3ENQ47QdiiYq7nWQtDzKs21zZ4YDkhAf0hAITv3LRTIN4xj03zgmjRAlhJ+8
5zt9E9q8eAmcLHU9mYM3ktUfRfHYPGApGyPttDD2VOC18LDpf2KLkOoxjfRH/otI
sVT0GBsP1gxB3OKvLw+b6hdNxcHyDA06KSGi7cKZO1Y7toqYj4clkG+VFN48vOXu
rTxzhgtiCngNp+NICwHk02R0mZ/bdw80HH5/H85beuKxRPjg+21U8SO7tXOZ/JFh
neTdsxmxnFQmhakJceKtGBIoG6YGkXSlPfsQLh6OxJbD0pax+Zn4Z6M0IVEL7tnf
JQUcxBh5LkQj2KZW/5dJZkAi+sETMjKTb6CnOG9s5OMHg4yysaLTURmFO2epZK41
qz61MU4BI8PwfmaZN8KPrHWqwA5Jvo2OxKt71IRF1SsmqdBqiuMlQLNc4zKB3Axh
cbP0eOd3m50SuElC/WA7yfVCNQR41tCYKK0xHRNw49GKML+jZXKVuzai+QQySoNN
+6lWFAQKauN5DO+CqMrUL/lqKjl5lKK1ZPujZq7rHTtuqFrAq0txIAGQu6jYGp6f
kU0SgFrWRci9lloaJEbHbqnsmOtZpYvsLyd/0CBl27yDfQpbSK79m7j1WAfXoGef
YXPlt3Sc1DmXyz9vsbmmZ9IUsI3KnVsThQV7Y76TpXkuRgqesifBa563/989afi2
YYKIV7NDpGMvBO9rfDwGf980XSWlUh1sJPa/wkdaP2q5CJMyngsUQAM/H4h1y0kg
ZofvTrMb/ycaqOg8Uhqz5daSHUImFOPQLGfVKwzFBRPTNNXiHM9SXY3UN+Z+jR3X
TZUn2ClVbx9xrvAdqYgk43nDn+LP+2fTHnzABN+vgu8U7/o9ww7DydxUEr61HW9U
gwYWRWlmE8ci5G2BNIivOCVq0AU4WrR/ZWzFKxeF0+qLPBkTxVwH+ll+v/VrbBat
d+lAXZv/9OZOuZ9DWtZEkEyh7ZVqiI+ioCSz2zu07d/ZaArJnDgfZkDuN4ywhKhe
FFf/yAkKNUjjumnTrBPoSjGbdBjatFQOZNQgXJ5bEW+Lgifx198q4iZcDDAGngjb
JLDrjFtWWk5N9EygU/c7I4ofCHwISc5NRb/YWCbCOGOgxuWpLIIKvm7uOWmta1J8
fWmUHhV9g5XJdCbAf0S7pX2UQSbtQ1rqijR1CsN3NIr9mxWs8C4tes/HoetT2wBf
Y7aA5rmMkQPx3+AdwOzgTk6RSKiENbXCokjcW3ytkteBFZhsV2XWBRm99091pe6X
YWG4yOffzmb1DhSHWEesiAOIswMwe23QHh6uF0KY5od2qNm+1vJO4mWy9sMDuSP4
cgi7tfJEmNcOJbl0eBLHxlMceFUMHOtEcbU2tDN50wertwfQYBbtNx7g+9q/pmrX
eyJXcyJkqgwAIfoYencOmPWDR7MyVmyfSRFjxmqlrjF6qU/swAdu32ZjIvFTnjNC
hJu/AfV/N/90cMcOP4pf/kJJXTxd7R2qK0FHxxJJcmhkhucbit8iCoL6PaJQP2P2
/6ADhqmNKXZceHH7uZUf4cZIyc3UbVGP+A3CHsFRoIYeabx83N0oQCKer/qyijyA
prhxH41V2ilpzyy7MZZlzrdUvf1NTxxHEfbXTY/H57nHyk6QBlv/1b7BOc1irNd9
eD994XAmLFopSljAYgLijbmhHUK5FI32uppOnhGiNEqh26bUN+NMX5cYdNEAnE/z
AthMUA/XPULmvZC+Z6e62MULrPHR+7UVldM7PDQ2JQ2jMiY9EvIv1j+z8SW6SxPO
7wJwD/P0nkpx/1LC8TIzIBlbjhSyNpDnsruImNc80//ymhXmpUKfLIk/pFEyroCH
KZTjvw1BkAyVKVFxrKvn5NipuJs7ZIaa3uo8RiD6lonic8z5Ya9mg+F0j9AUsOz2
Ry/WcKTY4I9n0VnIBNkdn34jFN8Guq/BwbqpyQLcpAwidFDZ3+6Ln7BgPsZxOlsB
nB22xooU/27FutwyqIgwcYL927To4FBkBBTimZDoz9i5ftTuhSP3Cqz9PQIwJnL2
dn7JOw1xnba23jB+EOMPITKoKTS7Hyym0FzK3Obg6F2L2BsaVIAn494aFH+DHiXX
fjorAJeMH32MjLXkNzKWCT4n0pMOxwyfLmmDK8R6sFodz5toJcw1iRE/C2LmjPhb
1hZ2KLVF+VJnmQB9QgHHZjfyBen7auOJ2uXnETdBUy5SSq3gvWem1bFjlv0LmRza
oq4r3sD/icXXqLPgO8fcmVAKHjjuXHn2yi0TfEGCCCRyZNMJIPm2HDm7zEJ7XJI4
dggNG5fO1Xl/J8BgCedThqotBJxLdG/IRmNLG20Th0MJ4vdsSLHdHr/8vXKHI0Oh
cnW5mDQjh++rszjFMjm5BnHDsVS/EFM9Cw/bvFgiLoqRkEV3ywswm7Az/PQSQSad
nnIxcT74rLouNEMYc1FB9RTrJbF65CRnovOjkuDthRiVae1lOeDHo60JdiA7mrI8
hhPXGZINAQlpm2KaE0RQCXHItfKqbpQea3hZ38TMpg5BHQdnlm15nJvGmZLipkaK
NyIc1/CTPQyX5Nd9PHOnKDDQZQe1lWn3NpnJVbypPcue48TsUlD4uy8lZ98VdXjx
NtSCNqb8jMDCV66Ss7+lJnpL+xXG5qH/+xW47KYwzkpya1dIku15uPbKdlY/tf8j
cQBKIKJNjS9SQ5mmDygPbjKYOC4Nhh0bjBYbUH6/ggmUbjM1gEXI/O7b6yOBpXd5
normIoTxGLl6fTxRYAfXgAEsthSWJSA+yH20dA2blK8Ku5GqsWSGSRouO+jjmxIo
mrJbDnb0w6sR1PEgp+zpHT1US8d4WMijrPs6JU907+4oNLB5p0Tsi5pN4sMy99J3
pXbqMFAy+KPpfFFAvmDYgwPnzzH3q8J1PYRawThk8SXOAIo5yJWz6CN6imD6vVuy
/mhg966vYDA5pS/tnTfqYvnL5Iop09zi362eb0Zsd5jDTY1Pjcx3wkYlXIRAPPn1
fJYURepXhXMcLvX563oecFuvlV7Jqdc8tvVV2Cz2yKk6UD7OWb9u9cXh6UF1shgG
kjuN3Ph+ms2baqBtNI/S5kGcjfWqt0bxshOc+/F1DoJ0nzGNYw7oeLjpvilHrtdd
EIk4ZOt0LG90pLibIwuD5IpLCG8Km3ETpbUsD4fpRldplFKHad9X4c/2SZErtSfA
zp0kVWgglzqVnHbQmc1jOntEEec5tdgZSBWEXAiymNtoqX19wUlZ55Pk4S64jpCu
TeXftXZX3LJ8URjlX1L9qi6ihflE5vJieyOYMmoYXvlfBH8keBydcJvufPloHhvT
PwJEvW3sYbxqHKq8SrxLmiSo4z4cDVRrOptYA1LwC3jiaYglgAU2C60JQ/4Al16g
LEOntQ5yaVKvIN4ncZkI1tIP1WhNecCAYmslsiYodRWBwXkcAHMbdKyK4236jDwk
rqObmv/2Fla4sXE+I++OOrgU9o8eVU1l70XnV2qKnN9tCb9MZ4GK2o3yPolDRLmE
v/7KEzfh7LsBxsfSrP+v5p0DYpjKRdf0Y9T+WsJTpa5F4/cNDF4ksJMMipKwZMPk
2ouFSzqxeOlmlozurKp0tTrjq2UrBB5/yic3orYxXabQGculgKRoSf2J3PWCveMq
ZSNAKP0x6kJdFsTEJB7rUiaCKo9Cv+T8oJsrzTCSDvAeD6XZnPLkCs0+TLVGwMJP
nuKSEVi8j3LeJqCShgEplQgZwry+bOpeAc1tKxqMRl9qWInRMCUVGJ59AcFn/BWR
QRNG1yCepKSGdvFXOp5W6gyUxRTdcH9MVeAF3s0+5NUBhHEd1OZrdX13cBOrFjc5
UtO0+ynER5jHLpsNX3UYmTMpYid0/u9hDw/R54F3tpGEyQdw8eKdHPlxGicGSRYv
lg9NdQAZq3DV4G1wImhJH1lBr6owUobrljJ6Ya4e3K2J/qHoNOjZrjtpy1DIHaHb
Vl4T5Lt32E7HKK3P7tsvF0oDJWGvgT6epG4Szq3h/hbC8juOmnbGQO348o+KZIgq
JxAnEwA2+wktVZ0UtjExQQhDHLz6O79W2gpCSkR76IUuku6xpld0UNWUoRqqJtxH
fcSHbhIf6gy4nJw3SiDRsp6fj7IF9PYvhrTXO5HRo1WB8L2Ynq3+KpY2Wi/fsc5u
2nLwWXoaPMEtQpLxjFOTXoCAm1FMOrWarUmf78YLJTRA0vIS1KwKeizlXoo9YxlO
lqlYJNAjWWMfzR02tVlJJ0ZwWCGINtFFOEMFW3F7xqmvZ8PE7zgVRstAOP43R8L8
8MWIqjW1wQys/SWtXLvKj+P5HSu2SBB6curjz74YWMAaf4lGaeRba8XHSLJmWrAd
7X0zh5raES5TpBriRaTvgt9wCKsbspUtgACjF2ejpcefrU09DewuomdI8q7qXGPW
OvfYRzw7RLEGJzyWPZIo5WgLxmecsF3P26yTVVslDe/kfgKFRvUUIDM7yNhzwkGq
65cSK8BghVGCIHpNYzXUg/f6TqoHQTnXoZWUaOc/e95OrH4E0zd5aXnmmiS0a5zl
JYzFV2y36zv0w9aS+GcbTTkIdHZ6jpvylb3MlmL/xJGlnano9HSnBQXjsRr6Q4e8
A9NinemNdrkqBSQ4jjiSAR9t5YL6RjrglQk9/6b4Ly4RrkY/Jn95XZf2w5rMqGBR
iPZMqwL/fCmBUl0IJ+Dk47uujXeGO0xuk8RfO74eawOn7POOAwC2OI8EQJDvE5Tt
5nNm6jtJD7gP/OegBQmyPYTsgb8cZCmWbKHdnita90G9z2PxZj9BYqs/TT6Onw78
8pHSP/B9E+LluQ1rToxhNppDpez6AHRe0S78hNPS6hkfS9Bc6nIyeKnfQxrolbgS
yaa+6gwQMYIFhcuy29PzQalV8icLFJyQtkhtgKI9HVfUwsv6scp1JnjCpGFEmuCB
2FnsOmf4Rf5TxiEvtZL93D/ZKhWfr8IJHL/aua/y6V1DAIDpavSDvgKd3pXYIkdU
11v2ax0IyepU+Xb4j5SNdCUKkyTwSop3Gy/TW11eY9c84Lmwo1atcdLudT28SRnb
hfEDIJhDKVTYobefh10V7C/P5jxdHA3MOxBM0mlVF+yMhZE54p7a+4f1t/2oogb6
AkYZi+9rujIeZhRt7LlD7pTApz2PEX1JTa6B58DnvxNlJ264bZYIQB++cS4FPwdE
KNKjTEd8Ho1wTxNT+vMdP4YTvfXSF4YIkWa+ZUDumUIF0XIwm3a+t6NHBMDwgiwu
wyP8eq+UR4zIb6BRMATHjWau7cZlZGDhnB590eF/Ifva83XnsLqRMFKj3OlyFhZD
TN28BOiHp9yiBg196PQJZOzkjQ0IVLpIc04Fzo5ZtpAbyzazoUnDyXkcjMSHXMIq
i+A+lPjuh4GLF1GSPZzRtrtgLlX97rfXktJxSzU5/S3rKIrV3i8KJ3QKbhmPLIwD
iiHxxyl2eS12GodUSFqlJU27xtgOei8wFhPS0fPr5/x0MA+s+OFAllhyCuhOkVko
5OrVl52DwWLc/h3TO4suyy/67BPCTfUCtVetwVsc+yxyB5a4AEURzdRUWpu38/us
wWb9P7HM0gu1Z1Eh9CAmDLK+gTRCeorhl6KKUcaO07hohHJn8WbT927H4Q1KswDJ
yXKhwbgcAPfbOrW0K0CRNwbfbsc9VwoJnPANw8vPCAJz0rsLQElZ0cDJgiwIyoWi
geRsW2GQ2sdDNIm/qH2Tqt+dU+Juiae14MW+CXKj6oBVoXwHt+ajN2hJGrPKH6TR
2ZQB4Lg702VJcUu56xgknoYg5A3d81rnKy9FUKv3ST6C5PKviF1RGxNn73MgYbta
NrqXvzdki4v80UzaArTm5A11wjWQofDDbU9TNGEbpWH39liJ4HJlJjOujyjxGHBk
XkghE5lBom0JaW6DwCz0hDfhHs4hFPQXJ9a0TxdgdlWI/EoNyemmwbMagSj/WyJu
uVyBiPTLY8fvVGsED787fkc1I4baXCCaMIhvIcSRsjH01K6577Sdz5lksRBFlyPJ
2aOGxj7KwDuVfWqL94iUS0+9GguU8RWTuCVhxk3/mYYHqe+MoDI8KKpZ10Up8PQD
LyIVHWTHnCWgYlx15U5HN0Y3bCD01LVY0g8N6Rd/CWagDuTgcJVzf52zxKoQXrJR
4E8/t6a5/BoW5mhyI2ZNwTEiZBaGMnli7ldI/T07hEpahPHSQHtBUQr0nVd4ryyH
4KsFUV/rKPxzlqxl5rmetI/7pqYgPRzgWCyeaVlsuoAwVR1sa5k+mtdKaNV2UOPg
NGcnKK4mgBDsPo9YSMX2PvuwntP1pchKWuK0SMx5I4//rg+Qdd2i1tZ7+g2g18HJ
6dM/GltZP67p3JLVAlwndpY34vJlG7CZO+Vmj6BpqFGwUtEcf2ynUkHwxjTcD2CH
FBU8aG0WkHkmTHpETIPwYKJihI8wQOZUTMEZdfONTRE4LZJyNUEXUjKtQDrp1GqF
rCugo11zfldXsEsEZa607Edz3nQc5lmsePm2DuAlLR9T8bsYKDCSyuwgWrlJAYeR
c8t5cYiEQK0IYHGjK0bDrxQ5d07rqha7/63vpDGzExnw9cx4raO64jhNnzqSJXo5
nEu766c6Ir5Vy8bQjKf0l8+2OqixsElXIepgpOyxnFDZn7FWe8xxhUB16z2c0sPT
WPkBznPbQMTh1LM2Xk+ZqIWXe5ON1ngjShgdIQVZjBHfSg1nl3PcYPxxhbFlLcYA
FIjd1PtAuPouBzICArQm7oM3aQBga/5+TXaZL2etmPzSlox4WoLrRb+seKvHgjp0
CVRREwBlM6NRmr+mTFedMQV2nX2pctVKCPlebj/x69RNWBoFdJPW1nxZz3g9P4M7
N0iycM71irPKuC4XnsIMZIi1xrXlGkWkalQDV5IT96P735I95f8bXD2ddjUJuZpm
xWWEDG6VfiG0t2Hmr3iomgo63CsuobiDh0945mwB6vMlD2AuPZgRWxvFnjPadE+k
pFSF1kVKX0E8pcxZpJElhrIz1Bpmay8IH/+V6HRYarGD1F29UunYL/f0fOvHz+zn
t4K5HVITrElI0Aosy5iAkeoGiSu8ioXzFQTs5lI8Sq8zwVhfKm/7RLYcKGZE2fG7
DetSCPl5InupTMRxNSWeULl2rSBKlNwEW3rqMEGhB652Zl23Et1XgnTBbfuT6jwg
0JZcnPkfTyWC/WiNnz+p8l16KKUV+Y1CQX8KdV8hUhVcUIsJS1DVrwvT+fOmTHTs
cYB8egw0ebPz6SqMAZ+qkUi/lzGWj8fBPi1fwcb9keSy4eeCQAsM1/TNdLFjtBxY
soL9myLAIQ40JK0wrBgOvnRemEtq9yrrf5EsB71fkN/lcWjCHpNNl8oid06tgsZX
9gNoIpGBrsTNuo4WUc+iuj0yH4eGJaCKADJQ1DNCxQZdK8sCvhg4i+8OHNs2EB25
TdvMcdxAPhtulaoyBFr13+Mmij6TfvNZCGbxOQ+mstvyqj90wj1Fk1lHyOx1lCvv
lURktQq1M4nDhXnvc+/wLMZloe3xKcjJkULBe2H3laPG1sW+IPVNm0Hh4FTmvAJ4
BXX7RkI5Jsx7tvEEIyRwbKsc8zRPK8pzh3ITWyO0JOn3bQf3nFJuna7aIBPN6tzH
Tx8sprp8f6ya8urOT5ukqMapgx/tCWAm9F+VuWFV8/XAiuBYtKumvdE4JQHUXpUL
URMSvQCfPTeqfvmRLOmVfx3p9N/DO9RCeXMzipWkr/mG50ulask/mkoK3J/2sVlN
uU9cgkuHPGE6Z+TLVnSljNfyJ/+S7DuYMTGFw5JdeAcGhTtFo7VNm0c21dwEuCTm
KdRexeBBIzUboWWjBbPTKfI9NNo2UdTMJ+yl8Qj1mRvdzkWVfidLe6YuUxvd67bK
9H4I+wXP0s3ZXoA213Cs+yVfJg9BPRQEpuv8/qX7kRD6k9uP/HuLGyIi+j21Yybj
oVuseCNAWVuFr8NkV5f00/oytwNiFuRTYb0DGtSq35rlj3QhgLEgvJZZTu4sVcNz
EMw4yR05IUiSJyRaNIxB9WudEuSH6kr3Bym0hJl5fmTin0qasiGqetyUTm7tVK3S
XTQqodZRRGFen3NZfSBNSHG6izfGqKf1GDbR6zjpvvlqvj7o2da/bhMO/5LpIUUN
uj3L1xO1n/r19maF2bt+uWFMVefh9RxjVUnY3KxtJKwJCMOLBAQkNTSx8AuQeAty
Ov3INbRS2OZdgAIxO129WxkWavfsy99iPza+61CeN9SqxzsNatJUz1Q63aenYX/q
ZNvsQ/+E+4rw0kjXUOTBT1M0jP+rswWuKvjc6N+p7F2lOoqH461bOzFlesQAfLn3
QG39T0OkHi48dtaxtN581CZo7wMEHiOxPgp8llIS/RQLZBse7Rdl6KiGaLJ+kRLt
mn8HwtDNM5PQ86T8Ybc7lvbc3s8d2IlG/scfiqM+g5Vse3SmUqh20lVlJBGQ94JV
z1QHljbJ22gIhEBB24yUfJFf+SIE17FtqAvLnVXPUgH85q1LOLdBhX0HHOomTZB0
Q+rR0f9Gfaw1Mu9+IHQxYpkHVI3040asqRVaTmixuJgBJzcWqI4sUjiFJislRiec
q3kOwvLqfN91iGeQBmJRNphY7EsihThieXDziw0qonv3maTkc69S/5wpqYmczKm1
5ty9a8m1mtwC7U+GHD1xiqB64pcqejSKG1NbAcQYZfTIpgB7YyJNZRc3AV11a7cS
79TWkQWYRpRDcyIpg9CO6dtecK0hRohwvVlB8w5REIFhZ8/ACo8cyawqFdesczh/
2i6dHNr/uVDOst2VRCgfe5WFp++6OicofNp0mfUD/Dnxw8Pmj9kXXTMVtVsAIXyI
MQ/NUMmFGkH8SHnSesuu75jB8I9RZxrYStGyNeeDha50Ml8MV6+O/2dET3W52PTY
0uC4nHanlOJTVNemf7WQQAWWaA4v8kUdmi4yg7F47FkG6khP1RT8k0HLEap/OxoQ
EILXOfxTdlgcXoRGaEBpzp9O+ipPlSue+vq9m+WhzR8iYHdMxLr1k/pxWXSQhcB7
cIwomrWB6AMCns6Oyz1nU3l95kcCcMZOu9Apwp4UiR1zdI7HRFv93/mEfo2FK64Z
m7UDxEcS/20LZ6bsjA4SWQz9EJ3vjkSj11LwGXheo6v4AfwmJf5bw4DR/LmLi+7D
8x8N2SUZBEWu3IQj6E3236Zp3gAzKJ0s5Lm8Yamm22+dHI3S0r0LgxmayryH6dBv
R56+H1NlwfQ8vae2NBFmWkHuMkACw3a1smVTqseftkeWa/j2fcnn8ejBiHml1sCS
L2dBvgJOjmtuco5S+vI9PakwJl5zSO++a3OmiYv4Lg4XGVGQ86G1uP0086Xw8Drj
hCV0h3gaWEHIG+yaKsv9kS0yhBElyjuFASoS+ybxURCHg3xPLc0KEF+0jk33v2Qn
pOtHsG4N4z8JPA57fNKBTlf+cWGYGg3Dl9MlCpz//WRrcQbcPaJaVld8UuiZ4sv6
Hw9UgNNYDFUhWs/B+yKJQWNMeSo3g9sgkXfTUHNNfBTY/MyjTUFYp5prsDhZGIpt
TnmGkadUcn8Cyyvvi99nrN2geqMCGt2X+jbi9TYissNztnwtcXdmYFuYlLFJHFZ5
CMFFlrZ2iJYHew7qbB4x9vLanVbSFZ/sXVrZY/ODkXGErCFPtt9x2DPTVupOEFE/
25+I1Zoc0u2bv8iulZBL+vx+fireV30SAC0OusUGZkUQifMIexZwM7+Q6TWMYaKa
S+S9WstgJ4XL9nAfo4vqYbEzwbGO7wrbssc3REcjEcdw+KR54rzy7x77drfdN9qZ
6lW0tGpVLmHGsrcqvHKezixDSm479OifsIU/m1G86CzAWbxSPLXUOqJ+vqwHNkKL
YM7zH8nXLoj5MLb5dkkszyfpqukvS9sCptuMzhOONsE0ezP6U5Lsb4lgwI1n2F9t
tWJ7J0ihcVdETuh47zgvOUMLx03NfSNfJUMct2F+Rc0TLbra+zDcWzOnr6oHvLUF
Uqkd2wuv9TctWnPpPI+nCqtxrs4TQ0ApOiEJiICTsu2O1mBbbvYCCVKmyFjUcZZa
Dj+yU4IByYq48lHjEA1h/mYVojb0r4+LiNZgwRMuqi30Jkz1KeZxsyuQSVtNi4pZ
Zp7zVlv0errSXQtOkrhHtMiPN1F5NMpjI5npbRgoC+4dE6sMMMT0lCKnY8Hz8+dT
fYJGtR3y5h97nlMLS8ETDz2i7BC6C2qOlBWVsMIMUwDytWvyY7DyvhM8Gy8nDdq9
a52EKKlaPOo4ZEjOxpYvxPeyOCRXVOU8SvXrNPy4RZWbwHTUSvqmGQO4wfdUsZeE
HBpf4Or6rsHAekbONWkeHIZr0Z0ATkSzAvWXlKjNshujNZEYXw7HY/Ebc2GP8pSV
2tr5DkIMsahjLJURdcYgVCuJjvallhJpmwb0AYyozgfXpgc8h6wUeagHtouK+GTR
2FC66p30+YFxa3EpnOAXrYPLM//fyI2J9yv5Lzs97Wqnf1dQMAUoi/nXzOjp01f9
TddGYhfj/f8VXwyVK6jPduUSt3pJGxosZJljTb8OBg8rGhAlnLCqNYxioVevRFB1
Ofda2Ue4JFyRexobMHWmjh4JDN3r1a0IXCySy7UeqG1vtaX6Avb/PJS0yd6WBZI5
6gzsFBrKja0UHHPCKaaxdRkkT/gUuU6vDb/5DllLAWfmbtHnozUoborGGzqD5r+7
ei1K8gfAIIvpfw0QT4X58JDvSQOHb0dBW27S4lq+kMFvInRvtVCKw9tYT8mOFvsx
mj9hrSeaPG8H32xWzZMn6haBa7/OpyZRnvPVoYvtZbXg7kNNrQlVXCVV9PxQuP4b
fjXs6FdPh5EqEeBeWRtuFesmmMYcrqyJUDqRzYFf0VgPbIJACGDWLsEjlqaBRabI
qOIPC6IlRZbhbaVympFiRIBWAWo9W9UEGu117kqWRfCWTj9vHXD0zh2bua4bFzeh
Tmft+0ZsVe1yidmbDriMxCfXQSnBU2lLvFiL+A2ECDiWA2CXxqYvaTNy77r0vZ0h
yryGbrSkNA85TsqFb2WzNgZdp4vqG+/hDEp0PESJjl67Vj+yQC5vwOAqXyyR8lZg
eFnNJEFS6EJ2aqdsyXTsiau/o/rU0IUyKy581KMyH72Jv/azGgo8mbOkiXKnnADj
tayzynUEhJtI5V2krSWqj+1iBGHLVYCzW00/6SJ+XG08wH1s6uSW5LlH6lk/BTh/
95NCdnpEGRQpsGLaEzrc5WBwnBEo7rh9aa+8G3ibVupS67IqrgOIsydbGScOcBuB
U67SwQqTBG1/9ENOTBAwtN38VnlRQ84Emg0VCVGQ+wM8uio3rp8ONLljx1VDwbqA
jvEKQ5dPTbzYMa97pm8CtbcKMj81jKBC2Yv2uTGL+pXmb9az1y1GlBw8JdhT1nTP
es2SHzYd3x2Kud7OPNRRdQyTZx78/AJ8CJlboRA7MXJf9LFXBRd8dxgB0DdWOL3V
jDtkmpGAOJvi5cP/iWHdiF2A4D3qztT4JX4FReJruu953yW1rndBL9F4Q7WP9sQ2
z9ORRzzQaNrj+QRubB6X3eyIKIbSM4ilhH6fPj+z592MkRaIInkf4Co3Mum3RpzT
oqBpE9ZDBOGOFgAE/JIYTZ4wLkd5wneqkSmYocqssy4ZdzXuNBUHvGgKqDI9QRig
PukAM7Tkvt/aojYZubalcrZfhePABGn9YOcS3esfIaa9fcUxTxOyLqkqTAg897Ur
hc71CMOuP+w9XK/XFQCFCD8tN75i7yoanVjKz4OtHYcpY9JSjmb1MW3ImZ2cSesK
Jnv+DawmreRbrcpY5xl4DhFfLcfqp8kSulCWpP3UJ9kI67Rb3+Mq6kF+GG6ntKai
wY9rIC1wBk7X6gYueOkEoZKH8PVyYWVswZQcfoU7Mrf9grMnaCiV/xHK3A63jwWC
ByGJ9xX3OEHzTyZmmsgX8luntHWyHXLpNDut6OOMkR6X7ACW0WuKOSWQclJtiaX5
wah2SS22r2RtpeNGm3aG0+HRvw7uz6ISM38Q2xWbS1+6m0LsrSIdWzhW7R/F+oDd
H04IIeESirbisupqrRylvH2cVCQufPilfpMkwc+Naa97KH6K5XqPZ9DkIZQGneh8
I56mlsJWshfRFs6ypmcpg0luetxohpWcGC92bv6z2OTxCpMNe/oZlxvtP6Oqf6Gf
pfc4UY7PyPjlCLcZmRceLfT+QKK9yEm9s4Uy6DZHLViUo3meZ1PuftdzhjMz6hy/
vaL7JMMA8xpDR4t6CTeXJUKkE5Aj5dm4Tid4WddE13gPEYSuhQmgKioogSUlvpNN
lEJAVrBoR2kKt5K1FAUusziX7MWbTt4pq+lNuGhIltWLKokmrT2xindKGqMxpPc/
UJ/KZyoMEow88aoGWq/99NqzxAGHf2sAeWuccsU+g8rZjB5ziMR+viscUqnuclmZ
BkVc4kIpA44MG4oAYYveInzb+V6wkecBAV2Mp0kROluo3IoERjV+Px66JDeCb3MR
4KZJ7SYkgUlhFxQVZNLs5NMYNQXjfroJWWFJhQRDHyehV2jaNu2o+rCF2FfjjA06
cDIgHakU1y41r7kgaiyeUhn9t1tUjb5O03HJzzGvAtmvRGSW4rEi0R76bX/lQe7v
F/Dt3W17IigR98/TG+mMbL6Ud0gF70Nain0FK7+ykWCxy7McLIaUqsSu0ppHErEn
DRPDZm79keEbcjNGDOPEer7hEtYUPjUMPy5XldAy+/PFl2gIzaN/gxkXh+kriyUh
OXOockTD1HTsxXc+l4D9Cj7jDuq+MlCc51KRsqKWPvRrttGtZGfwOzk8h6+Uhmze
EhHRgrs1iA6pf/ZTUzUMh+tdJaXEyO1Ovhh5auMoV4Ay4i8k5N/dyoOCM9LmKCDp
l7+G4u9fxjW8s9/uMJviUEchdGRod4Bn4EM3FAn9kIYDdxt5RP+sAYTAAFM4vFLA
Yv9pxojVQvLS/uqk/mEjyL7EE5vl1inheH7U/ZzE8KXutbO9P06iy186ZsH7yxuC
6sDSWnbBzy2WRMt0gSFcdsCEOe6hoNEge2DehpNQhyaBEVAPY1w8rfaDNYd6eiTP
ZWfgKsqA3BYldHzWFPGxyuSy42nSmRxaU3ZS0yj2/Flyls370ayCTCPyac9dJ6xm
oRm8X6741JZQX5MguM5D+TNTDPwUi5pW1pCTA4Up+04DfF9NV9/icD/wMdGUoDqP
HHhwLIbOJrDJ+UFs95370PZLjQvspKtmiwGdrUiCESKUQqUFbrc6WtelQB5E9KK+
2GBD8Kp13YVn7jVoitgpErT//h5Bwz8T7Fy1n8g0nECplMmqW0YUzeeLZycAsZrH
KZEzKXyoWazkcfX1tg6nV8qcp3l/bvVJr594k4HdhL1vnvMGvkDhFjce+vsO/bEw
AdlrWgwNf2A+YJ8lyJBMz8oJes6fju/rZ5jA7IyHABwKof18Z4eR0aN1efjfDNpR
HZvSNXHFeVEh3JXUO4lSeIiCszbifJz/lebov4bFdXdWLFVO97IMZXf3T1Mo/oTG
WmjPeZQ0MoSojvTK/jfLnDrNxskMB2aHkZjOxLV0x4inqxZL5HT0+9GMj+WZZ++i
yDo4DcpVOl85Qgb73BFUitecblHBuRdXgH4KrwzThvZxR4ciLuaoFcMi6wfq1BDh
UljnBP00deQuuhWgWf93O07KboPy00I359caAy9Jr9b29IOyJnufm73uSFAzGxaB
sAZ8zlPdggV1GOBnitDr8jPhxDN8kNimV814OdqttQjGDJSV0D/P0Dvw+sjYJJGv
NiBnM4Hj5ZJqDdkjxr7swlX5V/jq3uKUVkCpCYW1Y2vCtugqaA9AmKuVn1MwA+i1
kiCnLJR2mbdxGoWwoVATj3EMYEjInW8GpWakUbqfYzy45okg6iQxr9tb2/UP+MnP
rt6XxEXAKPhD1Cr7R5e0zW77W+iNDsxuIfIBPMd9Z2Fky2qBE/jb9gCbMOfyn9Ah
CCjXijDNLErvoyG1vKsJEGV3s//EL0ZbH6rhnAMJF8bWWu6oULu9OkCV6tk7uiby
qwM6R+jk1eMqveWOk+ilFk/bMEbxP+axGN1Tr183Bqa9MxHOUSr6DyKAA03uLfYU
7mD+3SkTuH0cjEXg2N5miNy8DPzOPKcVJ72285BoelluKq2UQPqN8es1KlJQAaaI
GQ8tOPiB89wvjh2ycX5r8Ch+fNHt0UpfKrmKQMueocguT5S2J8oFT6qUNjelOjfA
bw2xzn46Kc1jaNuGnUD9tsZ9sUic0NoHNh0ZOgBA9+0OoTJh5rGeaPf8GcrYnY1+
6429SjzI4CcV2nN4bADT/Curu3bG+XIyKoWNYvEGZCwePfBeud/xFm+sPdLZNxmH
xFOgrrtUn3xMr6kSzriQmXfOVcbcl8rwgedFTME9DEMR59cfgctrEsu8ycTTY4YT
OtpEbfj6pemHJ1JCHpdOMF1j32HCoCl1odkVjnF5fn8Sv1oS9yc7TO8v2qo191zb
rTgOhzSraNsIGuUTiCbjj3IqzdylHhvi7NkXwE/eSSPZYPxRugj8Sy5AaUW5kBrb
GXxAE++7Jz70ivSAoLx6S8YdhGrcW1SQINwXtR1RSkHZIA11GZILdoj4AcObkUHv
V+E0D9FJ2S+IkTM85AeWD0qncDP95Pjn/OEH3jDHi2pNCfZzeNKZfikdc8CdOF1V
VdtvfL7uBpzkzAgoPj+Z8X5iqUoC7n7/PE2Tu9zurj0tmSCAehVB9u6jgeezch1i
FVezQsz0jnj6vd9ghGlfh07QK2AJ2uyI4qGECAn4dheJprSqs+kRFw/TU0JmK8aZ
S0dshpZ9ztaK992ifP+YxNfBIu28H5rBOxoL8fudgNr0y+AhFfao6O+bmaNCw8aM
lZ68oU/5rvaKlP97owQph7BgO5fJTFBb8pI5FyLbraEfAOUPK/53e6SuqTCatpQm
4pbcARDNQdKWmwvGG8sj6R6W6LwqxuxenZ/tzMRIUNVBaW82AkuhJdfF5alFQZ/K
3wgpukcdQ8X2RFdMIqbbHFh6WcLdemZyP9LtlEFIm7wje524tiV0VGD0zynF8vfd
5QR3xaTUwuob1SJe9BYtJcRJ1hDlrDnBb+ccnnzc4/FVXuCHyZFuIWc/qwb5/iIR
vjBJe9kwbBNmPfDfS4O5R0aR3y2WWwWzoSEOR9vfq7eZ3c69jY1kgm8ViaedxwR2
vyR4nFHO+DZmpQ0m56A0zeTWufUyP6OpT0E01nqckniH/5d32GF54m5d99VDv3iP
MNbZ0QQfWIkCNIs8GJUWW3+QcdDF7aE6ShwGSe5+1rClKiSUHFVNsZChJ/bhqQcd
+dv95U5dBAh8jBJg80a1/HqjfW7CxPMmp8jyg7LoiUj6mwtl3lquRiF9ZpGjzzPG
dC0Ed3/Em4Zbsm2ZmilzfB7XaKMdSRSMnlfVb+jm9bHFd2E//sQU1s+vglj5FtM7
bc6ioSjHmrbxXjZoZR6XkHIvN01K2lfnbJXAvx+NO6EkCf2PS4i6Jgnj7003R7bI
FV1dX38uz/piElKnlj3ZxwQS0kQJag/kAwQ+Z4LbjuPEjAVjTzWKxBgOlHwCVep0
EXK3ZyNN+b3/IEpu5+FBfKfbAHaY8jVd2UOm/OIMw9QCRHIpaqRTbOCRR7SQY+v0
AK/4gHaNONeJ8dAi6GwgrQD48XoVCuDEVXnVq4KTYZ0tewk1+KCKoOE4+EEm8duC
MMS8TPbcPw/gjDAYGptguntoWc6Zj1/a2wr9JONuCs+A29O1+vru++spZuCpRzoO
pNPxF7bOdns/vMz/tK9FKq5d6jt9HPzjjvdByqWHvjpKOJ3Xogv3ShPAqozQHo5u
YG5e1u9reDkbsQ55mhfJP/R3KhELP/5K2wfFSt3SOiSYzgs9KRCy4i+Ku/VXMMzH
1Eltdnp1zKz9RWYPwLaFzXgLOKp6ChqkWsWX27LCpfqKgfRFZr6/+tivtE4cjKbK
ugtB32jWxlMq8f2QnKwDEC/0P/n62iMkQ5hpFONVCX0E/9S6VU1ICVE+tEjfpk98
kJDIuteEBAYEzsXh+NIE/Xt+MhhkmjnWxQ60Y6XoAW6cxsofYtZyeTkdTCpsfOd7
IlNfn0kJ44S5C4K83wly+MVxoQMdcYC2if7yBKr0pOusQGlPJGQxMoXzilrPxTcV
bgM1mJkksOODy5pU3o/zVEe5cjVFWWr7+GyDavRtdAaj3Y2kFIh2z62bFAkmkxND
xNnWd9oHsmhiS1Y20J0vWdtDRURw5t2haHEY1HZyt0V0X8ibqpn2ocas1lChBJoR
+dbnwiykRzCYNtYLDlBMekmdrc3yAx65xZBGEdnIEWt/b7vy9ThPHzT94qeIqbIp
D0GqAt3pHeacv58PaVEdaqR49ufIPh3oIrXJJmviJAPjHO9pg+lhK0fX/XHmOC4i
m52Bxxezz1FG9OuwJpjJvPS8ptnlRq2h3x0I+lawQvY57NumOWb9cmIZYAN6cwh9
jRz9LDRoTZFf95Z6mpizvgiYM21YJmahJYm78uQOQcpRg7ockHkpbAN1sjKZEc65
GLC3SWcKb0mFMSiTwKtgb1LmwbbxTrF/q9egr1o0sS0JMMKGxZyImlaOZtqxyEdq
krP0CWmL37yVrlmuiQc+Bq/dUDDXTxNh8oeruIsGQXukgIQ+BRXqS+3oQMXGasqI
5MLclyBHHZDfHP69jvcAdyNQKcFdgdvfqxu78jDYVVtj/5WwClfphPYHUTSyrPB1
EEsZsCxxYRcc0DhJjxzIgy3dRmbZsrPINomySsyf2F1ZIU7l5rZbcpuqaZiLKUmB
CZ6IcStY02XMfcZDb7dQJFSaYq+i7Pgkmih2VmnVkcQTMcfhP+I2aOwa9dKZCH4h
9hjbXDQpPXGRW7uBJXyIwbk0zJsUCNUl8kKvWZhidLo8FDzeNFuJMLSiORsrYIrT
pqfZSbRsCZT6sSjHgpKxVwtKPRj5nEoLTj9nrHcnt7ArKl3aUgeeN7KrqIEfFi4Y
UNluaFb/aORLZQOv+AhyDlD9cLkd8mczcZucafZI2xnXG1uUbzombuPZunf6V5GS
t4B13ZsjmCR78YVdAZoy1+xrAI62HUr2s4jhVoNMakkyoDzyWXp27loXU67H5cKm
UhGj8pcTOKwKfRZjJJsqMq9hph+p3QSxcCfLoT5c0i/IdsByMZOJCWNKKnhcR/0J
SLhq1woqspcvthN7u7PDZgxDV9O2/3j9rSYZUhQhqdebobLmjp6PpIuvz6XrKNeU
10BAKV7n5iuhJkIzOOkTYeuOnl29MXHcpUA9GrH6CricwT41XFch6x2sZle5Z3VH
ZR+BeF0eRcqgbsgNKaIOYWgMB1hcvaiHwW36ABHykkYH8JQR6lk08ed9f04dpXd/
BPsa+SOWJhv+VmE82KGBLgvtTKd2deT7BerfC8dxYgomaJVrrN4sEwIHDPWBavqM
BdHLAv8MpfqXaWHZBuDSfLHPSnLSUD9fRp3fgk2p1ZuQt6edhgGW0SjtXKVK5kp2
eh17gC71Tkg+5m2bb5wl0EadtAMMAyE1bdcNdf/7Blv3Mcr6agENtbhIPLPc53YI
IAlbyyEymA9KWFSURlzHJnKfa7i/sMhqiWhmNUHPDW1NpEYejAmxyxIGOlRDObzD
LxFc8TT4/AILow5hQ29SRB6P5wpyj63EGsOvQXoPiWX2I6vmULmLjgTO8LHfunlu
ZVz6Chg4PAz4/BzpaiZ43p9xJr1wtb8kSNvjAw13w7zAKjnsoKUu6uspdDWWqeWR
QHz42C2P5ViBf+gg2cXBuLuzkioe6gqDFypNuAHKNidiOny0NcP20GXcb3HxVMBk
9nR2sos72hntu/ZHk8Szi9Cf83J48lyP5plsNUFQAKi3lQlfyuBtBLp4vnnrj0lv
xy0gD/aXc0e5F/kCk8cZKKLSKxpoe4CZzvlytRTRjBM45UpUE8gV3CuFJ/zuhDxs
O5yPeA3uCyFF00HaQUIFc7TcG0pGE1yiiYouh1rJSLw59T91tsZaYyKO0+1K8qNt
OWiy6XAKQ2OZO9vrXaZKwdwda3aayXWvP3GSNBKUbOBp8dtt5cWgBkp90hxqwtZm
w5JM5/bLAiflYI/IzNAlGDNans+JlPVWbbRZcxPXeXt7doLXyfTyWgv0a5kUkvnw
+Z93Y3RFgBQ54Lx+axQmk/f+GF3hCcv8hDCwsstyCYY6G8EAbVIvJeqJnSKhlzXG
PmuCjk7b+YsalIDAf3dyi9yBayHBPrjHHIxqMkWS7SiJllbQTMGRNMqBS525MOd7
pJ1sxA8fZkNiNIZWupsZ78HwLMdW2MWc0+kwONPWcI9aiMb9rhD9x4ccP0kypkX+
UVpz+4bkjcGdyjdYer1g+zczYTf2z65UCLaVBB1NM6t8mxwggYSJNvR/I2fwLlLO
haYO/Wd90krt69P0MqXlF2/dr8A1Xnhtq/xTgNcRNFiu7flcqQ7Xk7TrzAhmX59D
vs1BpUmgIhel69P0CQiUWKhL2ynSHy11qPP7hCeHJM8vxrq8bW1eGMNjg0UwUh4k
Im6gkS3K3ZIj4y9CDMrWECPeOQHylUY94fTPbj8nE2Nl6xqK7Rl0/KIla6udN7av
6qOKG0UNaTPNKeGZCA+Z0Evm81c3RcYkk9S02kvoqRAWyeiod1OgzMM65qsbWTVz
kroizKPodEEAuryMZeZzrjhq6J7I0y1s/StDcxM67TD3pKnumAPB4hpuMNh/TRVs
LUGSJyRgghu3F/6siEws3M/e54jE1FwiatoIXamBNQkZDADQgRfFtWcfJM5R+U+5
SqZ6lgW0QSOI4Mbnb8EO2NW3m1dKAbEZbTpf+xm663P89a6SHRBopRwXkzE3+BzZ
KFMmvPpUy0VLoqoa0Wn8o3XtMwdy0dXQT+7p29Lw2wK3dF9G46DYueJafsP/BI6K
2DE1EB8k1qEQDD9nsNSyuict760DfBXJ0dhbSqsJvOewWnBXmYTkrarEnq9Btwpb
AX2dl6cymS6QFEjiPI89ruAclSEVDQZcYc2nKCCEfvFWivt0LNtugCl0QEhkwE2F
z3mIJs8qvu7UtGRI4d7mB7WLig8aH402VFuHqZ5f9cLXnUMSYg05eev9O0DEDhUn
mzyKIMf/+BNDQjvJPPbQ36KX14A4W7y2rpUq0id4693FqonLUAixntQWk3EeI57V
sNeu7Xjfk9MfOD3ydXEf71EwDWn9tXrOjxMxSZzrsf2n5eJKTBEZsohK0n0Yfwdt
NUs2A1qEq12CPiUdinMPnswkLfzgSyH/Dhn7WZYnsoLIAKqZFBmrD3jb0oF2PsLE
3y6dMhBqrElUdUcskGzsRu8UgxxdPjE3R9ZCvEwKvmlQlwu/PsJ1NfDjX4jpqi7j
hSrhT9VCJGqTaiAiWIky1lJOeIWmEwpuS5RjZynkiDyq1lptZCTz8o5fKbbabDrI
1MB6qGQakOc3IUFSMkDoHgqRY4pAenfVwvxU73wVM+mMqr7BhNkGo6w4nUZPGhUx
IY5Ge80coUnq0quRWJTAPS+u9Tmos6ohG025ptdbbF6S+DX6lvN3lErzwjIiNzuL
/JCLdSXQcOw0+q1/UkxoAqhry0TM8J0ob02qq+G1OGpbnslEEBVl5ElNyYQRUXuM
Z9N/5+KhlZov7c0We3A/hL2j9ftEXArecjc8AaSA1tIwzgOuC/CFTEw3fvPTT091
HiRw3a8gdt1BuhM/CRBzVTuH+Dz9nYeiWtU+miYWtUKg4Fg3eXtOhWLL2DnjC8Pb
3OKHlU48qCDd6X0QwmZANM5Kyh2iqZ9XBMmal/xXUCOILaS4AkZuybboM4RcAw5J
wyMG6YZfbcWXJgxINU6VdrcJ0UpiOYCvAfqd5UsPelgPMrCYsqmLIbcm3ov54F/X
cJIqI52jZmHEo0QTabkcW2/iOFXLprWP9UGV7enyeX/8MrHrarYfdHUx7Xy2AYH5
TRJpRMo24xKGedX0EK5tZEgaiGVJprWfY5A45pKd2Si1OhCtMQf0DCLSCJ1sDZbK
w9NoQpnS+UcjXzATF8EdK1da6r89QV1CW9AZqxAjpa/jc4V/vfh9WlbHCVRYOXu0
oEmWgEUKdqE1Y0Fb35OgOrg6hQ6fXkRNbpr8Lt//SXbnWX9ai4gPXXbSEAmiEaIB
6ZrbSoXMrmFpokoxGgQwVIcyBQE0TFa9jbTGzFKxRnEVaPDBq0CCUMjs/wYevKf3
6u54bnEjXH2+XFKXY7RxlPSofyHDEKXRvugk3q3edZwDQuAfHrkkN0wRsFP0nzUJ
qnIgynmhUu4tM/EYSx3YT4BZr13sBf/q4SjHcA1x/iKJcUTaav0A21WJiXXhUxWw
rB89e8899JtUr4YH80QmhvhIdQ2C+SwvlEUxSxsu2I7cmp6xmfjFJrPT9aL0M/RH
phXWJR2tGIN0yPuQGqz2nPUCzfOS38WedYEivIRdp8+rnOE0t3ka9L7iKVq8md1v
RQeuIYjGZIR6vG5yXfRUc0a4riV2s0kdGeGto4dyC+07en9IWSSCdXJ33Ek9Ya6h
2SAHyoVFJSNzZuzp6xlFKuSdfYNr5zBKrq6ZZPRSD9ZWpO8nyuLCnVSq2Fbe2RGL
qtthErvrYWXZ1lfnJsjNIT+DoM+DUce/lCxTez3pQFadi3/p2WdEkNxDuczcZ0B8
FfYNMAKHeufxnvi75/0zsV0FQywAEIpI/sPhv0w61Kb5/7/ee/qBaBXtFSTnDkET
tn03SfMKNm0B+vPdtVxZYr+xaX5Lg3xs2mCyUewgM/jnNlGaTXkvCk6d47Ornv55
rKNcSfvqJr5Vrotrf420Z0FGX5oXC63gmZ/fy4ZrfofD6ZerH4V39EHatb/fd2lM
jhRMzdU8xVE6VEhxQz+6LVL7glvFPCYiiEvf09XYwPI5faHt37bQABzjKuAS/W6C
e6ppKJlGPKQHqN8ZFfj1I7JAHZGFRRwV3LghS0P7Qso7iOQ9XpGb53Ly10NQUDSF
m9tbF6/wA1oIqvVDq28ZHxb1v3wqzzzcaMIxQ6UPpc/U0eHpOMgU420i6gYDjU4Q
esTDwxExg6Ly0mOI0hsXiWsdKSrpBPNiMTc4LOkKxVO0A7JMAGvT0vagB/xhjifO
rzMj0+TMDBcc8NlWJfcW66kYVYscW5AZJNYhRhbCwuqlwjzgGI4NGgByPnJPCyMO
V+oCmsrGojLfW+ciaaodECGVoIUvsMgsLYIjRTBuBHSVomlheSoykfs8WOw76e37
yY3Y6eKMyXcif8QGKTBvKFGoBrQIGxJXX/f7D5EtW2FOXPhLZ41F2vbo4aBpyOm8
I0sKKjw6ic5SHgSfzItudoyX2SQAaXC+bBSPSc5o+h6di0RC+21sUuYT2ybs4o/X
UE3x+R7gvv27IQMrb3xfYvi1XKOOK6Lq5MOGK9D572WvldP5D1Y7Zm+rZFQjXuxG
MlLpcXhWM12HthMrulBQq5U31MhUi2W08myI3Vsk8Ftcqr3lO0wH2pT00L0lRTZx
dr3GjOtj6HPn56TaC3YRhl+tS7y4KTDwTCuXH706yJw2ykD3bA8wQLtQGEhlGwVE
gLPB9zHEUg3Lzc7O44ePewaz6Skbnv3zcEilEmdxB4dmNmkb7IU+/UAK9A/VZd8n
6+hidj3DkRWlWbjPFS139O+zQ7ycugtrVgoQp1rbMwqhhl8KQbdjSQqOFA7Vs2eT
Drnf7DTlIR2pGuqNkaQadN0ZFfKshFi0qSxklFkuB+3ysNtnrnzKBQF2+TUYnJit
zIMdlbRSznMdr76GLK4UH+2RdGyhB3/LAthIpE/94OthVKpWlubAkIkUuv7Nk5Dc
cMFMB72fug/aBDH88Q5epacSZEjD6pybvpXPUXY2vywML8NebAb/gz4PUMNQ70HN
0r1zoZNkRfdwqDvGxEXXEA1xcJZiVW6omL+ieipVIsjYlPGpuMbHYGgNXcvmgL03
Veoym2J6hBoTu3ERkK+6BAU84O4Unf5b0IUO2l4O5Ahq/bIoZfa+pMsuAFBcQ0hh
AkcnMQ0u4Wo8GMlhWZe7+0siUaiDX8puC4WsPff3fujwt8vboMcImSIPME1/mb22
G8/7d+2rKOlKvd9CBoC0jl7JD6kYAkCAyZJbM1u6kXdBEayWPLZQaQVj7k+Z4jSw
IvIPg3NiD/NlOKT297mvanU8Am20bmz+bTZqRXDCIPMG5N15e3bK90K6+fRUUpTp
+Jyydw0qevZ4vxdqrRqk6CFUhyQheeJstWaIdhdodk3RPD6/Y3/IDDHV7EFCwFOT
yVHBLZD7NJHxyqxUWoYJ+Vhs0vJMSAc+fCuQCr8hP9FEQVP/8xDeSCUpdTj+5xLG
mMMWyH2VG83i3wJQc4jfvbWp10otgLaLGctkwSv7AS/M8+TVoEV9KpR1TCrD2Apa
0Yw+5p/Lrg4eEOhKlMiSSyoHi+eu5+R8YFUDCnnyuT01QuK9mqVCoMgpYMGDpnJX
tqLqAWWgoYpPto6oWqpjJRfGCE/e80jIuAe5YjDj0jaeji95Au48XegUY3lP3p8Z
GNguwsSZJR/Rbcl/G/UBhIYpREZdZeTYqMNNzfxB1N8WEbwQACfdk6VyFKzQFvFC
NpULOE6PNQENHJo1862w12OI4HxrWIZU+QDQpilfQDf1Y8ntpgeeZeuka0qlioUY
XlwfJ2NSzG56LCs2/y9VWSgI2pNq6stUMGjgBxmvl3XZHcJBrkVeBMYFwn38C0av
A7XZ+deyIC4ejBgezGDwdM/o3x8rfiF+CT1J5B8R7+jopmDr7pvkOlAZYoqCLaTI
+JN6e6jKn9luIQMlaeqiPyQmpUjlxjFyyjD4MItA8pEQZfyw8/Lu/yjtTATGscTt
Y/fmqQMpJT57/k1tUdZhT121kFdjpuaC98K8qSZcQGokvo23Yhf1bE3ZokOyUpUt
oiHDMWH/94bZmt+AWqe3xCLYMIYu8PQvdJ1FS2ksaCnCKIsbqB7U9Adn0oN+pfPO
R4T8Gks0XCnbEDH8zI2Rt1jZuRhywy5qZ1jRpi1DZItGK8bUJHg31Xd6QdIQ3EEf
ORg4TvP6RDg+92d5qjTWw00FkZNcFTZolH6LA2wC7J3fRbVZ4jBv3iL0PVenTDpf
GStMowKr0mKA3VzZFQmqIg6oF/6U5yJkWeQSgg+c0M4A+GxSiaSldYhF1DSjbRWL
Smp1DYJqA2XlSdLTwLVD9iWGJGrFuII9fy2R1tNmjNbRt6hZuT0OIxq+crbQ937P
mbrWKpfPU8EKdNzgs46Qg8i6VPv072f838VF+otsDZfTItpf2pDNzI/WRmCoMRmV
L2qKgPheDFJhSG0t8oGvZxG1wtGOh0JsSUeB03NHmqcivbUBDtozVyBco89Oizco
pSDwWHnUM+2iNaQEGfSNcLVmrtz/wFX1e7oG9GRyr1RjXY8ewMtGTJCg/b6Z8KZT
qDxwaM/tpDQRDpTE+9yW7wzEvd5YvXavaMuGGV8Vcy1r2xzGSjOeMmDyd/rvUNEs
wBNiUylgYH+Nrd49m4PUDNtdgCEWTn5sNCg7bCbNYwCTN3JEAGLh88AHUJCegLyT
8RkeK6kNEzQsLVtCA6oJF/WkyesMlcuRFhTfFLUTRVJx9DBoHyAQlJ7mTl2ESbI2
q7h52Qa2obtlgo/fDah5B4lb2THJRQW37vE/24/5J+hmeTh9p5uYxVbxnkOrO3WY
qrHJkaB7QPpeoRcvWRoL/1ZuDor4GNRg7kViUCSIwzxUHHippETp8dEAalMKFPWg
qEOYHDkyrD1RlkMzZGMvJz6WGNicIGkTBeqqbRxx0pd1hAM7Oq7hpS+/lE/KhUJ+
TnAel8D9XCqDDjAvPOzE+SwH+hdYNDw71xzoHxVUy5Q/Yzu/JWdu8GCwHbi/xCxx
2mH1/iAPuXgWeAUh0IPJ6u1Fo+LqTYCgk+q71OtNzgUVoSgh6i4eTtLDd8YtCHEO
Y6eO5wkfZxSRp3ikq8PSLMorHbigp/jR5XFtM4Sy4x1JeiCOUszsbawGwnH9racJ
usZ2P/ohsUfzkPgsc9yhVQa1TI+Tpf9UIo9SYGNP4GEHJH0NtafV8R7DqJPOO2e6
CxFQP9GAPHCsfkLUFdpbAlRSrxWHJOTV/1y0FJ2Zn32CgUp7LtO/2xs4PfEVAECa
kSIWpYIiFSqSL6xVNP4WpQiFeWli3hYpfzh91Toi/BO7C7mnlfz0YqSNsxj6aRiU
2fWXAXxzpBCzRQWAWoWcGI/GLOl8p0duWbGTojYk9oOo/0VOS63hIGXyeKy1A02j
5PKCZvg5YzclJAXeqQeAkzOhIN1waSXZcNv6AWlqzI4aHHW8oyh8NVivrvuTTRmp
2ZVkwqyVwmUVEHjQtdAET/TMmzwd7JD47nU6hs/XjCMknhi8LMZ1Oau9lnjnky/c
ZM2wxADdvPwoav8ESOouolSAWbOWYGKsGgN8xYF6z5siPgwErL0A9m+n4smBKGif
oxfycXJWH9dascTPT4t5baM6W3fN4m6WOKu19TQMV8O04TtXysv9H562NgCONw3C
A2jcPfolKxN0TvPsxT6jlkfbef3UM9yMXNN3Tv9G+Yl7DABEdw/TtHmLXCdPOuoO
0mhg/wC8ZZ2QYIeH+oOsrwisMBIZQOiLjIM78OXEGtwrPa8eshe6Ekd9LA4D7OTG
VwP3sjQrYqGA/hwUpx+zym/igoJGBUPPUT+4lnqqXEbElny81p4glxRf6qzIhD0E
exaNtDhoiNR6h6IBsXjW4vBqp3a6463KA6XOICY1QCQ7KOHGKCrUTgvH/yDjWVMr
Sc1Orelpq1tcA8nmUnZ3odMJ+/IV4OOEbgEYPFdE1hpjs2b0nTwYT3jEmg4OeRmL
NNezbmNaS3ePoRo8vWzwRV+Ca2Dy/Zn2bwYfyvSxaGzMARNTSq1yHnMN820ApaIc
XKdfTbo/VlgCOYlkY0ToVaNSYJgTYoLh9sGlcpF11TOvqf7kS6b02zD3bhV2t9aJ
N0O5kZHmiao+PI2iZ0CT9OyFoBnRlQdI1GzHeH+2VuH/HfF2tqHj2L67ucD1vFXn
p1t9aa58VDPxsvgAmlXbdUWUIt99q1Ip/mf9LF2ksrWctEEMFGliLP8daJuHmMl0
XpHy2vOC1RV8/OyNeFFzmbnN/lATMiPc6jTkMSDsxdjhDqZsIh+X4XtGvmL0dunA
hXzx7NqopD42OPh2rP6brS6ZUnMQPy3qUP0yW8ZsKUaEfWV+3IhFtCvYTTGhAWxX
4K21vTh2Z3bBv/021qcP6POGI/sTpznSJIec43RCvW7geBqEjBxA1xIGqJKsVh7E
P+5vFc6CmOyriRlYmLoegRQoOaVPShooaTa6APjNBg5q93uHD/35Y7hGkiEkSrO/
sKAUSYsl27de+uyX9zAHW2dW97yt1W5EnRKfGt//BOaPeeaBDEZ0JBxKciziWRaB
LG1hyF7hDpY1gDUSOLNF72EIUW96d9rJ4FUUsowItBBJk5dm/EVaJxlD1XcNf74b
ukqnK54a3hA3CxeSQ7W1rPMw81pPs9Y1gSh/0+cawn5FNVg39bkyzr6VGeCAzNBe
yx9Qd9MyQ6vlEQu4saQ68/Cc3IVHLMa8ckYP9vugW9IgaqXFoS5u1r8yscu4756z
F9XROKOmeQbYWmL/EM2EAEaMY/WFKJ4xEsZ3Pmil1oMZ372/JbPbNRaFvsm0FSUf
MfEZuAv/SD5IURzy2B/iq8IczjuYmh1zFs+g35O81wyGIi2f24l8iC5JJHhgvtAs
a8DmHpP+NnpM60paaR4t7x3DfJrEvnytqHMKmQiRoC2QFAO++OOuBj8sVsXn7lin
MxdMEKQ8lC9FbPM50uH5+Lk0FMrujxrMtH9TgKNEWbOS/hgNAUJH+wxiwGPN1Asg
CYn86ocYOYuX2NEx9F1toQIoDEIm4tzeTsnnqR6ZZsAMb0P6p4dk2Or6Bcs6HSsH
G+hjBcCIcq2zojQusCV5D5dO/XDAUno+6Q4sfzPPLZOAEeo+J1qfE2icyDsQdGvk
nt1G2yjJg4eK+hNJjemJZ+zKd57L7UBDlMDR/dYGRMJfKd/CEW9YTHsFT1EZRaNf
rFVFDdoHOITn8s5KybaQpMT1M69QV5tDy5UkVDKSLcQm2LM9xg1VTF/h4cJzrF40
T5lPphder3osWCU/RcJTywZJwgiM8NV7X4b9/NIgkAX/zJgHslzm7UGKC8O/IU0P
jF5lMhBzwHKRzC8vJNG4QmnHxrERBY90onVZnE2eZUBVnxqJVYaaDKMRRD8EQxEf
Ebt0BYud+xkTMh3lyoSfvSq+iM5SGsamP2oKhmUdsOXu81JvfRVAn7I+sld3tTA6
xMgZJkKNNj63dYGP6+23ChjBQ4MFrNU6AckB3d9glDxIpNQmPhYpISf7EUYU8Jvu
0j3KpR+ypI64KA0a9UUmglJABseUwYFv2ijKwH9yO4bNk7vH7jl/YIXPTka0miCR
4w7IuHza0SBNJHg/QrY2kPWJYzvbyZhvuTYBH7vO46SKV3ML4oVYXkEykgsRQTih
31NHzyjFRZvDaKph7cDxu0rg4tXsUsk3YYjIVrFiwyR2f/K3SNA+Ucxfd1Wr3fIj
5/p2oWKI0Kcoopfpoj+cW9vIYp/BiFfanyWCubmix6y/No8iKwV1AIxR5vzBj2Cm
m7LhbVUFePFUq6GwEXT4PgXKuw+YLKpRnhy1vEDBnZ1EcIKQOrCkIPUnWU/jlEMt
WcofXQaqmPJ532kfNaG90Ow2HPoREl4vZE08jhgXOJObGpjQpXGKt1Ep3aML6+ht
rKAfUTGXV2NGDqFspYD+LJyZC1XIok68LLXP95Sz7HGaLjafJUGBcgqz4fccqNR7
q6DNXSMziWF+iHR3ZS7Ijt3kLVuHnqbYkMJTzjRIyELqZ9+si62fQcff7gzAKd2v
Ev9cmhjmivKPUqdcAI+7R7oLX1N5VzZZpTAt0fGtKYiqyPlzsrWyNDRYx3U0lQv8
8pI8OBFtocBaUaJc79elV2rY1YEWF0P2V6zV4cWCH8aaO9u41DMoC6rzDgzdDOLO
oAZNdbe8BAFi1RDtNKct08VLcWTbjInYw682dSEUphGklxwxIhv9/9yWcwQP+Ayq
dAxijIzqWqfG9daU5n6xgB/kP0jWXVbHgySEA8KFioE/XwV5Nq/2/vYq0egwULKw
8lxzWsRyMXjnGmy/Fw922sdL9X7iubEUGo8RCP9UwHHjsoUgIIagAieaTJ3rhbDu
28t0zs/NJZNS2T6aqVRTP0fQWv9ly3BZg8UYM3nqW/COwsIir9cm3o8YzxeEavf2
3N2Q8pw52JpRjzLpbTU8dBBEjgLF2X4T43aqt8fRBWWoZjOtjQq/+XWfumQpSWfT
g7s/7gshWVogUNzUmbWHfo2nfaXSax/dqtcrnmviP2Qwb1qeWYEamg5QcfZKTAsX
wKN0vs3t3C5KWCrYYx5DSqPXNl9sunkZjCFGqqHJx4gFEs0K9eFnHZ/cBNj0JIv7
/kXy+m3yhcyHepTcYV/vz/sZnbENpLR9qZx9HDlZKSODSog5AJIFHZ5qF5PZ4KJB
x2Mnsvkdl7xtsAkqrIgjH6QFcAqR8p6qyFFoitbYHSX27hcQbbrGEHYL/LcdYXu7
iBW5qvANNWom7wzxuGllIBD+g1wvcRvy9NQdjFw7XLYcXC4hgz/pnV6mTwnFyIgL
seoO8Hh1cyOG+GrBkpQMTcYHyYZnznMH1xKDNcv5c6dsawuZ34ypkVASCJcxBm1x
6LntqYNog8ZqA/csSISKu7RjZWLD7+0oDwEDYv40olDmAJfvdVKz6GDxQMVzJvn8
H7eZVJKvF6Yv61luY4CgTKVOH2X1iwlLIFgJNurrBCJdrKUe8I7qqcuScVv7YJ9G
m6ZphTk7MYeu3yxrgFWg+R+jPPi0L4a/yOp8yn3gZizvbN3deNfp9b0P1F3yQliS
DP073psL0+Nq04Qqex3jlQDbUj86eRj65W3sf0kjrcQp0JVbdgRYprlCO6TA6WOa
lXuouq3SbTPP70iJjp4FWG224dY0f6VxF/kIpv6aekB6Z9z5hE1Wl4krABsf3l2T
F8wesTlHnzIiBJ2wDCXV4R+L+q1tG3HJoLN+MhwYE0Q1a/EnEVcf6nLPPlM4nZQ9
br7SvMWkr3csKgVft+i1iREtMuDbAFCN+/CZDNfZHYEDCbBAzLN8if7tv/r+wgwg
rcGbHOJULKX5pryidUAHhIk/Ipkp/o8imE+1Za8BH10VntHYqARav8oPIEu1twcA
ufvxOA1xiB41OR5M5PGZ+FTf5QBsF8kuYgOKp3o+n7WS9s6/vzbcNnXnULKRmylO
2utEe7X0cx555o9pr1Z3yUoAuq+XBKX2DVmwfhUi3JOnoVuAa2hjrTFsfoS4aPA1
DWqJHpCuxx0ZkrCb7+koUPazuI8A7fztUIDhQGAZ73ej/Hvv8BOBynzlsIjLhcFt
y4Fa7v9VHL+TOZjpFY8iCMKOok4+MQXP2rfUggyGzes5o05pWFXM9dMmpQFfmKN7
mNv03rrw+21N05h2dYcb4qOZwfSndU9U134ZoeKGQ9UOy9gu+BVg6fh6YXLMmTln
zAVoOQS1ygOWZ9VoV2fSQd0aytfwFZChD4xyS7Abx1TTy0ZxXdoTQ+6bL/FPQfh0
H5ULb0K5xtU7rTnZHPZ+8weryENc++cpHWzUMx0O6qOtYAmM0pIgLwTkbstzTbUY
iAkJaiNinJYfXzERGW9PqAyxRolPGyKnv+XB03GZExJIMVLmZDsczA2uP9jY2FTS
Qhfs23eWc7Fz0p2D0nlEA2KyEPN3K/eofdovCFvtmlfwLZeNkpv1x23nsmfzFv69
1MSVkhtj6Rc8mBwscs49A3zluo18Psb6bE22bQlGERBnJobgcFu1tG5ghJ1u8ZxO
x8miiYiAX/EHyX7EqhGva8cHh/QEtxiHVGNeClfJJKCqwKHKE85KEwui0hF0Y95j
Bpkshrd2bxjDTYBvhph6jRZlEZ2zT5/WzIOIZyMOQuPqepbkKA7YqQw9J/0CCG/a
WiH8u1lC7y6zec4/HI55phRzhUDTMBjEB200ucfHxyrBn33QldriMNgNIDxv5I8U
qT0bL0vIUGNFeDIjxdfvGMdbg0cQke+IVbbAGkg1rMTAIid0ZaqTTA3gRTpPJefO
4dxNxsvIl1fG0cDvE5BtchtzleW1pt7tGRMxgMwmn+dgIxg9mfaQWpp6v6EVXCeR
vIQoUkvAokh+XCPetl2IO9aaeuHgV6Odo8lGGJZqnzqW3P1OQsqHcsbTCdyiuPW+
6T7U7heKcycbPgUUqi3swFRkPzYpxD900oKsQqOLpbE5J227U7l5ZPNJtkGXUaBw
BZAQ4gdh9ajycZ8yR7tMALKSCJ5ptA72nwwpxQLZSLXilK4lCTSc9BjO1qVqbMuB
kqvCLolMnh9jiSufjju6VFG/4ZQg8YXnrANez0TIonf91OUnpOak8fHmIi0Y7mmq
AGqL9mjJ+LhXBzJd7fB4uvlUipXzvZsdi5zI8ai8lAT5AiZ0W/KUU5+B8r8DYbP0
Xq3ruIplRGb5c9+i33NhETdYPMgKvkGwW6QB3QR+ZYFuqFCZNqoP9jESg2ODIv08
Jpj4fNf5mLEEIpxXOYgW4G8HAziTigKZkMJIGGSwSvPyF44SeUb8uTJ9XwvTllff
J2FlCCkVKdapmw9p1Kab2VB30+HFNc91jQ1mr51pyGGyItR13lm/nO5Mk0bc1Dr8
AO9wZDhDVIVck59Luvn1PuopF/tRcPLJDrLj1+LqcK2R/dsyO2AaiLavOcSYDz5B
k4X0fzFUZIUwGzMUqpaGcNpSYC30Ddn1T7T4M7x8eCH54RC8SRIb/xsG32eEwufY
nl+1kq5WcOIFv3mxBn/4w+4Q1KYXvTmCl4B0N6CqlrnvK8UxV9o6KytRePtR5brg
h7Wa1ux27lzK3K9fkERrhsN8oDH4gMhPRMcuA6MAn6WmT0x1J6seQd58fwTmUlVa
+JOaRDbLraJwUezR6ieFfiHi5YWJg78vsInroIZ/X/e64YKPb+2FEF6o+a1adyQN
fXQ5/DHvFV5tpHVgsnsH2fpHDXdClNw9RDaRWn3nILZ2wbkqTDyuFTEkuhptmcpZ
3Rn4S9V7OovmI82IYx9HZZyflLRQunrXrpH10sAzCFft97Ju+chTa1ENWa+6sEso
rJ0EQ+ML4WFcV09nje5jZsR3VdtwPnV93/084Ki9ieRmNsqpRRkOhcLX1xr1MgoS
FsVXfprWsLWr6rwQ1jbCrOBGNBKIXhQ2ZH4L8/6jAxpBQvMf4xSjSAxlx69KRo7T
2juRI6C+Oj4G0oQxVfYa1uX0yeaZpPJ9LQglqKBh/kHhDtdIa9ZQl/w4EbZVnUzq
HFbnwf/MNKGZq70QYakWd3fdoITzPfgEH/FZhY47EvUV0943HsSCYEe0V9jQg971
734kzhUsIorjxKtTVoAXtr91UDurwfWDVy9eagUv6NHS+o7xeNSZE2IidWaVwnxr
ldmNgvw3oQ+lY3Q0SMR0r7kdYxt1Htt+qVlqSDzurwxbo/FWcKy/83jm6d86Sdxm
J4jXGnKfRyOViSrzmvi12EmPUUAaK3YsriuwBcuOe+ZNgHN1AVYZuLVCY07ckRDP
sL/QxbMe7ePEdv/IDNl6+y4mju0cGgzjbpNdA2XxxWBAA6+E27FQv54REMNfAesA
k7eL0EVpoZe9yoRnN75nN6XR9vvNPElIA9yfpskQ1zMWbdFJq6FBJBiVacBK5t7y
+jKhlSp7MOiuq9J2twgj94hEHqUioXSskOfxy/jBWtDPw4C3Q7XlaEP9jhlzX1AV
Cauh23CLrSpVWZ8Q6Ptl15Drx41KuQKcTTDLY0hvz1+X0D4/aJd/cieu+25bbJeS
9aOYZaRgEJhv7riw88ApCAoMdOzlrhCDSyvC20ardFoH60PLZaNdtrwHFupiMvVc
Os1LWR24SCZJo5vR3ojYa7rEcSlErdSY9z+diP7ueKp54VW3j5J1C6/Maff8iyT+
0jKUz+/TKBJUirdp1WDt3dFA46Jx2xxnDMGTF3E081sZ4HIxQzviayz/UkStssZZ
EwGnzttu6QaocQTy1XD4Hpl8h87MXn3BOPd/wq8TQX0g7grT49zxcDyJyOWL8W6k
1mW+8EEi1PgW0d9Mmjd8IIkCtybB9+JAfxeg+YEeW7NVEgrHXs8AVWXU7INJ//pz
X3jNdeLUd7ufgsy7znyu+2z7cXhn3Fmtw1HST3u8GY89I2G9AdBC68NtEKMIKriw
4tvvD4PkQ1kbTi57oowhC6lrRw+Sz6jk1BmKWPypcMvfb57SQfduDGvx8M7mZqbw
hLw8esY5U5zkS+SdPqk9rg+coF/GMhsNlg3e+QfS4X6OyKR9uLVYb7yACOTCWftx
ozKRH0HTtLSqPHJvcZOVaWAMHl+30VcvnGF93nLmqiC+ITZN06Pg50XIcTDvCOYA
12zplzk6jRDdXCC/bKmcCwe82Jvt3uinrkY/jjiKV5AtYQjfGRzbxGo6Q8Xcchmh
eyHbdsdmncPYpOSJhe4JIrzaouR11S7DGI5HNI5ZHvSDLGoG7yoQNqdYqqCPAIvL
MHG9lnU79sthc8pcKhdZ48PmkLfbEvKNEvB6goVkbEFwKiYFKnRShIDTGnqnuzEk
MaHFZALy8yGLe+j9WFHCe3jq3w3b5Kbyv/Mk5xBqryLAn+SSju2mPq5dME29h0yv
HsamTp39Sa/mYuIzh3Zq393yA8Yhwy1sSmS70032H+kUObwKyENr1Hoh7MXiKikC
xqtYhj3Gf4bSMngtqGP2FoC7S3qwXnEjoI4AXgoAVVZ127BIj8+6otTdbfjXo34s
ViBCPDa/fwtpCCvk9FLzsExLi1F6ydRXmejGTMFQPRvuMLnFcBnSp2bVeBc6mqRf
JzE+BoPpfSejnjROqnrfhiK+thAd0LhTt8araMrUW2mQTzFuD3I3dHhM57wgF/l/
FRw0yg6Tmi/wWOQW1bjhZg1/iRY3KYebUVsGYcsd2G+S3EKxrkH+GNvUB+vuZYvj
4N8YxiMXunQjAr+vGlnEyWOXwrafkseSlNmjrKEdvbGgjSq2lP0aZ+ABpltgJqVJ
m2mt/b0HeAtd2VhsewYx34nid6n+9b5dJKFuCI7VAbjuXRmNjdCtmfF17a+HqTXM
7FQa15z1MAHAw2DSfZTi321l/TIHA+ZAyEeGQUVNvS/z780Zq4i436aVKnLNTFsH
g7ZOzWiZ6NTLemldpUCveFpWZ6XCyCNj+Mum63EasaV/70LM0S9fnJ7I9gqTsIRY
Lb7+XtyUgm+8HuH/I2cHRUIMLya03BoqJiNYnqMq7wX/WxyxuuuNjHeS92jzneoF
uuBSPfy7biWlStYqH0i8r7LFyFTY6TQtTojtgMSDOJotNKfwSyoSuhGL+uvIdWXQ
vJGGV2zyfhyaYrkXiCf9NDHzt1bYWrXl7ybDqheBc4xhYGAi2HluNmO2vD/NTwzS
FRPzu+QhIeGmBhNgqWwkS7F9wnUD9+cZjaeicq4Kn+sH+asVKlxqoHpGtfanJlv+
zdBMIa2GvDPGIaNMo7iizpHGdalmjfmDSi2NQe/U4kRQ2C7Vsh0yw3B/49fmHZ5Y
gI9v9jn/YzJwNzArvid2KY+Jw2X9TpgxWecigu7MN/3AyLEcoZJaAWMPZc3RlX79
HaMDsLy7LxoItIs7/DSJPUAvCjWFbMcf3W5eLW86ETr+7dmVGS7yPGtg9qdwj/xJ
b/TrerHeoSGRawzOex0ec7nW3Norras9c32bl6T9BAUmzGpMuhMFYR7Jvt1bjHVF
vk1/Ekxdmvgo1B2iLhZDY7u/G5rZEF0rvto3NxpGX4bHheU9ZC+yIrl5WtkH+Zu2
Qy8HS0JS5eZmuXdzqSPhLNeQBCmFNSP38LSKTKtKwAUsbLsgyVgNpw56n2dA1S0J
/y84PwFu1+EvbDGwhulzDo7FrlsnnucWgu/YSXxpnxj8KqIzTZYRJ//l5mdZVtaq
In/UzNbLGIFcMLls+Njxf5Vg5x/+JjgsGIsuwW/YJW3G3TPZGNB4GY+N1Z1p9wWR
7VOlLkZGFWbynluWhjlsiv3wsDGvNik/olMz9ZHoelLi6SO/CG5+UG3VlNZa+xiF
EPQt6z32sKI5eye5Zaiva2UMsGz42b7798u14QJIUh/cxmRdbOfSg424SSIChq70
QO09yTzvef2NeAY39Im/VsjVTc6c/1Vpr7S6I/mAbeEuhG8D37oWId86ZEhIPNKE
2t2147I0J5uuXmthOcaVId5qUfueKcTSfTViGg/6CV8lmQRMz8im5KaZ52KsJVuB
6oHooTPeU5RLwZBYQNVL+eBEyhfdnf8w5/b2PsU4Cy7/f44j+Y9sziKeO5pHR1d+
smiuJuc8tYRc/4NpatZIkdYqnQtMUVxo0ofkrpoNReKsCTCLlUEjpW/nK6bm2rPh
eGYtkkUMyiYkPs1gbypn5AvK6y0Ps2+FWXCOISzMmumuA0Q8Kng69J97hMX+X50y
8Xn4b6vkHVb6xXi98d1YKfFCIuFZ1eUt/pOD84VakWUjve0Fbp3blg6Jkc/OZcTL
ejobM60RA+lkX114UJBVUq8DRpXYeYHte5rYaBxuz9u0RG8xWowTZ0jUmCMpjWsx
43f/LZr5Suc7EhmMw9CRLxjmQXY78+Jg1+Xv7bogT3xeqL3+hImgjBvQFOGnUsic
eYsOFKqJKa4J8pAWHESDVZdW4CoZeo9hchu8bIqZ3DcJZ1JoBmFB3y45NehzTeJt
7GS/LojwWrW4T0MUMnuwT28eJVxLtdZbewM2rIhFskii7K4m7TFTg/HofAIcFtGv
jCOmiUevwMijujpPp9j/zN7ZP0sGqc5dqS5ntceTftJVNS5crEDjbIWfIl7jfy7d
6l4M26/X60uxFepj4gaPHCJZ5mf6SuEXnQCmo0M/EQzBsyzL7/IPUsT1Gj/O4rcO
jCAyBGqojwzyAvSEJ3heW0HVEAlZCnp4PYpqoNCrm1u6evXmRgNlu9mbkVDir75w
94L8SD+L1MkM//OT1iGFw1yTcenoJzebrHt/evO1NY7EW2ZmVlUyBAApOndUScce
bU3erZJaT6n6fMJNKFXc8wBp7s8OhNyvtrAfT6owBSsvSkgAmI+C8ZZCWMkBv3B+
JbtVszEWjPyxvvcp4dafvsv9nnSgHisXpDkkrrRih7awItepOKivaRcY26pRXWLs
WZ0dZtAJIVt/RtMzwYbMCPQss5ER26dtKNSDcRqBtMDjUiSH6aJ3mnuLlCgU5peI
RuNjM34W6r3s6+cLJ+W0qGsZ5YVOWKaCu/Y2Vsg79CIdFWN6RYJzf3eF+f1zsZtB
bTnxC/vq2MB1vCvfNBPW465BOl5wufeyeKvVrUeWD55kcp9vw4Pbo0red0tgVx4G
Id3IoFl77BxpbIfEtpN2tiGpPTpy1PBbsO9ipSUhApcQ4dEdTq+ZmWskIremN/EF
Pqb1XfpT5PPzhsDxRKmWQg0UqCZnISeK/YmzO102EnIcU76NkiH2sqx+wJ8b6HuS
wPf+LeqXDIN78N63j9Pf19A8EqZNYUGRVw2+bfLH9YvXJ4ssrKFaWNcJlHZ4BTiI
6KdcN9BVzQc7rsdYkp/GDBtMc8dvWKO346SFIr3fPCOXlkCu1+ZsE2WfWhx4auY/
tk33svK3CuSlZ+B2Jz7nMJx8dxMR8m/lZSyEPTUolzgB4zz6e2CsznNvk2qwK+mu
3n4LfyY9t802HGXQwq0uT2azzQ7a633/SitkQ+42E0bk+5u0DQHKsTX50F12G/rX
j/dhuxzfXVNTN5kfJLQEL9ouasl5/rXZBXzdxRw6njVAjGTenILQ3oD9YTXuMaai
vXfQxQuSk+qKhph2QEYBDkgaHDRW/W1LHDHPBax3v/aPiMFsfvWQtNVuoRRhY6vv
7BM3tpyFGYksqE0O+AbBQDmpDnN4myJMS+4Jba8edHfy84shCzPGK1OzUzFv2S1e
3DyzqP/syFIiyCjGwrcwGJM2ZQKgtFR9FsAkXeeymyCjzZ3BYmpb4H0uLlP8aN6F
/ctslQIlDd9/bYtsEQS0AeyN5SGl8QAZiOfxl/Jl7l5vUSMPc4jjpu6j2ecemg1F
H6602EudmB6iOVyzLykGvBZLyJdCSA6o3eR2DLNfAVWll9Zz31WyoTZwIroW0Gqg
4NNVloAFOdN8RUrWANN1DkVRY+R1mQtO8wVQkPn7hkROEDxG4x2cXvM2IO3IMhHb
BImrQQnUKjJG6isn5aELdYiQZ9z0Xi+MK9DMu7caC3ShabenAlSRAPLGzLf+D8VO
fylL4Old1QTGnt7444hzvgym66brAbOWQ/IY/hAkiDBQSZN5mtyfQvFxHPi96Eb7
OvlDald/T4dHS8FUVwYpIRcNecMsQ3CZJqVRWNx/ZXjKQa5aL57DkGiCKpjOa+Ke
Pk4+ZDNXpWVJyuIZI1ML2PedQJxJa/gXqHZB69wkL63ZwRJu/aLCQ/KZpjdWn0AD
VcKOAZx9QpALdhigWYNi78auMnS3/P2ULxmXgrrlHu3BbmezIBqDmeGP0qH8gT2b
DIR7Mb+PcVgYKyx2S68qpmYvgDZ4lx+T6n4vDPr+fQB7rStyPZFEtJ5VBBoYqv7V
AwA+8vWujiTM0njOMKbPO8F1l9pghvGjC9nlbtYYVyX67n465CZ9a25OFFQGBB9+
lO1iHjEMskM5Chx3v+ouh7x+eZ7nEaNHNR109xJBFc5CFGtm/oRkLomw+ntz5VVH
aX8BarMsI+jnRf2WNeVmgAJW0eBgGnvYBZKDAHroz5Qk2/0fHhjPwug03Mg6l8Iu
Y1gKRuNFYGpc5IUA+g7FOlj1Jx3ce5S6HnLCbfh5vsbUfJ6Co5vQdwU1+HBEYHxB
rEH/bHEhMzR8g2sPyp/Db/3TaO0vtlqs7d68daXWqr9Cj+WzBLKt4yqHefmXp3O5
QIWH0WyiPFI1ba/nSkweRMJIyr7SAnInNZEV2ul9jcW5IT2GdWg+nfRbtJdD1nUb
uHpMyb69EtBe7KtVsbchD3plooX/4ueiqVeYipG9ovB5L/DvbOqXemtALZuydcTz
WYFZrumaZPFM0iE8EedRWSN4YbT2u4IY1zC+sLfs8Nb/bNsKbBMXx8uPasGfqk6Q
AVEZs8d9BVJndlSDOQwAnSKh7gs34+idYQ505lXqR8Ifodm6wSpbFjz73qQnZuNk
z95hbe7Sbtp/fKkabaCG8ierJt8Q2NCR4XM5vDDs+G7hMvSlr6AX51DisbZ4xGTW
5WQHn4XefHZrWTGC5zCs8a0IQhrwfQ8Yo1qeEqc1nSJ6zb4nIaau+0BpWIFltCLk
kul7SLnQqSzg6VHwuLbtYmkMO7BlFx/4s473NQIhoU3EOAsnce1IEI6gmdZoWksE
DeTe7CVDpLQjaaEF05PtLvtbEfXOvgtVjpHUQxFtPblwGLE1O0JTCArg7Bm3VZii
sT7Ohopu8J1x0de8HpnKOwggG1kHXU9jjeUP9A5RSYB01Yn2VO6GSilltGtwLhdM
/1m5tE8uLWwb6dsyoSwgd7j1lGjgBXAg+5of6AP+Pgn+DU4NzmJQSJWbQmfHv45G
HzIm/Rnkx2MusghF72U3pDhbFoOqHMtZz2NDY2ujLteWn1vukQPBPHlxySPBEbch
/qs34qRPfy4Qq99eo42ms71TnoAJsQDb8wwc5XYo6cTbzwvQcXBqu03BAdR4G+KK
tmjX9VohVEjs0epbEY3vFkGwQru4HSrJvZxMZU0vkoBCtHK+6TAVWMjyzJ9uBXek
dS4W9WEjMIhlXPdIHEAyikyca9V3f2WaY+G8qzy2boeMfzHgeI6eF+UYNMKPvlVJ
/2XMgvJdC9zMOnXZMw2gey1ArGxzLotrSEhNMIsvePJxKJ7u09nG4rbl1RcjFuM2
Dr9hj+lpYRJZ+7p1Vw9+iQhlo8JqbOgz8egTdwbkcSXYOmy7ttJ0q3OwhOfJ4lKX
UkMwMC3GFPqsvP23wxX1TZe8fENcSu3VrZQQklcGIfKzlJKSOgvdjktXA8P/JxET
Q/FG2D/eNJO2g49jMYAksWQ3jrQozTwW35s2ARzTELPFgmcydPSxqD7Br+MZnpjj
LesfLPmEDzXvu30T/2Vpjk3nuV85qitcti9deVB46bdh/5mLmGv4yF7QaDbgzVz9
3lG1xF7TpJPlY6QTZ7P/vZKn5ECPQGuU4Z49nl0+qbmiDYmanbXzHG9x3xz21hTp
c/Bjg1nybslbv14F25v9xy0yTgql6y1OE/9BBiZel47wUmsN3ua9etpmRDpGBxHn
Tm+uqVLDMi6KuWSbj6mJU1yZXIy95cMxBJZ/yN63ipr1FkvWpLA+8hcnV46FY8zD
sVYnpm+g/bQ3SQjFijCc2tSNszRzzJrSRW99sfanutXaOLeswJPRMamDe4dwzjKz
tawLOQIbs5Ip/9BBNP/PCuSF8Hm33MajG1/JDlZ4+MOdtqeMyVkRUda8CNPT+zqa
rCvLrlQAdFCRicodYSCrjNlPKFMtWPoa84j8dS0SQd+qTsN+/lvzRYfsVOCEm3ss
H8xyDE8FJWqWx1jzdYf7V6uiNV2Jcre2Vxed9MvZkARthZDQi/qJAWtS3KusOj3Z
dk4kBFWxRK/hHFXQXyok932/1Gj8U3wPDOFLDnhmCLwKFQIiyKi6TPq6p9hvrac0
QfnKrmXvmiFEq7fIsiTlTrERDtMfF/xQphvphCUy5a3weZ62/wr9/XNy3p+ccEkx
1xSvvj60Ov3VpxWBvGKw72xwJrhhReyEg1y3wXxrcFroRtDe9j5IPfLkl+Fe2HP1
uZCEXBu6yZZV0mh5nwnynwVOU6uLKSqqwCnFjel7WCnTNYw0MC4gZPxjwAeCbybM
jxIxlN2ZxX48UOguYwGpSfCOFZM1dMVYgPZfYRsRgdRWjPKIyBOfVy+gs3l0fB2v
5NS/buS7I76j401qPnzP/nFwa2POIl4lwmRFDTnXGNoao+m3lAqwXlRq512OUwRA
wtZzOBx7refPyEsvrUsj4pWdaAPigDiKPucCsd6PPcAioAPibA+aMaCxz/2ZW6e+
cST/WF7gLFo7+QMouYsqWa1PELO1/5nYyHgfWI4PPMOx9ZgmCCVpPF7xVosuVmHR
Th9K10uQB9hRj6BeH/jMQ7nG21oK+b5BDukn6IdNZpcQLNXYzltD5xzKxKR0opAi
EyXlU1EMS4+0PV2WVnl4kCPSoSnbWp7cTr5MxtvsxymsJDPAxBE3lJ5w3n/BYgst
nKF6PrDTT76kCVk8tCA4TeVc+9F8L89L47uWk3/l9K/gkiyYOIMqiz6jIDJDsUf6
lgkIoMXrGKfCZPI1rWeSathtNOJ68/9QGeBGbn3kjV61PVc2nYMSbD6DuWU0XewO
2bZZO/lMVnwYJNhd4HpxFsIIq1IrdozSIn+KHoJzxd9A/X3TfFtEW/+igR0qKqSD
6ZjtEhG7+RJFxBryRQFJYYdvPhoSd0YkPqTTWRrsVrQtmJ7qqOsl9E3lxWknEkj4
k/Qn6ZLrSWsAV1eeL/spMRVK6m5ipwFwrEHR+2VQX9J9zJTw4OFo2PWGp4GniZRg
Gt2yL8PmJSbT20L6PvAfwnXr48wb9L51mIJc2P+4rzrksSFbamxN2NGzsIAu+Pvz
jsGexCqk1uRYZmIaOhmxpgGw9wXt8M5jU2TiLBlsYMIKbu6S3wImUXULRmXkHX1W
me6CTQ7aZ5akI1AVGzgXM8iQD83z0enFmd9MGDGARETuSL4u7yVBVFi896t/5pNu
qQr6K63MW09FIj6TTs44CIUYow/01e8iU5W2zHW/hQY8MmEYy4kG6c1fgDa76Z+j
iLN09Yi5e8Dm7EpArnaWMO07k8bm8AAgOE2dlKby9wVTkXWcLVTy5Jsg+8e83tpN
vmFGjBpXcc1l+nDNBaQ4rUIpqbJveNrobh+mvpzmNpghBMRIwVreO1HVHWg9e3+L
BaHrFvcji1bDuBu1125D03TXW/h+THnRpmUg3qELVC2WUhxI904zi06qcAnaSfgO
UoeGq+YgR3Jsw12aAqHAQQkL9IV1DivtuOHEw3CvPtKtJlG6cQdrtzXpKvXOLbD2
YH4+f+ejrvullyTVKQd7QldpxlCRXTT7cJZgGSLuva1EKSJlldn0PWgl2Uo2Cu8H
BT6dzZyQZYG/C2NHb1xFcqFhnm1q0Hg/ae+uFJoIv+1OAm3zOxGPkJSjq0krUYn8
KNtHXgGSynJhD28VTY3JBjRPdf9RJ79O9vOtUHpl3xa7uHYx3wYSUdab9sLFTI7A
4WtWu7pWl78g2K+w4G3q2xUmpFQJTuaVsfGDNRljiHJDDxBw3OzGP0bKVGtZAMuw
8n2fg0RMdjvqEE5zo0eQSp49pxD6r/DyII5X/eAWB238XhWR4dOkpaHq2hLS6PZS
9Xto79l+ZevpeEPwqE4bLVUj92R2U4d0aMGJXDTjKn3tseT2biGjM5pVc2kC1aib
/QN/XDfP/19iBsTZijNZGyeyi/P5wldzN7Usfh2BmUnVJiPDpxqHN+eoOK4GtD0P
odS+zTnzwP7pUWD7LYVy386SGmGnKSjwo8infmXrM6jeK+o6Ukh+O+ksBZpKHixv
OlmYXV4TdYvwMuOVGU6SeD1bZb0CVtl76w+agwQmiks9hXBsOtcoCgJetYUyBB6S
Ck54ueKOu7xYSp8lBlVcJmISMoMRhM9Up73ahpsJF3hkKoNC2TVG691PaR95lCF3
SYOviVPkn/xWJEaY9BEKSTSIgQL5lbUoWuSg784pUyxSn1DLllnEfE2ZHPugIel0
C8uhEcAhhahJqOvUrvZsVWn5R6Od7xWLphrat/XzETTiIine4Y7y2TfPkpl9ZxOi
KrcE5OolqsJvtdqh8oKd9giovUBrVG4V52cH1FX+VjFSzjEoevwfXwHpo8eYCkUP
8qdoSFh5qCuUF3YWTq1IzDRVEoL/paXZDfJCpQMi2Pqkmg+ZYgc2w2lyGzDl6KEk
rpKv9LH14pDa3r3W1BT8qBXe6GCXT6Yxn0m8M9Z9c2piOQjAw37DU4sTBj0aDvI+
SomyfN1E/+2qH/7x9EVyC5/pV8n3srcQJBTiTrEU15u2GEcI2ExCTrsdThhA6Xga
hVlF+cZs6HDG0Zv/hxPnyTRRcVX/H/tj6W9Go3PQD1DN/bZw7bbxmtGs5BRP+BU6
OlQ2dTySYofflNif08hGaiYxVBBEDDQMiVaKhVnPhouF+5qN3A+Mp8GMrrNT3PBa
iucIHpTRNmMy7x5jZkSnFrmb7RA6luiNwReTD5Dzu9pXr3HkX4RyA+PtfLUUJVFm
39lvFsG7Q3L/dpq1M4cTKZ7i/swSuCKUf49NqXF/JwSJP6BuUSkRZdC/bw3kaEJx
vzgkpYdLlvDER/MCbV+t9vnMN8+ugCRDy+u5jgQmsjx0gcV90oVhXLAStVKsphqi
OxWZd6XsF21s6iQveMbBThI5eWvWRFQbgZkbGBCuD5AsAP3iqMwZAH0aml+GtFoY
po9/Gd3NOI1fdfHpIIseeproizRyUWp+8LDRg1l7FoRSxqo+6l/j8VDIblniR99a
Xf1/EkFxn6+DPjHIULB0JOwWM4PAfB7pA+VA2HpFeupuQuLFJg8DggylgD2Dhox2
a2qVMwv3GmiV8yqeDhTWHs9BxNAG5Oh3GzHSLf2eqC9pZhF83+7p3DXTdiWEojJD
8ZeM/qcnOc0TnJYwSopjvHZ/TzKGg3Tn2C/a3suOsimxFyToIG/L4jnCLLDcyCU8
gRkOkU5lefdZegum8yDx27PLw/7YC8JyHHj1vlfTFB1Qrh4x7Y5/dzA6jzJOjsJv
49rQ4Zj3y3Vjl3WNXJJ487VkbOyr0K0cTxjWuSSEqXqZjATdadd+58SulF3zHU1+
dBQQZyo+bduxza+VxlfqMOKerbkHwNnCGOyJ1DkVmsaZIQIeYCY3lInNQJp/R0+U
ofnsLaQPo4CLQOOcBjqoQbiQbuJx1TCnTLel3Y32WNz/cfJZ4WvA9B3YzLxf9DkB
geDjOURE27xD9UHem8HfjX17fEgll9UAYhoH6xmB+R3hUtIW60wu9Y4ssLstwvnr
Z0BGqVI6LHU/pk1bRF4yJpOWb/1Lgi6IfdtRBCwRb5meuQ37FjTJckAhBAH81J/3
AG3IWijAOfLzsOnMn6QUsUVQX3iHAlHtW2Zemo6seMxn0hFcxR7FrY8OiTRJ9rjo
VVhxdg9PrVjSVUnfawJAvQufvm/IIlYgT4bImPNGf3Tm7h3wwQ0/U81Re3Lxr90F
QxYwqBMHKhaZ+X14PUSRqg5/3pB59yHc26q+s1VWUNBZ/zeU+uXoT7hhrfrkuN5u
snVSm6hs0YA1MROJlciiYsddSJT6Y265EDe8V4bEJn0hRrtUV0OLg5PJFNuqSQkj
Zj7Fdi8ZxBuUq85Eu250l/HgoYInxNcCgKQljA2fnL3Xahs58qqtPAHBufb/Eqh6
5FoQmNYtKvw5AbswqXK15VOxn7+rwsT0n2Yzf47F0DLxVmWxRQ3tusV9o5kgY4dt
3PPyR7BWMyd+rRU3TbApRCs/qKw+dofRdBVaK974fYPm8rS2c0R8oCW4NsJNxz26
uYrbccKg44/GluK0oXRToGRB8cHBKb1ocxiyut9CRkfXNhxJLHLABFsBlj1HdU0l
bI3duevm11SPHD4lxzVOWwyZT+pJCdOuXJJpI67Z/dTsXYR72R3rA1PSkRLvPOlW
xP5pcCUHuSdTiJ7CuPFEsZoRZOYSaNhaJikuOittjXp1lkbs11hBeT/q8cnDhc8E
xFROadIAyppA/RTY0dU4NEt/BrJzDNfxIcMD36y0zGWAjMoYGRov8PnTMqyoMqq3
KLRW+U9qajjIeqHcNlNLWT1m1bgpT9mGE6Qb0cehPrGjVM3JONPVggnDpGHo3HCB
UBlcMh/HCk2DV/5VbGwaNWbPFJd78bMst/u7OIbeK18O7bzlITBqTCkZDlbPedD/
8xnat0ECktWyXaUt6cp2YQDdKypfmZy1rKqGP8fSm+xSclmw3TUT25VOlfwykX/9
UXUrYgU/4YSu1ST4URHpUGEjgsFP8tc1NSqzfA/isUmIL3x7KAunqmVxtQcZa+vM
fBbQsgug1ahlNmdrrD28VP6gLns6p9lKh/McDWz5rbPWXEvrnqY3/YAbAebLscxF
K8G/4EOdaNDrTgNsvJvKxn+ynNVDrFvjAAHbAhcL8hpWXn511MerxqU4MKG8UB1u
da+bcS/2eExwGRWAHvM9x5065GWO6iUT+1ULP9kH0Tye6NBcVgBTTgqKuVG7DtWE
h+KECZFkoxRsReVGVBN5PrHkQbtF9Wwul5o12FK80ADkQTuNLi1JVjWtLf//Yw4F
Shx8l0fD0fvl6s2zNZ3SdyP3ve9wb5A7EYkNzia+Z6gGG8f4t2zfJyGb43FRUadZ
gj6JlvnHtbZj1u5VV2G0MK99890vcGae8keRJ3pzmjdNJvlUpYm0IRMBXs3vxn4a
PTRVE39XhxNN1MxKR68g+RhfSfc1//hPco2B4M2tc2/wECkEUr874+1ZhTo8CBTx
l3/GrVD6Xr5ATVHJ4ggHe/LsJCt2kvN0XGLId4Wn3U14wVxjlmY0Juy1hPnP68Kc
U6X8QF90YpqM/uYWNe4b/iz5PPwy+p/meDv5E6TWHl8mvPvLbexKy/hC2DKbgz85
e5fabUVUSKrT8d/BmDWgGBUrNSx3moJw7ekOfFJgh1OSEizjC1dUkYCzx6RNwTIQ
t1RqWZOIAQzEL2jCmVMD3rkwYLX866hgmfonNj9kJbU6yx33k4j66UEf0zBLZxEG
GnZJrTah9HioDdzKUro/NpTLhnimal0Kv+STG8/kEQ6w2w8uUVzkEqU+ODswckqP
y/dpJ9YXjpUTuX/TeskgW5+XbqFVMbVttpyceh8GSqVPot8dSAFRrzZAkgR29TdX
0twOJhGDciPeh+DvvuAWXPSh9uIYrxSATl6nFOgZKL0a2APhDlri1J3B1j4DONYo
HuITFek6E8QUcrJZbBDrTUCMNeccahYoqALaIOK/ZMa5TcBnOrRP2ll/d04Lg35A
D4mU5Spmj1ZDsCor10kKBey6wnH6bDeysVY/b6jNJh7c6N9LSEqEOnXOeWOnZ0FM
JAiENeYpDnntrWci5aNsmmTX/nQmL3O5FdGp+LFybYWxuycLROInRh6uUjR4P+pE
95wvSdK9AMgvzagrtS0gXOUHWQ0DDcR46sNAuRB1l1XUEhk1N+AUqgS45KOMWuo+
B+UKUU0pHos6/558JPug8gZfdj6Fw1ffe26b3Fbrd/jTYznz3K808ZiTTZ43UxTF
0gfXYuXp0h8CYjB7Wr4JlkcNzoV9R53b8t34bSWVTM/0wh8rOTFbkQnRvB+3xptn
Ncmjj2wma3Di7LwjVhWVXppv07njDSikPgq+iMIiFgwC+ebIiuRK1pQyhQ+iGWWs
Px0Oy5awZaqRwwObde9CLHwfmviHRyCcpoDiyLDe5bpA6sBrsg2YaKr/sOXHYyJy
X8f9SYATVynBs4x5pfH3g5Du0HLX7K/tFGHJSrtcxQoIqAPJ/mASYiEdGb4EagyF
53fmD3iv0IkG8pZVx/SPXwpcZzrS4agiCdR99nF1q786XMW7CDMDpED+vOneYgfg
5NrJ8rCju04XBahZFe1TokMjcpb5C/p3avlN09fah7r4Zu/yCxKsLjCiyzCXSwFl
jj9aIp/JDVzi0NjGK1qtmfXKMCzs6T7hkh2W5vkN3N+cKg2rocuP5DPFyVq/LWeS
gnQsgjH7SXWdH7UctUHLaOmy1Zv7MbVSNSgJaa+e2P6vdxL6Szv3qtWFkOjubHZo
9QB95r0fIo4T/r103YA+yQTadsXtxTlDVWcCcn7rLRdqNDD3QFPPzzOea1WhvjfN
8oc/ntaEcauYNEvW7JF8aFO2a4pWD51IF4+2caisOwT6ycmMeKMJJMK/RfuMbrZE
WgITAdRWv+PUZ1o2ynkBRveNMgKOS+wE41VHbLtfvTDEBzFZO0sy6WK8MVTdJMRJ
VAdxnLmyMW3+wXWmEMiHlTZVyiyTXNPbQmRdc+wdVK7ZUCjP0dbw5rjEgl0PpUlS
sKu8zgnRqPz+9QuJB5bRYQbX3hNYiQAO6Q0Dp88HMpHUKuCOhAa/cZB1bebIQwCk
wN8+/rifnsg0BhMUwntY+gk6kRopPI39aUxKfWXsMBx8tXp6SrPdJk9Cs25bulcd
fyuo+9LjSOrNI1OZob2h3kJ+4jRZk2uOg2Lot7K6yS8mmXoN35bbsP5b6QMs5Unt
4mf/HfWkEh4IZzczHA8cuCsRscyZGEOSjuRGUUuC9XA0xrBOjY8sIZ1Ji4WYCCga
6kz3KnEI8PWmrBWRJNSVNemcl9TToO8AfhD+3rSlSjQyW0J31jZN/yDVGNATfKB8
Zn/reaRUwQrdPckHuPiQPzN0dH9Iv7kTn1nL4Y1Y5Q9JiEH2PFrOeyMc05I6HPx1
29w10mHDPTbPvL0xEyXl4JBskmn/gSqROXqxQhMUPs4U2bo0XAHRRFHmywwJ/+cs
AHjbZ+eE+fA+cC/xBwtAouwcTDp1kft+LpLzSDvpCszeX4/kh7gSNrbnEHri73wZ
mYobLG/+qm+s//QBUHLo7wSM3eYJUk1P11UvKYPsyU3s2OUKCyvRjTgP6eGL4HuC
7KvRu4sbFCKf32AP1TujxLqtck06K+3RwP87rsiENs6eSP7YFhruxwLQqsegJlCo
ONNYH6wR5Bi40ZPed6INE1ysllfL9gQikOaUggNONwPIA3JGSZjde42XRgZEaHWT
e2k5WMabtNcWxWycAvz4MwqNBtgKON2evPr53aivMWaWe827Us48LMgFuhsCygeW
sBqInvwET464poON8Oq1Nz2uOHrRoqjfZcN2ejEL5gA1N+bRffFdbzTySul9Xb9q
upcahRSVmITsYcPmUM1BtcAujlBMvpcvikyYp08L5jZ37r6PaAm1r8NGfIK6m/0v
44mQpZHQwiL+dOIRhg4/UjhxVE9tRthsn1tIb7oqIy8BWrJdRU/g/h2WKP9UM9NO
pzuxIMQdf/63TGUCOsVLAPxFqF7E5fhKdkReWD+yqArQhMRjt40BbAfY04JhxaCo
maH5Iz04yDqKZzP1RJY8jdscuv50ycOj1M5QBJiWXNXSansfbQAlii9dAHV8f6Bi
r2LzjUJ2CsTqRx1VVm6CM5meT8N326tmlDmKTAZ4bO4Sy0HvbV511NC5a4x6HUXt
YUaL2TRJW6alk6IBXwJdjZ7UtAJFohiZOmGc3L/MIH6Riqlcsk4YxvqsbVPcpz9j
QpQK4hufPcfW7ymSnoB1aY1ahNQvPU5C+F5UDDduAFVVTtnFt41gTTMS2nCuxhzo
G4rGJr60HFDmzNGvvalVeFhvk9mSA4w+lgYAk+QOgx3bhGqfmm/Lr79Acb9coCuM
77XKynI/QUpr+klBWvZBMPaTTAtgADRL0RVbyE2Kkgm7SuNoxYAXTbvHE9m/fXaW
QY7TLpnlbk5rRsd2e9UHStfkm9gFczy3guUmvyiqMnd4fQAR0HvMn8D6ALEL0MtB
G68I/X8rsYtjrvz0em6MeX+CLtEJhF54DAU4G4xGyfHJfIoc7x1eWB1pa/CpUFRQ
YlRYHDMwPXMi5Y4yGy4FTG7BcE+/oUqBzCPW+TwZzGTA1bir1gIvJIkDoslZCAf6
XgGREXgm6BpLpMrblXOpXFUcaTFnwOyuT5A7nK+4doSsm4OpQCruRdijwQzGCypA
H4SijBKIbl3xxeJwHknHlPJlSTjV3GHrC5Iqqp2eAanrQzmX80QEATUC+9a/BtBr
ZWeCPAhpinjgWJ+ORNhsw+M4xKlN5Ocbx98f0wX5vsW/dXzfaMC2VEXrwIXOZLXH
5mYSlRLQaQSpC30S+Gy/Eco4xf/fRdSj3NpJuFL1O0pKJ+T5HePliVo2XsSl+of/
DdCQUymOaQKqHlYDp8pqGrFbV4A4VVdoEN/6CyxvVnVWtKnYjRUL8/z0JDP1R/El
rjoTBxZEtI8WQA5/ezYdmTaLW3WZqnTmKtSLIX36ccvWsQfTI4OCv6JLntJpQy9f
nMMXA27/BtZPRXVEBUr49+qh8Sqy5CKYpMfTm8MLhyWuv/ZDVBHzSkQmo10upWh8
mOyUZhdOGSg4xO2fyEZLDxFCKrcGJM5v4vzHU9ejGdxc42UuSgowpoD/HCsgzsyt
WsieWR0CFzsvZqFZd7HjKHhYk568GyycunNCV5bR2m2yTPAoI3BAK9xId34TdUSe
3SLuHLCogvurGSqgndaAn/ZKY9HjtlH+jIiVLfgc6g2202ntCVr4Rka4Fw94DSjx
l3Q9zeF0+Vcig7Ys0c8EWK06I9srMaSwqY4MMYyhkXGnvET3aGULQsqXP2cs5x4M
Xjd5/O/ETrYddAZQQ8BdHXhJVkPB2YlxUXAQUT1QDRUjBl0XyFKbCxujr1xhF+ds
G9KoGkcgtErvnXFX42CexcIhIDA27QO+dj24Bmot4Ti2nl4MVz1A4AHlF/dymeIr
Jr6/PboRPcXGy0jCt4WdEFFidtFfUEMjW0PD1V49IMm+77n8o+sk9XpqUxtr+zL2
Ca+LjC3/Fhf2uiCm8gvrpXYFqel3HCYcKIrjC0xU16gxoe97zq3P2jwKm9MamWOp
Lu9SyKOyc6f/+upC5IIdw7huRENtSQNTp2ps+6iYK4U2PK2PV/vmJtsiwbcRs5vU
n3t+WIqenmcgj7gCdMinKwzK5k1PCWcmCKHRmHK7lPVFgqJCbQAEGktwbw7upoWP
/udFUwyM3C53VC8+mPsmieb1zOg6tvTlRjN7dOiOWjt/AY0ZBtacD/29ianjLEGx
2BPMH1LQb0zIBEc2Z6BxF3ihS7tjFjXQSokJ3I47xADeoF5bVxUEHp90/VBvtL8v
HOlMgvd/qBfsjaSOX6IOuBHpz04HQOuuJ4YBR5B7ndwtGisGXh2U6VfE3LbqKDJT
vioJtuslIbAwcWvFg8x8DStMIwsErDray+sM5J/Bh0mydAqSyEFOOVhV+SM+3pRw
3IdUjkfqlL/fCxo3cpedAdyzbwRy044s98OjNa42bM45Dd+itw/ZlIevJp45aAlm
kRAruEdP27BVPt01i86xD7aTYs1nLXkZzhRycQqPLMnzpP1z/GtNFkNLRf3O+Zdg
/oXJwjcutcuIKyCkmKgHnJdEIRSoijHHH5x5wsnZrxaVVHIE+SxFGw6NEWBndKxG
TsgMaZCCgyYXn33P43MFQ7z+XAmoOpWrFh2EfOIlHRaEwqDH6VgsL2wpZaUovR22
iTyg3ggzgaCxara6ojCIjuqJTLG4f+zitoKs6WmhoKczqpzQUaxiRqhQUlCe0nQp
PJxA1RquSgmVmmqvoJyIVlLfWMUDaS64f25xPJ/jgz3s9fKuheX+644F30+Y36Ed
N9R4DB5U8r2zVScDYm3/ew9r3VhX4We8ISw6gw8GWTjYtjygfqq94wnIaFPUxTH1
+lJXNetzBf9n1yT0r45vQEmiNrdH4HERcd9JKziS0m0Rs/jAR6rdNIN4K8Khu/lw
zUxzO3angfIfFxvnuw8A59IoJetRE9AtOUF1DOqQTnj6mlnRCKXQn9OCRGTFxB2s
8CTPxkSh9e7Dom//g3J0O1Xv3aaXUBRVQbfAxtB2UxLrRg0RneL5Mwm3Y78d4thC
F9A2aLFOrPjc2cfwM/veaW6rPJEx/qJ2kOJyuxoxexYxtADDS+Z8+a2w7GH1FkDU
uGIC9zaBq5KRv8RCodEcCGxEXx0ai7CRR1y+3vGC+W1uI/8gY4FLGALpiDxwXJkx
ZnMVgjxB3C9/g3kHYkYTt0eVy214cx2ZWlTczGuVVyCwpSQzC/jcvThc94wq81Aa
zmohPjj5WAOf3tik1SPluWCoftJbgRudaZRSWRDUNfsI+bVc5bj6b2rFq4hyHjkv
c6rBzUENMoc0+LWKojyrZsBQ9ZBgWowI4WyrkhmOU0nCVBk9yveZBkgGlHoTdSPw
11f8DWn1A2KhGqODhVU7w0UBKcjycABasbkxxBZ3TkDFc99T39tu4h5GGG7PpwjY
g9mLOJaPXSKi9Qdx1sCK58MJNXxP43XzJbdmYofZ5xgqUJTr9PWcGxInlJ2PmrWw
3UWD5+AnTiHV8ZNA9N+b72RcaZxMxW5qPDoTvZoCEUSZ9PoOPScVfM9FXpTcU5bR
2nLoTDY3SOjtJ8h/EbO3jLtMlugEkQVPY526HGacOzBPap8KV+C+3eFTG6ii1xEv
2qxy53y3V+QRCnu13oaaxWK8k+pbuW2OH7ToL3TmpPTBA5XCQyXtbQf7RDYtqH3p
mjTjiQ97N6G70qNYO2m9Wb2G/fnA5Zc2zpJWI0NtfEa7Q67wQ3eVA3qrREpdW3Tx
Ll09CAMFkhIs2dAprBhSV5NXVqrfQCaTkXQdlf+RX+S9/LC4Eld7fjfs4qD2Ycub
cmLduTMkntsz3mglUYBqMFwHMNuATsbaW82fZjZrnVH2rVaQRtTiDeoVIxv7P7KK
A2MKKrN2ri2HiwGNEExHJiUiwpg1820r9JzoWrYIuimKhSL/B9qerzvWuUy4HNk4
43RUsrrZJpvRvFDE8KZSNBuTr08HXCRQhDzcm5jFRZpNYxmLrayKBbYKb+iRpHXq
GGhpMXcn9j9uOdIkDVKE1XHjtjSFnYj4s38fjNX3sj5NhuyHNlbrLYoBLSEl4PJp
RndCXf0ooy8rsDuAtsBDWA46sEE5mWWiYipqXt4ftpTlnnFIYRbL4Ehm6Rq2ssW5
boRT/7fjDiEn4VLSbpCjv1+nOfbrOmE7Gulgu83gbJdgy+/gr8QGry000mkZBCc4
OPc6CW/1qsVeOTc7wCqxmBYCaWv97twt+EUcRjl7ouoxtu+vY8GbmdkwDoWjxcqy
fYPas0Fgk4j3ikTLgMR2R18gwemHDqQY98Cbv4LxsZOaFr9ozHsHrjseaOovTdPs
v/c91hn9jgYHf+wMiuKi5A8bRQ5qHVIpaPY6a3jojqexEIuY9Lde1Op4fNP1qD/t
wObM7BQrJKV4vgZekvWmq7iI9WvZANv/5D07nWhnzfHe82tOIifwyeb61e1GdfrF
kHFfbP4/HQ4Gp7fSDC52w3gCHzkicLYehOWK39xl1hUt9v/oUgb7RS5YRTFbe+jM
QdlydTuGXIFPiVL3DlG0dbMjDVmrVosxAq/VRXFh9zeB0zikOJCNZVKecGxF/ARi
j/wwm9jCqkH8xwEWeHV6RJAnb0J2rAN7bgpWrI7oUEcr4EIrC93sXz37sw6WQPXX
UIYKEd0g56G8OSwPXq8SLEgJhHkf/iC84fZGz1Hs9+QZymjyCSC0TRnTaqN17bLV
VAC3SLMhA7r1LMOfmzF7zg/+pOO4dDASDkmGKHM5ZueLukyGcOICUlK7xR6Scf+0
CHpVL1kFTQ8ieboBUn27dc4Ku/q9oibFKxULNHK0r6dmOAUW9yzkueQzKyBL1sIF
iTjzSr+m0iRnZV/C8I7kf+2H1CbrSCKpR+tfF/3fvSCk//2UQvr1ObFdnHBLe5sk
47UuQ5n+qZnohv5Mml1WlIfTZTa1N8Rnl1NyIN593ElL2mZxfZ5wT4ga1kLLeOmT
BiFK+j72wcgMawAuav9rqEI4bqOL2nY89CwAxytyD5/5wivqdSyBD9ShVa5b0N0f
+oJezAuK/ErFs1GVQvekFsHS0BbM3PpBGOYLLv36aA6RzLjCuTlNY2KczT9Sgbo7
KvkG8gGEycyjbkfmYRMYjPJV8Um9yTOnmPWCsZfPyRf1odnYfOFjNZ7CxGxJvHzx
2sbjqpv8wiH1Rf4WZPC3kUS9NC5XP3CHH57V9MeHWgzf1g4d131fXYzMbsuO7S5u
e4ODHV2iSG+CGisXivHKpN01PvV5XPfu62Gkh2nL1iFyCVo37KhJdTdpgHBCvMno
9OUjex1ZyB0A07FNVwP9s9AVHU2I+tmO5z2zwJvYlHaKrwi+4fFefOuxng9xIiHC
qzwIqLG4/jjZkFPSmFbdL0PRD9nmlKUWnCh86tn76nAGeDRdU3HMq/0b9aA7ZO+7
nOdx9l9Lo2VHLyItG+Wbwl6L9ccXOVkXFre8HXbTxfGTqSf1mnNsvwn27LldMVus
y2NfJezRKsoZ/m6uxVTo1tIdeFlpk/XbvZEkiVrAmPffSDQqhLgAPme+Xe/vNe4X
EL527WfL7AGxwX2YKsGkgAzYJmxaNE3wZTHQIktKtaaMNc8wMfAIOmwhSFYOL76/
5EOQ7EdJMUoMJpWyAnZa57R1P46xMKhy4B+cey5oPFGDay21ZBnqc6JAQABX2fFd
R00T6bEZ6UwrzT8aaCaW34sHrVGpdIfiruZx/tlnLVFGdG96zzyfuXV+vz3QG7Tr
KW6nnhCjIxwgbY+Ejm13dsN1Ew3ytA7QIbIwwDHckUUou16T9cbmwS4hM7IOmPgc
y2WJOf/p54xHAdjyh1vgS8cncjzaFNrIDJQRZ1/dTa9z1szEl9LrTStRhK925N5E
JyBwo5l3Hc4HXAA4dT7RoKTIydvL40TdCYn7HQPMfuCW0KW1F+CxkAnsmyQw05Ni
5TolJ8NLLfAghKNQLYEGfD5+si60mWbkbkTabCEkBUVlss/E142+NdhXghgg26ny
smjn/fwxwZEsPg3GDRlGL0YRwcwU9o7fwa5XmZ7i6os6UFGNxOvF5pSiezgRcswf
T+b+AX3opbRyu/Pq1UwSbhd5YuV8r2mImNM9Nb6AWaktvDygKPcCbHpHFNICjK5G
Cislj1ljAYblQiKfOjSQSkawm9qKYAweKYQF+TUA14nC+piVY0MK5wwMJI9yuTJJ
HU9AkcQDegZV2R8MkFT0NCxyqkUh3gctHuEDN34lMaMyYu6EZ/TeaOqV5kNY1Yv8
Hi0U7NWa5jD6iFUyYJpk06lbd41C9F1WmIrm4dIMBtyP83JCoB3UfhbaOgmW3xoT
h79LKJK6tlOfJtt1qUix+n+HSmYTThk7v1zDulWwHZqp4SRDQVU6TAnlH2okV4uU
UGWacEF91XpQX1vpBGN0AmsnDtNAjWGfwG6krrcYpfKacF/yhPzmRcdk3jMFqMIV
j/ytEqASCuYN0yCnbWWOULxue3ScpXbiBg5lFAxh7UFOocij8ScEcnP9yVS8Bnqa
ZRJu39DLC3Zvo5l0+66Q/tQXa4VkLgRotlDxhqpAVcEasqjbr09qlGIIV4X2c4aJ
/K/+WwUDf3JTIfadOrQXEIuGscdudXLcNT5iBGYeIBNZe3acbFCGSLFCIacAmHB0
0en93iDvGa9MeTYpSIzgLgGJGELD1Q3dVLuS4eeIve//KQNKFFFcxG9DwMhwabC9
drvJ9/UOeIiH9tsUL2p0Qs9dfS4HE6SPcXrk74LusPQFtofwKX3CImwI+BQWR/uz
MqF6EYCieVdF82T8QtU1FDE/GRRd8BVeRj4gIO0+2NASnjqBkXP5Pakw7DWXBv/5
wWFYcJDp8lJ7sGL65t0q1Cj01shmrzMHiEs0MZw6WBoSMo7zJnnxcjOIbJczS4TP
Dtp6NE1nhyxwNziiOeg3FqnZmSJpaZOXaM+hYtnFfAbtYHU+JYnNTROJwg5s4Fno
nB2rxw2p2z+3LVzYGftd427Wbs1Yj+ljhYS/lm1yw5GZjSK9Id9gDn4HvyVeDEty
LOmNGPKrc2AmcNb3/OLErM4uYuv6MbtE7Ft5/8SLWI6dBaKTt10xqu+tCmaiNn+3
RNo9KUMCtF8JZU0+/TiEIKihy/S/mBBhhAUcDZLBJNGd7+6jdsIKtjtZ1xtS8rzc
Z0GRDwGUPoZ7CUXoZYi5Ph+ihwdoPEp0ZXg0Z2pgaNYTmygqRwcIPzMT6ynb//e5
sfZt5eUEo9peLf/JhcumBT7n7lR7QdepJvfhy2FKIfzctiosUfZAKVATJ64CkSYZ
UIABHJ2MB2CV48G7Ig9RrYYMyrIvGea+sM+Xf7XVVM8Jipo8rgig+2+DCnM5/s3Q
GrQB6Azuo3UVnhyAkHTM8q2QTu+CLlFk6Wr2ahjU8wIJtt1601M293CG1s0JSyed
I63yjxCkZHUV/waloJNiQsegDLK99hBl2Nhn0lB15g6Ev0BlLzQYcBEEGi1ypbrf
RD/gDm5PETGdE8bdV/MpnMgQY+7gwtjm/FoaTchkLqQddnqEyulV5PNNf6xVDeNv
gjH5f2H4yWOPg2Rusc2DBc5D/MXuWkaPsrJKvRkSyV2Ph/LhVCrFRuncB77X7TLQ
GdPu5zim3rixAulcYWNEeH5z2+cKwdU94SckaD3tym0Lc3Y6mpw2uD1ANaFqAIoI
rINYEGRMYnCjYBCgnxSikYc49JTU72iCfdiOYoDDuT8gPphxnYs9Sga+yWYBOZeu
dcPxlDbHpoKB6PU3N5zRl6wOzdmYZfmH/HxmPRFgUyNIY4UhhIRV0ur4mT+Aj48p
n6qdBNSnm4Pj01N5JSOsUkNak1r9SpU8Sl5L0o1nF3w5IlD+UpDNMTsU94XJGBMs
aLAqn2bZWLrbfZ7x99Do6syHanMuG/wRPky+GuN0Ve/vbPN/fdyMhTkT1c0kX2+M
OdDeq2vTYHi8m1aDTijmVp4yEV79u/u0K69ZrClGxkcYXCCKFgfMvvEMfeMOZEHT
kNjJZRJp/vkLNkc2xjCRml2DChwII4f6tBi7Tmrrij9c5rsrdlS6lO1OXKyRw0tO
VRPsU2i9VDCG83MtEsgTw5FnaE3h3bPeVOOaHBOPHgLS3L5Nsymp8WWLsVtdrgst
+WLWkm90brS07yUuVOz2u+QbDk2M13TGQ8awJrQrmN0OeTLI4qqiQaIWrzDyV4Mp
bmvio4YNHPfCpY2WNmeb2163/pXNszbdUcyJIssQRHLSEYVBwKE1H3rbH0rGzQqV
vo/Oysikk8HWaaby06f7TWXvAqKOPiLnUjQGrszzGrCPHK1yfnR1KvkNAlniWTEU
ucVFW/zrnAqMg0/oUI+LRCfCZqTRd1IQHJF2kbb7Ua8PRNrtKfsl8r47rwoWS4ol
sjc+sERrhfIsMt4/9mJAPwtpPUwiSghjI3hAp1REGi39U94Ff2R6Zm5dsfDcbN/w
pEDE30WjEzA6BVluAtPyn6glMw/jTSj2xuvuxpeYO389I+GdC6ko7N8oQ/EBMory
5tt3UibCZqkV0F69Hu9Shzq5vTWfx4FiAFec7rgfDokR1xVl3A0TPmJDmD5/N5vx
nPj2djntlG2q6/R5aZiaYo8Aw7jEJs3BqriFX1dFy9as/XyH2U47ee7lcoOx8ToK
VfNZSA9MhT/kwq8YFcDBvBxy2goC6PtRzCDQuLA1SgWDYzniqfkgHLA1NT7R/e+d
8Wdvmcy8hD2clC7NxF91ljyr9Vz47zSdeOpLcbr6648tB0xPjwTXE7D3chn38nCy
tCvtIm/SfBXAUjomgvxCfupZPPefsEEJdiG0O96XQxfEEOwDUjgnpE0fIdC8uFb0
rYqo2/NWlR+Mg5KO0R/Kr7KGWZYnCHPKqZtC7KB+JF4LyDLyFz4oRlE1DGsgiooW
5ufivU9OLSZMHTvvZtUrjWMgcp27EN35bbMPrazUquhMv3WAspZrfhH+DHAo2XgI
JXtfg8yVkM6Xp+Ywzkh1/+1Pnti8h/oZ5JvJOMEh9O6FIhTW0TLjIH8/3Qrjf3k2
OpS59tyZXH3zHTpOMTtD1nY2X5AUEfjqP3IWvT0WzBmr0Opjls+MkLW74eUYuWdS
1I3fyEvqDPwYXOK5JFVPNvPYjH+riXmWC/QpjaXGJUqNBdhkMedr2vs3DsHhOiXR
jsXCi9HR2G0kKuSTmQNn62KeOWoKbfsdPWobuHic4FKep99wcS2mAbJn9k4D/XVJ
cxq2pn1Z3y7uFnsRN4kM+iQ4Ih8KA1WVXQnSSGSq/oRON2zUEfv0UQXiLoBT9L18
2yLzjjYSk9+2FBBsa20RHJ+NDKAxsfYRUgUiJCcRbQH5VM7UrZz5cpPrKfEhiOkp
GGvWoDtnlYu0+1LA1FCBJpjo2PxiKsePsDC+HPk+9x+0E5Vbj0ioXmNuptviQFIE
grpa8ahII3KoL8HO9Ic7zuDgMIj7KiOcGE+wblA9bgCNEWPFeZlxGrV/Uc80PRMS
5K8E42TrCYRbnM3AXiVO2e2vh4lnwSU59qHz86Vdj2PskET8YyVuTb6nn/ulu2+c
/+nbX7xE5GRgWBvwewS14WlY89YwuAKdx/JnH8wO/HBprcfC3a5cBAaoFH2oukJO
4h2+tn/GljBhzrkmlawgPCF230VsTLfhBRlLn5+aX1VW8r+Ly36z7DlXu2HyernL
S/ohWC2H49bJs80l4RVDL6oY998wL4IMsL+ERqOp/WmcbUDcYd5iQw1Jq0URxaMR
5a2rnqUEfgtJwyvRk6b3Armh5m7L9NJgyod7yiBKMFUSrXy8kxKdXO9caEjB3S4H
Tm1oB0aX6ssNPJf3HB7ad4xmSdoQTDIUMyMGkjhGmE2xURyUfsE/kVYzq0vLvAp/
Bxpj67MXf5jteLpRGrIljlIeoGoqOoLDGb2TUYP6UVf/vJJ6UYmXRPoJKkw0n9lO
kcKgY7sgB8yCGxjiObccfBt1VUAmQVA189YMY1JyBM/EOQ+wUGlHB1sRuibV6ySM
I1k884XFqOQJ/WVMsWMZuFh/n5Piphm5cIqJE2zjfqJqp/3pQ86LLat9mrVxMST+
jTiXi+Q73jcuCzAQPEzjZksSRNLvpyWvwSyp6VBs5zDAq3N3rdPY4EZmMI/RGNSM
NHN34TvN9BFIRV4kybh2WLfi/erHaj7P6Fh6zeAbYxj44pL/b1Lt/fUoOF7lemVk
c1eB7w2hnE1mzkF2DJtwEc81octkZSOutOM4wkMlIaeVrOcH0hR0mWIVM3bhKH+S
WLOoObIHgUijpbHikk9aFMG9Ng94Kde6MZ+1Xs6JhtwP+Dx4YNq2pK5GQFtR47vt
6PvJScBIfwOp4lgA21HI2+OWAEQDU+C8uOzitedvy3zoANAKtTvK5ggRuFem2XSp
s9R5VsIVhZSh77ZyhJS9uBciEtmaI2P9HszQadVJaxlShJf1P0TXvxSp+UCx4cwT
muA/imMAXdaVsZgj1/Mj2wgNbmWeYRGxTxf11m85ejXjfrkl3bn4iEmMGTfywDt5
2qBsZW4GB7fHiwpcw9N5WkM4VD900f/nWR9c/Y7xqoFtWvCV6cyjbgL+FdP8ZhN9
6kr5eSP/oqciDJhpruevvbYVtJ6ze2ETNGicXm28qaVEgXcgbrppdq0v7QQsyeHx
WsKnicaDtWXfHYkAcSkzhjNZMkKsqcTmXdDKTZmXFxLe+/Q7aZN0CjYWDMxxYDg+
3eAKNo7uxbWtGq6NRUOwiLf0MUK29wo77cULxVqP1SAbuUXs+QzsP/6qRMevxD+1
ZbjNAGhQ4pZb/LE0A7kMTdn38Rt4o7HkvV8EFSXpq8NFjX6iHETnXNfyglwENJ8K
LR2ZhPecb0UG0BGRLU9+6v7XWPfxVE8dMaXzBLl4I7ARrSH/dtNzozRrV+UbeX/5
xR95QEDSdU05liEMd7uB/2HMPD4WlYV1uSkKnzDj+30Ixs41kdqfjDzhW5Fubqp/
+PLvjbKyKVjmPl4BBp2QtRq/RibOlT4jQRph8hUMW1nYhqd9wfaPJmanzlDnlW5K
mZbGPfj+uVXF5m3Muq7TUps+00o+DG+i6bjDAeBR0ecrrkmEaUuBGsvslkYmJi2r
6eJmn1LjCNMU5Feu9QQY3UyH9eg+FnUq+PahXLly6FWS81/Chzy6/SSlg12LOu/G
OYUH708NwYKBdHSwXoHZ9BPVvD1MwoUk2pkkaAyCYNI55s+JRh2WAh11F1phNxVM
kS3gqRrj+oxhXEs4Ikb8uGnIq4dJ2bwB6QJ8mce1kfrZ9m4GwfldvRzs6/y1yYnM
ek36gLSthDsZCm6LK1VKGOSllz+Z4cB1PJV/FTg1T5t096eYWOPmd9YZp9bkFslo
ILDKm2tQCWmu78BAAYeU9vs1ypTU22d2rf6cgXJ35lJvwq9x0MrTzf17GPSQ8hks
ynWMhWqPx7dxRbDk6ZxgETrqTKz/Qz09lVWdAfYFKW+DfbDmJB5VlUKyvcSzL2t7
4UH3zMnq6r7MdwFsb+g8adzP6CrdOizaRrQ5np3y1UHG1VgnplaqmY3A5u1JugzX
SlcEKQ5+ouplYtzKb4aTNm2G5pHRnzZ6OZ/pDOfBQ6AdFhKEg3BuMMySs96o7gt4
oasIGK0G8ykeDJ58uffkd0X7SBcYu0ShXbNyi01VC3eRd12wZFxFJdgzL/wzUBiJ
SSUasLpDuSQVJkYWTkuishrdWuDPqhD8+QGTuxEJvKHAjrrvufZk7F4Skg23Cevk
Jjy/VG3EUsGiI07GQErMIcQEBb0CwTB2KRrWvmEHEKxiFF+6DD8GcxkiuhxiCqem
Ei/O0j+0Byya9Rzv+Za2Yjs9Yre3wYeh45yPTi29hf7jcbHBwaHBj0/olZhmOz3M
sKCaSLNTRjMfaeiaKAcVPlleqo2TLdSjpLsEJ2Qlxvi5bYpKXr2xk0njOUrZVYv+
9XopeQVKODLh3Qo5IkfGIcKj4ne+ACz4e17d4alkKA2l/axlVySo91PlpxX5ZTjg
awMpU3WUVI+0nspDwyJqe3Rj7hzRQDMDMhjwQ29Kj0BVmYHmRa4K9hDXT6oeJWch
ykGN9o9pxvN1Jl4xgLrWU/XAt66TpFUxSI0wpR5UAjqETyd+7UTzd79BdprfNiDd
eCWcl6nNdeLV4a4secySKEq2e7V2fvl2RWtZ+whR3FLOexk/rjgeRQpb1GmMzT2m
8sJlg2lLIp6dkjPDZ/S3mn6ZkXX1A6IPW/2PlJNXnfv5xU24USxQPWXeSJFoRe6e
54LQqxriUUOwuBUmao2LpYef8CqSoXfKmxtuLkouuXKIpnE6wQvv3OMz5fDFNhJs
DehpUhwGfrR/xNrD6c75SWqoYqgJOut3uEssZ5daeZxjejyMjcKPAPb8muOxMKtB
0bjK7kp/p3b6Mg1WUGyaexDFsMA8d7INIX/mcqEMUxHZD8nMP9ilg8hs8NbiGNq6
NaPGb7VApR0EsBKZpvOJbMoSxr0/IzCVFXajo86IDEqRtgS8bR/1yD/o1AZ+P0OS
WnmYe+xM9GvosEk2EYNG8SsLxUPIq0jkYr99tbtsN1KbTZypk1IWWGYvP9BLvXWe
KMMr3uqBe4P8l5LbFw59ZCHpASqmE3SJ/5+onneJV6uYFZ0K6/wH07pRQ7Ne7RsS
yh3j6Zu6kbDhYnIGqWT4UgF7Vzv8nRSCEtMiP6mU+oAM8qSghJXDG4l7yVrB1LLF
9zesHJBK4rJfvEsjJWhr/lSZ+TLWRYg5NSRCZA0JmEbds/1jbtCfYLbsGavnpH0L
Vxs+SQaCXsnQez7UOyuMq4EFl7WrS/aZKVkIcSLfLPTwv1jLHHCeipMoYiJb/W4M
0G2JYLltgY3onrqjk6ptul4TlscLiYkPupbFC/sxLBLnohP/kv99rm91q8P0KD3P
T3uh8l0ZIXPGEi2XuuQzPB+9hvhBWUNP9o2yeenz0EWDzKWoIfAICv2e0KR5xWEv
uskOyTjAVRqjpjajK9TmB6I2gE+rghYP5q4qVD2kXniUd5jVt1VbG9qYFDFwpHty
iPBLrhszcfOPuJBY7nJZ0fItbWjIIgq2QGjRSIbYFr72yai5ruXu3AGpDxqM1HeI
Ki4YbOCrzKBUU72vXsLR+ibqPYEqDLut27QLhHfWHr9hXItRYdVaii4ZpemGR/HB
pEOHReOoZj8KWKiKFPeZhvcE9Dm9jLTDQCFgYOvV7R90o6DF+hnRiN5+Qs6TghEK
OLc3r154JDkVKTin+N88tXSoNAFrWhxbWVm+cftGXNOy0TSJgA84XdxyOR9mWcYR
6lxgXRyI99OvavpGOGx0M3Uak05RsTHVLCgIzQbpjEoybBxbfUmyEF7I8ozenX04
1fcZ6WeYb031MswJRN242t44xxpDVXEE/ws8bNpEj9WByfTtCaqIaghSRMVlkNOA
XgnnSG17fh7KWKn/3depbUi/dVp0yc/c49m0voA8XblGyHNtyIPJhmgitDik1SHG
bSpTyOXtFNTEDeD6BTxHY6wH9MVPkxvCzHnDem6TjHwz6TZHA2GLXa/ektyaeHzt
dmlc96sYMFQDI713sk69xd0PN665x5P+0aXivUx+LD5drX6O8HwSl+IGU6a61Pi4
JXPdKAlROQLmXs/LgULc36HlSjgLJtYLkU4n8d79h5eE6cEXoJ69TjDH+OqIG7wU
aobgC0X1dix05Z3bdeGVidR6mN1WurwbEWG5rhXlOWWvfEzrSqVUUURx7B3dxud+
Z4MHKKM2hSwXBcggJv7IDn39DpaFONN2SmgLkFst4Bbo2Z2UHezWm7Tzouic41Ps
MTQUNWMCXXb0RfSIx6S/Hyp6r5CKxnCp+CQiMAXnqrswdCEOryQvpojVrlxR65mm
BVJKt3s3MtMSqfM/IfBBe4YVNwM8aeL5wG11XQaxJJ87pkFwBPs+zJbnBQJzI0rA
r7ji64fIK6VWscdNT8HCnbjnskRzSnuTqIvVZ1CI6nCJJK8141e/G9BJM3jp78/h
7PGtCxRchH/3XWg5QcApD9B7Y6S3pVTk/S421QaNJoe5/sUL54dTfSOybXkrFLkd
5+uxN1d2LK0zS2hcgDFPqqfrHnzPWU6Z73VrOPER/zdi5q6v1qChE2tkSyGDo0Za
lJhjYHRbvQWdXu/H7PfrRsVoiQU6vQavXPTi2PXD0SPlXZ0DwdcfLAkFE7xdb4r9
kMKn0M84+m41e+d6CCOHzJJgOBPoxOnoh8kUPFa70GFGtKbE3YnOC4+BV7VmR5rW
e+X64aELEPZyeU2Zm/qVt3LCi8qF+pWNoqJDhsU96PJXNWUjbvpiBLN+kUWXQeM8
IpEzdLFaHBR7HBvtUFpGmn++jUdFzHak/0cLuptF39TfVRHJRJtrhHrMGb3f1K2F
ZRwv9BswfpBW5nqEdRm2xKlMpXb8AZWdsU54AR2gJ5gARHojspxygCB5a2LAdWC0
FlRLLVNQqHI7ny4AX+VVo5uREZDSoRPAuDlTIX6lvkWZZvH+4YIAH3UIzoGjASHj
HCSpPIuuYRe2eTur2aRIO5Du5hWLd+sru+m1fQaGya3RLW8J9HbuOzOTYvr9/0Wp
RmfgUlE+Q6/yB+sE2wVGq5BvOydeGyIltidkLqMaMPt2z1ZPLrqGXMkQEDSh/oFx
RQ39R5jTz2p50YaZTuBkf9Mb70UiRLJ0J8yILh7l6MJt06OvIiCK0v+27ohjkxwA
3KNwMduPb3J6Xtlg1rqMmsdkvTY707ZYaLadA5L4tOLajsr1jGL7+UVi+OJlvtoQ
v8GvKGhRIaNC8ceTkApKFY4mDXl0r5dnKRz6oZm5S4Kayb7Y4jNNjVwyVhr9mMem
VQJ9aYnHpk79PJxxlVV8qJSQNYn6WxjMW0nzz0MePKhh9Bxbb5WO6EZRIZMiB1Ea
iFqLwODqMjlKLHxLVb95Ir/K/6szC8x5BEoY7j9dolPCUZYG2y4BNcMA5NxjxkW2
oJKbTz2pqQi3QrwKT/II2ZNKoEVII8cEfPOyYTFfa6fg7uHFDCtcD5E//nfpvf6R
DvXtYrDjOgTwDX89xexFm/l4mtEzySX89hAGKtfgkItfgYzJ42f4zIH+UZ7o1fLx
E79MrmSez3l/T9FR7HG4u8ikS3oznPjopH7dtmQyVBF/vXkA76Y+AibzyQ3A4ozA
wFnJA5A4RMfXJGEhJ1bq2MTeblZ1mknoOy2yzW0TKRhQxnE2ZKGTFu/qGfCMfbuF
3X/zPjy+Zo29o74nCdZbbJIt9X5lclRCuZVG0XLNKaWWiTKDeGK/U+tJf90QlncP
7hHti0nPIUnYiS3tO8CAxG8figHLS0Q6wGu4sPTRWdtlJ1gryriLBUr9Nsyfxj5j
QZbO1F9dZJpVDOhdXwxLZ3MGqs4ytw61OhcbbrhSjWSSQCK163AEQEhU2l8sTqSu
Oclf6h6BLZ5MGS0IDCT/SExS41voQqg/LA3UdK/YYMYlqJmxcKruzACnRkZcnarB
qtobHk5hw9wBg7xVh8dgV1CyfsWWgM0vGOcwndjiSWNp/vfsztan8NLZIONr7CT/
YVaE2sH2OCOeT/2g9rdLTXgCKHJk8A0AXdCEJ1f1QsUWCtYpNKmldJrrEJhWCBgb
kU6NKmy2jPiCxWxzSuJygWzRFa+7YRvDRc8NLGEudGYd5FL+Rs8oRsQliEooRMyO
jKpSytPb+sbB48cIewFju33YRNZU11hdbfBzNi1d2oH0ZBvCWuaWFBeSRJQny9RU
R9NSCgYCWMHf8EFYApIWvcdjCO19lxiozr+wbPEUg84/RUbr/pglFeKX+0OiVEkl
kf8ZrClJKcdxt3sFl7gQYJZ8WRlg0X1jWqIdpycKIiQuNB8SVncDuhdsQAmOOJPh
xa3sFedj+tTtnd9m60Wad+bbb+mT+maIxK3l9r3Mi5x6i0WdyjQWg8igjXeYe/A8
nQEa1H3jVOIfI4DtoJRErX9I9MrpXdDNj7vxK3oOKRCKttebJUNby07ceuN8HHtY
Bvk7PM+SEJYzAJ/yyVldfmlXumZoGYVlVbJUg5ma/Vdso3hG6cSMQMXxqkrPP/1u
RSGGBBQPC60uySUWP+xgky9wz7yfzbjdF4XQOi4QtCceSVWBMXVlGIaS5Vcwsnnu
xWScqn1+ge7F2WGW5oDxr+PmYq3A35a225DE3A8/2b4Bxg5sZ3zETfSck8wdEOmA
a2Mr9qabKYd5joF4oDnyLm3j9+DHpN9pbpyYKqKqGKHktPLo/mfQ4XvTpTUIpFVc
sx5OWDruCVV1zW39nWqWWvxk4oqiKhXDdnVJRyy4lw4dxta2ntXf+5zJyUmEFdnK
HKAgLITlzVEl7rCRwJpW13L9gx/CbO98gKaOXP+yMdFbu5AobHSxlXpA0pt+3qle
SS9t9hfv0gXzYOId+57SxMR/F+bO/oUmKHcZkLR1bF8dcxJ5KVIZ3hoPOrmCtRml
YErWB+ronP6AG/K5eOdJ2Yt3YqHu6DbsbiYeNgkGr04HArA3y0NaD/XZJMFrgm4y
vwfxu3L2P8g4BEqQ+sIIp1u/BthlhPu0atBo6wEwA2qhMcgz3ynxfu6U7/0Z/MrZ
+0wxQMSqxWtkuOnngCpsy3y79MW3jYf+odSQ9jmjGSNFhjDX+0ZZMq0b7cx2fhaB
49cmotQmdX68/nAv5Ez6VSeAXxDuV0CMoDSA0p7PyZC3WMFgDPJ7byy3rrxWeaI8
KiFWd1+665NMRHHvUJPKlo7ATJNVGXyl966Py69nSjeWiItw2yKFBg4g3vg+srxU
nY72p/rWHpWOeBLyZu+n8cK+kqequ6exBMDJ1V0PjWXM4yDRB5SwFSePfphbpcz5
N7W1h2UPJ7TFmn2bE3hpq+xTIdiV1HjSTACL12gliuk/A2MiP+wFkECJQ3xj68pr
J6sN3oxJnLPlfeUs/tUx65jQDtjbtNQeNREbSc+GqMoFaDHFkC9CEg6kXzkVsfQW
mIY1M1BVWrEM6qwN27GA6f6bgOYpBnItaHpBYLRB89uAYigLJehv8dGwyMmcOzPE
tAvoFXm+agE6DPSo4xChLJ0ewo/IttAX7o+EOC5j+hm0dIz2LSjeUTUZsBMBEwZk
eZwfsjDrwh4CQoDR8AQK6qoMrhKIy4cOCBqV8Nib7Ptyf+9uDIRb8a4zlw5foGKX
sQXLbh6vdFQ+lysFa8+9XK+NzEO5vmXDscLydHQ7IiCBzsLtVjvv72nalAUDalAH
qFuFYa2dPbdI9exLN0EEUzwuSFQxuv4JJlMC7JKtc2NLISUTJLNNHNa90MGcHKcd
IqvOKbYrmTB2JDQ/VDobakyserDC/zoRWSm+0XyDMtjxRJICS1bd+fKKTpsOUkeV
6tZPY26ux00zgFEhuZ/In/h6a9Ylsl+ODitUfZ1wH+CcxLuRl9TEwYi3L1CjjENT
rO/Kho1+jAw7tkZNo9nm2jfwksbvDTAU9PgmyEVdzwuhgrLKmexWJfdGUXVbohep
CmO/ERGwMW8f4b6hxdSZfuAmO4wYz8MZZ8JgfM4XeJbAK/4gKDYCEP5DxNpjQPjg
CQRKYfuhlzUxQLsEehC4Dx2006RIUpU0zl9QpoMsC9U7oUMJFfdcbUAFtoiakKm8
MYEL69WlQFh5BQjz4TVel3cUHJousLpU8fT/RxgBS0ucNrbZQxWqIThZoK7u/SI2
U/ZCQ1S85E4VnEOhULTGqD8hDgC6qGuyolHu3d9jWN7VogauLQ/BZ+abFZFb6U2/
OjWKKsscmIcG4qjOoCqARQ7qfqcsc28/8sjarl+KjqnDX41X47N6Egi73vO8Yys7
1ytwLAr2W0MISIW1acGvM355B0GzuQY6eI5KwbkCNNY+d5t9EMNR3/5ak5iReKb0
m6El2EdHy3Kh+Hfw9xmdnhZAJEC7gATFvfpjP0QGiqfb2pT+vmamJo0G2HMiAKKo
EwHuGYeOAZ/32NTD8fX/YuPSmxH8F9MR/txU4N+vbBAAdRNzmgAyeqm3pD3gkv5z
FNgj4E4q7plpe+LxcspLDAbYzxOMgxmLKOBwasYJtmBnHqjw1C1gzPl2+OES084O
Ml3dflUAkEMt94Sr7yo54EtpPD3y9EIVaEuBWpNw7I/RMUqNWNjLqG1e2ADEbrao
CxN7Q1PwolR/SZjuA2BvAdc3jI29y2xwa697+bHEvmQoF693V44wTYnlCqaOezZN
Vo8QMJZ0DRja260cq7NRjRHAxN2BeflzL3harLWnhKFCWn441QXDY0u1/l6LiB4R
tKUMOInfUcxV23xlgX35A0/n1awHkpeIfHaha6JOvlIn1DXmFjuh9JyK3u0MQr4C
6MYLMoHRf2sxX9O8h/jrLijm+BW0PRH3qFRshbsXvTonPRDVVNrJWJ/wU9Xscir9
HspkI9zClGi/V0t0AbtNZlpuSNwjUn7NmAXdScgvK3h9mx/L0JG8RovdQbPDgbOh
K+l8fFOgd2+gyGzsdlTk1OTEOSQUD/zq643EA5RoeZWcA/OxkFTVr6P043SN39f3
eGOv7DFQBGEfltHkRg9WC8wg0k+harWnfDwVk+dVq99IlYbeF8GpW0SyZBXyZ9CV
1n0wlU5n/Ljo8V6Hlk8bVmnxDSFHNtBmgUPMAsKBs1AAFH1zARcSpDAxWXo+XIG2
hVVOkADk3h1B4+AK5VQmuGcVH9lseI9ipKAxCACDHLPNiDnm9eajAUlkjboxe1Gj
vaBuhpAH/cjl5A3s9olRI65r2OvjI2Vy94ociEbPjt3UAtwFbbG7TpCBkk46d24h
J2KJdCDBdCAa0K2eU/db+KUXO/FYeNtnqBCXBvFFjKzpD3F2W+tzmt8ZN6M2CTZN
0iQhX6pe3SuWFuVCW4Foq/8JLnoav8N51lpZ55Hg/HVvmCUiuJKm9hF/2LEcH3Z9
5TzRbklVRT7pcV6babatPtt423cWKY+6+rwa8BJQ0o22ohQxH2sEswNGqJ5b8n+8
EXpCy2euoQYA3XrB5GprdhDf01ARlz3S8Qy29YQFaUgCVI9Q/E2ex1tCq+wELzuq
26D61mQ+Sbu/UI6drsKYcaaAaFjBR4dIhCJx2tBDrfcopOLJiHy46dsO3TlSiwLK
TkhmvGboeW3vPCHnqDJYWN3WVjGX/uRwBXUayVe8RXLZUxXeOI12SAaqkMVkUiEp
OkUSaBqKnv45mBUbIeAq34+0USVy4JusJlj5DxqgcwxMjh9ZZ2kuCAQEubfftoKU
jqt0TseEGck78UXMZAXAvxT88LbgzSiePELHChpi+8RlnfZuBTdu+ZQmfEtfsltT
h9bZhaBxkswc2fBiLDSERRK7xGJKheKjNoUE0uQrYd2jLGhntLYMolUpXy28eroE
uv5K4a2twkvndepmWW11xD0NJ9Y+hIn0OLze6rQGBlPmZNiTEQ0kRTA1G6/PbjCD
UA5Jc/rJh8E2py/bOzGCF/DT6bhtzDRYU2ZGsEyabLQ8jU23XZ7GIryHOqzo4oRv
RDp1fS+mWjEzpK4HdQmXyd0omGqbSSTRprNUoftncDSnMtGtCbx4aE+egQ6psQiE
y0K1PkKd1uzJJkJihrWC3yacVYj3RPrlw3vJvBXLkKdOGEOF8pqpdYxzNwHfT6sD
VMVS82FfYKGTqlZw2BbRxD2qI0LU3BcZc5m53cfHcW9/p9j7Vq5F+i2D2jDgEJUQ
coABYyzd9hVuREun/45ZlZFec2As7LB+JHNY07tuVnb5RTad6hZsmbI7bxQ5DLKj
vynRjHURl0KDlHBAMxE1w+zfZZuexg1IAyQOomx6OffvxXdoFL6EMZUbuL8aRi4m
j4JnzPZ6nnNBZIriPqU/D8g6eAK+ojBrB91a3vFSNyFmSLNeznRR9NRRr6qUe1b/
ZzNoLVpvkY78g/D0gqpuGHUUxpA9HRuf6KmixGC+hEPyPWpxyzmNFc6yDfrTWU2A
QIlBZZ/p/sLFgLqvB7KIa9SymGK2cuLLkA1vB6uW2eGSEaZ0PFKfw5B6Kpth5X4N
STTuOCEEis4lTHF5qIeZztEZy9UIs33dQQv8jwqj731wYW7oe64BLMj3oiJ4mBnm
0uoGrSzx4EWroQ1V+DdelVHJ6TMx7v8cdAJNndVRmMIS0BggZBgvWgdcEBgYCgde
JQ/aO3zwXgqNgPOVuLCKv4mWwbHcOX7Pki/HFWY2tWHPz3sm69HZtcvw/9+mU+I+
ClVTiooKJWzBqwtnk5Of5oVS7XAQkFGjZ6RKa0+6PsO0iy/2C8CdR0Mkg9d2Jm1j
JFwTp1JbKOIStLf8nfVtOjUNr45Ce1CU94suKF6JjI+1LsaM7nbrksdhOEUx9ekx
QntWQ14SAqZVDNTIQy8BlNNgxEa87MjuS5VsTIxterBc0kqMbk62Xn8kCNn5yghg
v9tNEYZLMONksZY+uI8wuyUy/2LW5zIbkFUr4J5RBJg1gxeGbANc2YSbVLhu5i7D
i7k1i49jZNd+ytTPlszdlBGjU2vf0lckFihQwWm0AETeDexyJFAhsdQpQSc13ekb
VC227SkGEHD/ri/xLSlsFDursspHXJvgkZuB4thVI46Is/5Q7KKqsoXZ8M3XwZLb
edK6VRP2J+Fa7QdTNJC+wZfBElIoHrs+y/Y+6ilUK/C4w1BSHbFBC0v0OBwDM55f
kt8S84o2sCLVBSTMU50EtQ+t3+h3a28zF/nxLDXdEePZild4UCuHVjzDzt7TddvB
IXm8FZkzwhHpZR9mtuR/EWdK9iPUk6VV+LYyvyIeMKNv+WWu9WFwvEQXPSNF7QaX
aPx2GA4oK5VuGYwegPrqkUOWwxsDNdx8g1Sz2EpYvzVVyxlWm395NlFL85XOPn05
i44eYI1VlQpVkblcXx/l9sjh0mk5PGPFuQQy4biiydbKUYc/LJn6ad31FOG/QirR
jWQpfXddgDODzO8UW5jGKaUx0bIuyk09GWIOF9hotPRqEpSGgyQ8Mk9qLYYoAdnG
XR17xBBflbN8TcOc5KWpXuv3vsbibTy+jSuHPg8UVkLnzXImhW/smYHb/+VIoeHO
GdRFnEixkGvvjjM/yc0GSAgl9l8wJjCLSgN5cwnb/Cqul7+7iEH3m5ZUmDbmmLRM
cOkaGwnpg99mtQlYepwWXWD/ntn6s0OjShVe9IWBRftYh5u00lT3sZNZIGBS76AK
x01Jm3qevUtu58myz6Qc0wSgjakp2ZZCOT1UBfN0VYifTPaiTXUZirtB1HlrUVwD
zKc/fYCn8O7HYKkxbBl5Vc6OB9iVqBb0Xwv81Eidmusuclq5RR9GALjz+RsodYa0
7r1TSirZg604rOQe/pHKcP+Q9zP78zhvHnH0jyPG/TK/RIyLHLNFrDfXidq7d/LI
k9Abguc+LA8YyXD0ucvEoBr6Z7B+gI66qnvO3tLW/DSbCHQVTxYkr5V0YxJAxTDF
y3DcfIj0UNZXJ/WmbQSuJ61ooUOu4XfgWccL/Vs2LODhFPRNl+YdcnwoRzFQi8ch
Ss/QZZEq9PemsabvTmZt2SMbAVXCNV/Xu7okTJW6M1R0xrPp/cWnBLJjsnIsXjxb
cJ99Uc0ik0AbN0fqHCKYqnQgtMi6rhuHIWimpuyZ3au1U7upnCcVLV0OfvNHOCmm
G+c/gCXVUvO/LKFt6XpTAO2VK3+PoOx1a0/hNM5aJ0pDUY6Eycy1KOWuF4LRIYDX
mf4wcdpvHTavMBOTC1+uvoMaATaS7S4w9AYHo/ginqwBO2O0q2TCLqZLO0bFhECI
m94h8HlPXZfPxbp2UVPA7EmFecqFYq446NW9qVhDgnc3eSa5rpcfB50nGl/Tm2nE
59cp6kFYVhstmfHhIBB/04jLjXJuUSlRwLw8OWdDS4M9050l/QNi36BMPOBWjkJM
PwpXjETbbvFe1ITvqrJM5fm3Au6MZDx0QGcHI8lMFGZgYSMS015h1sqcRlIeX9K9
lAXLQrC44a+ghbNMYVPq0gcaqGSaF7HM+2QX4a9BQmQyD21zPh5YIFfFrqY/9Zx5
5y0Svq5cSoabQJtfEswBnwdWMRa/Bo+IIw0BpqiU3odg2N4Vgda+7a1FBpsIgJiL
6XcfoWTisIi/B1OBs/t/WJqPmi8JMCIX4njjexiptW3Z6rsiCKlZnzwraAxko9wD
apeMkSUXbIANFVQYOpVmOSGGF6DtqjGNnd+cP0H9LaRd4131BcMDQLhRd5ozbQlu
juJ8ejomggvLINYe6jxeK/Cv0wbjWKfFixAQbygMkrup2BOBgVFIk64tJhS1IL4a
0z4ALIa3pR8hOjY1XO8VVnR7yz+Gy5O1S2XC5Xmteka/hSmXAdsOJWNwAOUeN5I3
sDkeOhp3wPageY/4q5etA6NZSUuKr7Pd78Ub/vx4IoblG4/1DLrFs1V//AI0RoeE
vdXiPHqjve9pg/x3qif8o/jn6gIgvSFABYOc+UPF/cFpRbthOS8dmGYFsSJCHFes
JJy6H2ivSCO8D2aGOVp2/Zuasa2wVop9+RRk+/ovN5zGSoWyzEccIQdwsY5x0+kl
LvqWiLqRLrzaYbh9BrSq3js1TWFFaAczCSj6+ww3WKW4D2OBDdJpzfYwY7eOH1+r
EvVrXVLP7PYlsuEaKhMgzt0O/oy7MLNqx/8V4h8c5ZZFCrg9g8i3VtKQS6u0JdWz
MLq0jesFQfz4bovhQcvhuutdQXtawhg+1UIi9UMQs9YcBxouuQqM79UcSi7yGl5w
U1BRpFDHy1xTLrk0T5PswaPn6egJObblfMJXzda8tyMr1vwHj97erG6JiqZWBk59
iZL36BgHuX/0YL1mb7juY6UiIMadKB2F/yUhgMEQdwnBV8UcxJjA2b6/2Uyg3c4V
bSWlsU9wW1Wgr0m0p3sXfvoCrAsiY2fvI8OYlZGz1NNsjdxPR2ZQUun9AJNPGKD7
UBD+B/RmgVzGOOrifrb2R04rNEJ8YeJ2WMcFiZk8XWpTi8pSU/1tztR7XBt4MmmS
tL71fae7lrXmaGjCMwxsXiK7Lbq4cFLT6lo9ZMO/1tdxl0mUyxmps5GcNyBHjhs7
p6n+bMxRggCk0crwUPZhZFzc4tFZxz+9lhVttmDU0/sXcd5ZMsiCSkFr39z8KC0i
E9MjshLe/oSvkEfWrixnp2keFTb/HYL3ehp3U6STHLY1KG+X4ZeW22axXBZfoe/C
6HIgbMr/Vcsvj3AKrwsv55NJ4Lco8oG8YjOnscsKi+6/7D/lNVOhOtMr6Ha/3snZ
51VAS0lnNN6Dj/voWeqgOKDoZgLqzddhXLR9wYE9I/MYL6RiIBOoOyQ1uzt1fp7W
eOi3OD3v3/oFl0cx9H73tm2DH7Q6E/oKLH1TYa+w+He5nyRj12NOi8tuZOngbExl
j/Mt7M9Ny13ctQtjKO1F8R56ugTbhM/GHjm7bD2mBPrI7QbOP3snoJoGKsrmD3iC
fr8t+ndUUVAA+PRXSf0Ieq6h0l45IkOtbmwRCBh2Mq+G90aLfjkpzmqVV4Jt7PbY
XPb28Xtl6dEbInqUTjs/ZDVUiEU8VZHntlo8Zm9bKsIIeP+pYXbzXez08YOUtrBJ
+ppgWttUgVGYWJnh4hz8F12+2JxsJLtaTW7EHsMct99tkFrMyBL7GpCHzJfPRj2w
Mk1CijzQoqKfN6paIhQ20wApWMlqazECTRJJRKqnL5tcNjhx+CeC6oyju/uaN8/1
neML/37V/HhrC+K0jz0jLrnECgwcS6AWyb+bIRug4YPVBs2AqVT/GXTAyrrCFi1P
q2HIT2YEySlTooBI7NERAhZ+UjDH6dcEhONvGfctC/1l4cubVYrpfRcKq/oaf42a
AwXQ11U/Vh52zRMoNcUH9DZqYYce69HW9aFPreSFgY5L8uQph2KlvxjoO0svH3bs
egHle3mF5hNUCSKqTOWIU0wX9XZ1oGMYs8ShWxjMt2K2PjkTlAiro3mtAzeimYCx
CP6P6punmtQpn9nXwnwXghAZtZBAoxdO/hsh6tIKqKUVB4oioDffOrWZ7EUwI9ao
QZ5xa7xQtvPoWujjGgQV/Or9M2aLzBpKmSlQFfNBTwM6AGfAohW7oO/oSMqwrGIy
SnHzS6XHU2S11/SjonPtxa6q7dxv+nubxHZQ3m8mqti/ZDF0qiMMMxgdY3m9gHxZ
Bd1dA4d+dB1hV7y/kQ4k4+4eyifopjrnCnyE8Xy7ehWrvzllPFW8sLTQHYk4VFH4
4+WGA6CmTaPua9Ls76CvGaiEF8V6cimRiGsaxbc3pNLeYg0QeFcyQnlKfFuNM5tf
QP8deN4uqLdRPz9bZwXuDhsBdLf3GvPeS+CQ5SCrDFM5++vjq9GXQHcOnX2m3mpo
XjColbGEJXRcgTUpuRB+k/H2gejyI4C7WrSIhw3G2riI4Nh1Kqww+VF6MSul8y4F
ASt5sPwb3+cH2aB0LKrlxvqhukwB4FoAAvt2jILLBhKU1hnSlTH6iNfg3PJokgNC
IpxOkUcuYIu1HFMRCxWmHzTaE8iANMI6fGVxoeD5XJOr+LBvHKquRscZwD6CrK5z
QdmXTVZaIu1USkUH7fhISbUljHtc9Tvaxjlh1AXZDMc4NOvSCiolGtwfN++WOBJI
JIM5v87S91yvHN1V4nC9IAEAZK0QiSsbHjgt/mxvBr9D3ofdPMGYNxHMM2Zio6fI
awW4AJHSlHZv7OrobLnp2Re+RQknoYH74UrDNh32RzwbzZynFE6q/gyDtvFZh+a/
NIXIv9OcwlaEr4llm0DB88uC1PGW8OtFnhAp8ZGQAnptTLaX4O9ko8zBdcOijO9Z
DG1OWpWTraME1ivzp8K5uYV4pqGAvfyOxORfQC0X3uGTKr490s0lsc90mx3eouTL
aWmJSS9hIwtwUr5Wwc+BLOGX5fLhQahxhjwp6Qa0EWw9h4EGky1hyUcRk3Qfke2s
ZFxPn4m4vijIXd2i1YdrW+BUNkVPmw/pXUo00LuzWmOsDXZ0uwbiyPg/xMMk0Akt
207lgiFIr1NSi0GExLc2kowQwBroizP3F/vkG1IlU+DiK6MIJBG4eNN8MTtFm/LN
OnoJijiXa4eyo8gFErNQCZfxXKpUAtkK3YT17ISjDTRualDEu9i+mLqWm1eUdohf
5eXhxVGtcwQKT3FFYgVgHSocaKrCxmwmEJduZfL3KQr+EnMjZrAhePmiT7A2o73Y
DneP8xU6Envgg3xfikycwHAckk50RAfS6PT4OYKvPBl7YTejA4WTrqTS0bouviXB
/qCaaZI49CBzDEqtNU09cCRJ9PVbtTwmuzxK+Qq/FdlozHssIRaK1lTXOkwBLHVN
JYZw2VXHSmDPY38Pt8pLGHAMUp5aE4C9F8Ab96mxBivhBq1gxo2jyPpQQ0F9cp3N
d4O71IftStE7hR9EiF76g23OIL9cLKeTnCg20uWC3UupwogUx9ZXLPetc83NISdz
fo+VkVYWuwePbm1RqOHuSB0qST5u+Ao1+MWvDSrSZOwn192nTpdDWqVQSfz7KdY8
b7M1qGMMyi9BXu9HQXGD/JYzed8WDmHB9UPwJZUJ4u5LY3nqAVNcPZFYGf7jKOfq
47mr9HHq6QoSMklq6SWTiI4SmHL0Y/HfZUdQezEK4WCQzBDOnyQ3HBBp+wlo0oPw
wVYrq9/+u/h4FmHEuhIptQDQ3VlMC88/RpaD3Mbht31/curL1mpoDvC81Av5XSd5
B2iY425SgXWFeeDJaEGOT1Xwy4rGrHBzP9KAqjPsqFEw9veyHIT30eqexzLEezuD
qd1yIFVIephgP4fceJGaxgI2bsbG39Yhr5+Ga+avz1FNDAFdx3gH025eccibLrPa
OGYgR0R4CWGwHNZB0KNmOJ9MY5kna0pWjQpqUwofox3HocduH6JEYFxktlXczRgr
iOS0dBAJU3GaWAH62Oa53Egu/DkWRhagZXCjiuLG0EcCH+ahrC5p3+Kp0t231uwa
CQFGoyEAv8OfgkFNITDFTCEiQMFVzaiMTVv+u78junHoN0P+IWoDMzRaTzwvTDG/
yVMccLWSlQQCA8ZtYNWSLqpAIPfGpvNk3cGRM9rZuin72cW6gYN/j8qMdwnsyj6K
6uamUiXBolANcBnaRM7O6ew2/UGTqoRzDUFThl4OmLgfxiKAkS1wf7JZL6Vyxl/U
mPW82kfYJVTgBzVCqLDYmS1BRULyVuHlV2mdgs3lm0jky+UMRLyq0Gv3v2ujHZ7W
EGM9pp+oDMbGHQZ6BU67qkh8JDmSEi0YfACzlszcZjaQ42b+8PmhVtlLdX//5L/9
3TQeyj8ENfBnFZOVE2exsJaXWrdtuWNylw/FyB9iAM/uDvr1BLJUsuc1+7MvgU8R
zhX6Dgo5ZbDUBNfFU8ghyc0stHGNWlWevByLkSYEMvZxwcQwqWaurJOAa9yIdOHH
7ItSfDQYiP1HKKzoM/dp6bCw67J7y2KDexZyLvJ6q+z+ZrOaOWgxyD5uOC+xeYei
VWlZWjR4U5xnWb0U9HmHtF0wtyuWHJE2oCCCKkb/kyZTEyEVmaweKs0Im8WesU+c
h/YHb17cXFdUX9Y99kMlp7K8K7KXfKpAEOg0lQlPz/qegSkD3RoZ80eaQs1/QtBn
wpCsJsE/exKu5q7fuqL/bVbEegwcLvPccf6sjYjVRddjuDQ6O6FfOqMA9/h/30hj
qE5SN3KgBY2oIHpHYGFg/JpjvfXFnhygxnRto0P06QO8neQM68GYwOI5Rwjdtbkv
xtYJm3WQx3dBJNK3aepeC/AkOiFpA4NEFPAWgWvCUVRjO8DY5UXig603tn/+vwt8
wHq6Rv522Tn9ZZ5yKOdS3aCpk0AQFFkBb7nDV+vm2ZjEZ/BFuKANX0w5lqOvalWt
JIzWJfnRAHX+eND5bzpSvJ+/9RtZXxUTod0aI+dRIM8kj5jvKirkwVdk57VqSmRz
Uo4OV8AhjQdmC5VD+uWRjtg1/xuKAHYzZZ0i9cgDMJXLDoB+XBwaLmaqvpQw6qq5
p89/Fj7J77zgFYfEhq7i4Wql/TMRZEQkeOvI4xNywTXHbc9PXhQfj3FccvAn3+hC
DewKbfbAQP9QtXgwpCqtNtM9NDyboL5Y9t5Je07gzAf/kBd2Op+6BUCIZWIrY83e
03DG2y+OXF9r3tOXCQ+IHbAQ/RpOaiqxyz0X///p7IL37rpVtTIS04cj3EHzA1AB
3LkSux1fYNxim0NB345bQH6xYkHvSwKgj6JYnT1Zf47/LsOWAWjDmg9fFuBaWqVv
myV7a8VBalerefD+1m/lM8Nh367qa7BETXfn/b1WuvBpChViONCDzA3eLIS/IpLi
FDwvcFU4PL/b0rgP0MhTo99IbsNBjSbC1wTqO+PBAE+aGX91gKQ6Xzo/49q41dQh
rdYTux/nGYR+SJ2AdobOgYMOKhvEy4sH1Sq3QE/cf1Lot6zeB3vEX3gHil5IcGSm
LTCiWIzQkbC+zPzBdrF8We0HfDL5rYcaLbZ32pZ9tCQ4ljP+jFiZ5mYlLTfxma9x
29s6AeiHqPLi93Qvi9I6aXG/yYdEPp9zcfsOoE6upkZL0TI73etRJ06ANZUICM3U
m+PnHVi+GUV/IJszkzfnCgkhuK7Ble+FlhA1+eq/rVtxfK+8X8VyR7YFW85Lu75B
YxwoP7bat99z18IxSBDGMCa5B0edGv8o5t6Au9JUOII7BGwB9RqWg6qaEyrDkM5S
3LpYKsEMyrdoU6kV3gLDYpdxFPopAR0tKwSrD/EH8HM6hwJ9xwmcbd+/Vi9xqJFF
gcC0eURSqovPrjOZA1lGdVbT58PVYMHuv7r0kwoh6PXwPy/Z7FA0cjAlN6Qpciuz
tBzU4IqeyHUR4YPDQ6lMWmSteoLL905LCSr3xYPbhiYW+GhUdfurjw+lqvBWJsBL
wZtwgtXLHfxVZWeXJFMF/Y47fthXSuUPFzz76AA5Peldoj/4rTEEJAMp2q5Uc0pu
CWvRu2QN5nFfx93WEu1gM+k3KCzitDFQfFUuNnI33QxX2qKYxgCYqpfZ6FIsVjec
dCiNWojTkwSB2tcgMNTDIA4gnonWR+ZjWJYebTESeTyGz/5ZUFJlMdd7NIRO9YPD
YTJb1mSaLeG6PQWk/Se546GSvxk3vpU4RqNA4gGAe6rMmHKcJhyvEjUyqqafn6hO
RZo7MJEeSM6zPpX4j0kkIFsK3UYj3IJU3jLkC68gxGzIFrVAigFuIchPmPzr+Z1W
UzPCXibZgGEVH7QrJ5ZR3eRPeruphZYr70g13oXgIWYcZPttQG5cO/q/UZvrikFw
QSkIp4HJXypd70k4JmhuCBrWpOub9ULWT4hZ/b5Z2teBo1BAw0ohrriX7wm6mzfc
QSB0xEX7FO5N4To7FqCiwbmhxnVHJ49j2hQGoWxFXT+bKjvlx8mO1wSQ9kFisTNI
cxzKmE8vAD4oH1k6MvrGmmba8ipHJui5t4DEySDoUCfFPmXX3p2YsQmPV6o/MFOV
RdjuQ5TKjTUse8Z3CDilBe6uOpjgNUVn5XEC1Oe2saUQzkGrmWHEN+l//hlsrn15
yexIsVcRswXAhrmIHOb4s1Pb+Man/5w8B4CJvTYiTvhtckTEfY5jNVS6TpvHDL7A
oYUVmEgpqwE+UKzBrDzwo6lKDn8YGz+DXD9ASgc/rnDDFIrE7yQs4khSU5FwDnY4
4Mk9kWjTvfs0GASiMoOA9DLYE1Z1bTQUXs+QVc8YBq1uJ5B/PbgY+ub8CedffLh8
nVKO5OQE4LRCQTmXBvOIdKA0OkQohwWePSpvJ8P91ZgJP0tPsgW9pVbe6siTr6to
bJKzXoOxdFoXoe6mg1QyMH/UMieMlX2taVGEQY7mOFU+FI7sQbTfWhTfhqFWbjei
xUcj5Ro86mUAItLG264rTKUQcdakXxa6C4iiG415L3Ktrgywy3D6/2KqCYjki/YW
GHr56UzSLIJrxWIqIYiPXJpNrIXKylisaedU+4+aGcP8uH2lOoIrozpJCxs2kvKl
u9SZPEzwqG9gfoPoGlFzRzljlcMg9Zqg0V/6rpiqKf4enaDE4ByTEEaKgC1lu9k8
KBdoZ+LKpj7k17kqOnxxeuKwpWCqSCg5uiO+4N90043QzMgAQleIhbcUEBKqUCZr
OYtyT6dPV5D/a8lARDQFczt0bE225J0IZw8ZJAFfdh0vnOJ+foayswivcgDz7xch
XgVyeCbjHuYO+T5lHecPsTviTze+1eOAjHt8bskGWUdrNKlxE0SMf8IBqW6dMeG2
ZxRfxlGO11lDFCh5IVEdKdSY3uoZGpKTEjlRK8vp20dxDDJs3Oua7ZHBfQeZyiTq
YEUuGcTKNF+tesRSbotQrlyvy++EN9CzxfxylCIthdmOvyye1Kl+0mDBoGztFG0W
QosZf5szhDMk4Ky/nXsKd6hi958N7+/JUvH0C/jRbz9AuaXWh8p8u+oKDKpjZKXN
aP3/jiCcPIayVQHHu5p521NKSF+0zhtQHHWoIgicnORhm79zHl6TeZmnB9tT44nU
H/DvmKQhwR0j+RzEHFRvB7J8mt5ruCCLuXOvOmIoNYlftXNSU7wG7KDVTo2tia6e
CyG7w7R9Uboc4+3IZAPzCBIn2dfQvMjuZ3id+UBPv7S2uu0KiY+kpCubADLBLqZi
vfai36KYK0NDWW+wwcy4JCJO1hPCXkaqQ9EbyRn1D5QDEK7bm9xTn997NhyUrADm
8YeuVlXNLniGybLhqD2N747fHHb5BWd7dlxkdjqz0WwMd7GZl4DITpPRgv2pN7IA
QU68h2f2KcPbA+T0TG2vAuJt7WNHMc8E+fWPYy7AFFscXnX7fHJiLSKPbI38JqsU
VtQSP9Rt2acClB08kKvW6eHTkyDMUStIt7DoLmBUd/4vW8MMuRdNB+3m+9lRgoLd
QG+AEGG+qopvINhmHhUB0lKchLjWJnpl6vSXhuiYcpKEK8eF+3jzQgUC03QFcfYG
jsYAp/+55iXAOxNkcbVWcsX2pxC3wK8fxjehCkmuwR5kXrumGVNOyr/aQUkwtlUm
7xMDORbBBAKOQijoGNj9TBTYsNwxJ6TiLeWG44c9gaZc0MMnsXuEp6jPWl5Rd2MI
vabw24EDMNc3HkyYgGzR2mXo7FNv8hSUFLlkXsokkufpijmrxTBxVr8G/HiayG6C
NYFnhV2GJSMkkNK50NtyJ10ylE6wp4wiTqhyTOt+zWBQMCAMJid0gV3aIdHUuG6V
1rs2TfRaVWFda253LoQk5e6FmYbnd4KqKfsG4/gNg0Z/JRMHttQtahG3/h1qSskI
Y7nNS2dg6oYyJhQRjTbgmxTrl5dU5dvWiJYgBDNFfBT/f1o0eisVunfXK92WNU6b
7Ji/lFTCuwA8zNZGMJiqAhyOmqLqgLjSAHd692ugdIf9Do8gDIU26XaavpExBo6/
0cn4LDOCptXFIXL9mpu0hOCREOqD26go7tUi0ufQcXx+HdyNKIF1eg3nCWhxqkSL
ByP5xwYBq6k/0k49pF+Ck4ng9kNvPvf0YaPB314/BuhWrLYmL5vp4MdxJD/pC7de
pI2gk9xp80Obn9eMxwqb5rWT9ZiAJ4o8iSB1X1a1vXwX+PaPBYOpTS6JY2B5vu47
/rJFgMn1JMNGeBPpx7rTO5WaPpyztC/2x7pzPQumkH/BY7hixCNfO32yJWr2aaB5
XcmyVnAygfZb5llDpp/zSPEYDS23CslWdI8A2S2VmGCcdlaSk18WAtxlDgPf3wZS
ZU5j4/OU/BmmRYLI9prjDBbo2Cjv6PBcBPROzbV7JZPPcm1xCNbySs/j4qT7hnP/
9NyOBANMCQAUglFwO5v/AlWJE419UzOHi2jFt5tLMrnABJijTgw5C08DZ3SE6rww
0hEifQ2eZfOGoR6RmlPsLAOdn/WHvy/hZQgiWT3RWtuMgWGaEYeavyCWMLQ6KAsn
zA3thHXjf3DMX9e7Zljf10nP+v8tfZvx2G2S0t5/wzyHYFYTA6KEt5kzdXCMfVWJ
h610EictoazEI1b5hMGu05wmm+V0Msec6RoIZHTDXdUh2oBNop4viflEgoCC5noN
hWHPADRqK33ToLH1TIBv9elu8cbQJ8Y6J1hiBJw15qIaCr7KTenBEykX89ir7KR4
AzTiWEqi4a++ExgpRmctcwYN0ecK2lBro0QgOGVgskKocmAoItVa2/g/y+RDnSQf
16iqnxg9q9KBoTlSFavkOLztLpaYiRC0gywetPJrDuiQ6gc/wDIVjFxek3ggb8hf
Pf/p6HpYG/KlTDSzi6cBgQSl8vqbqn59f8rBFSZs1FwZwnFRDA7C1F4E+06J/sEr
ex/C1OTS6x1KHpEpjDZD7JVfGf0nvgDE9DfeeskdAdKmODZKMieniZsBxyiVvBvr
kk+5VF/D43+kBjCGH00LiusXZR3gvhTrjfAJJZDOXK3iWdSa+JIJ1CDx4GMc5Yvi
19JQGz5/SNRkhm0ieAx+XHKBCD6LH+i4Pj7M6sFZLzkRNTsGGbgeFwly/7NlTSW+
db1d7zhbyead5u6RP7bCcgHOd2XRL6svgTE19RF1WoOAdPyXaNNQ6ZVeTSXXq7bt
S/QO+eFdj3ZkJ9AeX/KZQ9i/tbNo2XtoKMYQgbnegxEqUnDLeMQ0vkhl5V8CjVld
vh0MBCwXIzIQkUOvJy+eeNyXP3v7vNYxHiIMsSMXFanPRzKlZz0Dzx4hA1AWp9ZG
RBWTKYB1RpsiY2YkB4NgjvSpuZ9QsU4DBmPCR75JKlBmsi7+tfgzijEsH2KAAqNg
1zN3L300AZkK0sopzS4qMgDKsmAGaCmf8VpXyDiZuem1Jt2zO4lfYcQ6zU7zOgib
23o8DQtl7ocqy8n7HMEexjfYUtLoFy83kP+LdtDulFjLEQgzjpIK5VAZ9/8+SJOq
ggs1gk1E9qzTr8MdLY3JO5K3LesV4hFSkquPdt1ScUd6XjOKS1YV2m6XOVAxRjBI
Bc9dpQ2wo0ikz8NQkX5pQq/+9M/6blcFzTMwRTgN8Lyg21D0dIiRptmgpLcCcBW8
qpDofml/H0s64wuOK/6NHtysi0dEduxX/U2CaB9rrbFVA1n3mDIZvwb1Ab+VrfdO
oeRlU8QH6aD4gFr9A5859uvd/RI4HfZrVOCgOoeVSD4WWWSD03cRKF/G/GMCuhtM
opiUYZ2h8dCkLxcquk/ZnslBeEVjxHaR1GylMXgwPwHqikSOof9FTXVmzCHVYXLR
tM8nEFjA1uR+7B1WWGxT0k+HG7yPoN4LQoosrnjRf60GqojJsYixTD7WBOjSGqX+
Y2soJcAU8Wmj1ZWn/aod5Pu46AzVjwVvb5vC4izfIvCoPm0F/f24Z+9DJEfJtmlC
tya2yTl0yJ9dAV67MnaGv2j0tB490kjNmShB2pJ0LENNeggrt0l5U+Ilp0u/hiXE
892ru5advuRqYNpZl/ZLa3mijCt/Od6ITSnUhuPIjyFDdBCzP5mEhuHj0roPiDjV
zXZBw/s5rtBYDT++3MmC4cXM6ht1OUXeIZJ9lHu3zjCvk6+vuen0Tut0ekb1no2M
FUOfEmkBsxDoHFXS7XKkMtEunT6VhGjsJDZS+9e7q44qYMMIbdidvszK3i0bDYiD
STE7Vf6qeWQG0EFjkLmAwPo0fmApER0ziC+pXHBgMIlbCHXtaXu2PtHSVk8uaIc/
FcKOXcGzIIWQU1HGPfZnvLCdgg2NcMYYMcb+rPM8u0oRTft5EhQjbY2heSg0BmpO
gCmptFqhu1NeTebjOFji67MXAfEEdWczQGIa7FS8Yc/b06ejXRkiBDE0ZanpCN1K
KcidwUeWfCfaQJTCK8M4OWeN/73+NPwl4GXsfGe5glphx/dKe2NCipnbCn+Adk3f
CCISf24VVlbcgPPcDhhgCo6YMqqW4214fiU2byq799mAvPgOs7WrqzJSOXSlfiwa
CI7miPQMch5+GUsXaT/dmE9eygZoCKBgLqcPeYbst698pC7EdVJRcfXaHTrss+JV
4zOubBjP4VwNjgpybQpg15Vysxq4hjxTMkkvYMmTO9idXIC+KTABNMw+V5YXTQxH
UIiNmO3PQRnPbTc+ud0CfQUe85XcLxFgr1Ul+OwtsBHUBGrLbiL0KOuzfBKM74t0
exQIFjPOftz58bHeJb+PkzX7XVxuZGs6lgNRNXOpOeonhMJ2FiPPOV7PihsmMUgU
Dh8Xfu/TlmOe1ki0m9PQsdlkV8U58df+TDb3QwlseE4jOW3FmFfVvwz6VvwWcSF6
P/y2g3iWjVie6R8UgQ68yKwE/10UnWNGh5PFUZQt2PwtDZ044Sw3dwphNsCT5bgU
ld8mFIB5ZJCHc30rcH0zgm1DIxubCCi9S0SwbhdBnh12oYc2q/xGgmbgGFAvwHOT
pJBCa58LXounyd1eHl7Ckceur825e6m8y3KDzYy7Ztfda64akeuC+ate2hITtdEB
fBVxgWdjSFw75sTRn55nd62/L2bLnOJ8egFImEYbs4eXR5T1+bb8F4L1Xwxcy3z8
W1N1xITDgvCZdzTCG27ZgL8mrHLpIqPHdimqx4nB88xnsiF7K0uC7fc4fijrCYs4
pOzIICv2kNAhOl60s5hxvc5LPkyD+U3oUVcVqKuRVMNz6gG/E3n0krhVHgb5RxL6
EZZxoE6K6XkTa36LpGatqgBA/w+nKGgpna+BUEtX7CDS/eGLbXbvNCuYZjgVzfSv
SgzIiDyMOLiewMYtEBG/bNHwqW4FzjLiqDnPLrMxJbqo6YneZVI98fwzkpMfxZNL
POHQNasrRfQxufUp2VRBYYt3ZL7YacCCbtKVDnjumW9BfF9+Jv2WOj4LGr2zovcl
oupRTxno6V2zwzi0vH6FUD6at4gvt5dDhWr8XQgADvTnno6t0UN30Y8CPwTtK7lT
VQnKZyAlNeaEn90ecck5hBi5lGLVKyzmjcNPm/uQRl4+6b5zyJR2ZpeYGwFcUUJ/
mA6mq1RNy/UelOVkfI6Wy27QRgj6W/SjBPppUw8bQU4RzVjz3HKikreP6KvD+w1L
JxmEtAnvi86NKNwpx5h6tuE3nDfi/eTO4zkLxx35lHppEusardxNGPH/dNV2Hc+s
Q8F3+94Av2vxrNSZDlnmkcFn96AxSWNC58RhtJ/j7em0mcf2Qiv+fghECkF5eJDw
WAJhF2U4H1inPylvEkcxzNHdkfrl4LruD4XiXpUZVka5FDXjRQ0X02unkfFDMNWk
m+gzvjWXk86B3PXJu2Qdq94W3NQOQX0HC8UNmK/VwbMOc3QLCh4bpPX6seDd5dHz
QKJJcbKclxNDbwQt22Fu2wfv4ZXxW3MBKYCF3yeznmIcpAu84zWroPNWsa+zJdOT
cnx/UT+vCnFbYI3VsQer/zmw8lJ10tWZd0m6dgJUWpjSURnB4TqX7RUNzunYMqns
tzHlhvSY40ar2okIKlSJVDrlBSnz1bSDFNYcrP0GrZxVLBQwDRDYPsprLHzFNU76
snZeCIz+LGpYEURobHo3+z/fkfrpt61CuNFZORbYL/lijuHuyNwcglAIHlAhJ3k/
13rYyYjMWpNuhUVWluzgYchUseNVqY4j9wsoTrFuwqNR7E9Yv/V1w3s7qsKWtyk3
8iTSxeUQ/2F6zGFvE9B0NsNofs6aAFG0t8gSzNyped2AtJVCJwta3uYPPZj52CXG
nYIPNc2Hj/Tu20ziui/BG2c6aUIFi42u5WobKeKy61+onqPH3wmRJHf0+PPKeGWb
sHv/ELqUHIHWqMkMmqzmgAbtgGU9ZzGvmQ80utOiuikD+MJbLn8c2Eyf0wDuEdsr
bT/vNpjPleVSaKtTEHSvRNt0SbTaDE3SQBK98XDBGWAQiTQ52FLSo5lW8EwRfu8R
MlbZatZ5dsvD0RXeyQmoNx1Oor9VddCt0cBEXxRj7TjL6wAew/xMboqXXX/Dfu5Z
E48vdtxcRNxX1VO0j9Im4xpO1apys8n9xVLeOqQaQLQGWTdlreuO5LvhVXoNmxnd
EVePJm/Ir1tAZC/s5xMTLRUuqv9AHQsyhVAd4Yh/JAl+I9rYS0yNyKKea3MjC2iW
j9hJ85sw8mvgLOEKa0ISRX+H8q8HlzdatmEcNemnGlALDa5flyifaCcI1t4+9+GX
HbdZ0+QSD1bLSUc//cuTq4x77PkjD7Vf2+bY2gVUp21xAsj+HOEE2oCMTBDpA9MR
lWrducuiKU4zytMindMzNxouoouLalkDatv/AO44ExW89KEW8Ip4uyZam042ko3o
/uaYghLSjbPqaF3ivknkYr+dsRb/DpIm0C08M9Bc152w2l9UbV/6Snelc7fyqZ9Y
8xOD11iZkQbOcbJQd14OEVE1pce/jZGmfYF4imDp1Q0U7guZaoGkQak0K7OW1hFu
EINAJwqKo7VVmrIvY4011DJl4i13lj4pUdT/jqvUwtJaQioD7OkTH54HWzr6JrP2
3Eg6AGDOZakEDPMoLbnKNW2yFieVsHftz7pTJd70OIBE09iWeOrQ1fVM1hnkx4If
JKN1G1AFaMvSKbkJqujUewz7zLULVUxsZhAalCNEzwjjCpOjZwtvZrzAGBJM03iY
fV/NsJY3V7MyH78MoMc50w+rO5xGh0A++wRQtG7cMglaVCytImU0gr2TOxptUdL6
Cj0G/9ruiy3G/p4ARrXviV6aCNy93Dx8xMyhzCLpK13z2PW5juMCKT9yzKZrp7Ka
xJ+bWxmzQBpYApNXXi6eQ9f+6pgnN5DqXF4ZF2WtKt4cLsLkJTfcVmfXKixSZ9Ej
vOa4MW+32kxQBBpc9uUbcCM2781sH9wfi0/yRikv0W1qaiBUKTGeQ2bFEUzQvNut
QjN1DdC6Iw6mgdbsaBVblaeffKCGGADLw8NQBURzY9cBdLQMLMqIRmyagayBJKLc
/0zSApDX91b33mTA6B5azLRIJKWzmxnX6td90NVRZ8kpijpoNBqwpNK5yIX/gd09
x2u7Ye7KkIiitkR5RJNs9hqz+mwAM1wcxCjqqDEQV4RIXHK3nFKc9FjpXMz+dt4u
i22fuo8X1vtFQlhIZ3p45alrpsGHmx8U5Ba29VfKUeEagQ7S0VHEl5jFP4iq2FoG
88YqF6dSTQyBF/W+mqGWZO5QruBH5MJcewFJjyuccxy6FJ4FCvct5BOY5qssbwAh
TNnehU+LR2BWIdOjkbSMYAoNlYJuwUeKrZ5TpkmlsPrFe5Y+OeIzfThd+G0xY7oQ
O0YLeugcZxhbRzRpFnAOu23ExEjuJWm2xjKgyoO+h+SoS6y2JgqhmDmLTMR8k5Ub
mgSZXtcqZoMgG4+pT5zPGqT1mhXzz5fN/7jL4/3JYLVAZrj32aBkX1ud4nTGLWPK
fhbbMIuw4Q//3PG2ZE9Sjbqd5czz2y9vKqxbMDKPk1t4cjNQMXUTI0lMnIJni0lQ
j+N3pGoaCSlInXSvvBkf2Jbmmtb9WCxM8d+IbpFQHEe5r8EmIf/+sn8PrDGK4gCe
x704o/YPhK4eFqYIvGrtE/DSvQjKsUOI0HLMvmVd9G4MlxL73OwFcsknEYcwxdWV
DytvQFb8C3+LldiG5NYV3KIHfhAqwfsuEpiPSs36fV9HOXvf1FKpNgRk1RL/hgyN
+Q1E5FaZ0D0Q+mXwdnOmR5R2h/2h1vZcwRnb0mNV6Bo2RZUm3BYYzp8nyDkwq9BF
6+J5tARfdJLs6nQPPHd+KUmKaRHYrl4IMQWh/nKHBm7FYWbjtHvIDhqWifqqNug8
5bOz5ML5fzTRjhTMmMBOfzhkz4ABPJm6mjPgTkg2m+CF5YAj8XzRRX1qPzB2ozDV
Qz+WdGTwT0aZ7z6G7Q53w7JDA8Rn+wCw/8OsUTdag4PsOjjhZGmqPH3oawNn/YbC
mV+APzdkcjfd1e3sQAXAC4Pu6N58AcAZrcDSwWqORx9hbBvcP7d/YAZCcLJA3Uzj
30qdqaS4ZAOCKzgMkHh7uVYiaHdnoCoqhlFhBlwiWv5iU8ZIQ6rPlmmaY/b0mB8L
0P/NL51ZPXe+aOrk0wZAlilTJhRoPrxMFFgrgCgDJULnwsTOU6uDzRhp5wTnz1bJ
Ht5vv297u57VvH01OL38AAdwteIv4tS8ElwZMPM7Wb7bfvEdHkoit8wZVLexz83S
EAoA1kxcmoz3ufa2XoxFIAdAJCR6bsa7WmWbr13cw8BLuXD6qMAu0bxCZUBNPAuO
e2dkRNfTGG1bdG1IfcQuMz9Y6FHoogWK4yrTSk4OSIZ5de997ru4G037BCZB4XCb
AP+Qz7njPq4nuzMU3taMm+QwO0Xty+KP1k2sqcP/iR8vvuT7L7WLj6nwcMSujKaX
7QEroxslvl1O+5qPv88Dd/cDGLubkc/1+hqkXXXhQk8jN98m+frCvnBB8QEWv1S8
4iUrl/C2cZa+D3De+BduDRK/+mF5CZLSY/5nCSTUAJI63UZFmylwyVHTWxgJ052u
oblesHsqPC1EqrhFpQKfCUCxLfhjrjs7tpFqBKypKknoETsf3K9it+9DARqqy/Pc
nSaBl5WmkkpFbjeKhPZgU2AELe7T3MEFk5bcd4b1uzPvSB+HNWhHHJlYaBrisiXM
NOOPKYpPXY8n7SZCyWwDRU79LEW0pYNwAQYdIz/aFLHiNKb7LG/ZWS89n5M2XY3W
PqgoiJyl5pazzVS7r8IihL2d4lfVZxaVn7v+dH6jvTkolcRv8czRdw9eq3/xxwtv
VPtc+IwvRS+rE9xJ0CkzobYtUP/mF8cmO6tHnyJKpAOSnkdzv8ltqqjzqlQHNkw9
ivGiimEpqdOqSRscNs8b486VrGdq/UYWyGF0igN/yEaWyKm0iiOBFO63qcvnoSQ8
FuF2G0xJy5Qvxy5MSJ92QKHIncZCM8uZM0yXEiyFmDeoRcGtI6n6AcEbI96k5s9L
0iUHTCx25Y9Nyrl/Eo09u/L++s4kpv/7D8/yf8iquyzKMtyXb6X81kPtQqzRu870
CJkBjjNsj9I706kTFmseONg0Ii25Tw9lreoupu8Ffmt3IUDWo0AsdugBjK++1jr/
Wt7gu64+dLwZJllAPmfHEJuA+LGLfP4AWu+1qB9Ms/aJk5yCGDvgbKqIqboARklG
SOiNYBs5VY2EaR678GptTJe5zv5kQdie9NBLJauuHNLt2quls9HDda4jdRiUsJgp
uX4r8nj4r1wMDXVj7BwMHmHvRUMiuDKALXcGCcuqLs8QUczZkN6hm7B3qQb7gv8G
lD8sqiRScUyDdd9JswLtCktOsIHykpOdb518+asIWOA2BMOc5jPTmzd8flHT27IG
mVJ4IeMBJo9nQ1QUrv61gcwM9pLP72xw69yZpzwWUV9VUA5mrsMankfZRUkx7uJi
Kw4d3SotDpJFi9AkV5Y7iYv3JWvQKLu5kK8zzxRChRAV17rBfVxZEwHE7PNGW78N
7LHdYC9EWGBP8CtPPEjoNAGvbESoTvsOop19P3JE1jCyjRx5ZqaGF2Ws7CTeTFk0
d0PonP7w8o55a2Y482a2wu6h7ZCv3iU/I0PlMpq81SWOcLQcd2/kAvro+IV2Y355
qEqkJLtkQbsBjnWVoHYcNCzoUPPtp6ijdxllck6V+6arSzmZtgEWwu2L94QE8/XT
AV9n/kxnpDW3irCYF5W7O7tVpaBfePUMmAya0pr0CGNKTeuQj7SuGeF5q5dk8LJB
71oS7YIIh43Xy7w5GRSYlClSm64KZRSBF05ic11w/bHTTtMBLUn2yEkKTWQsgVlQ
drhCGsedfEemDcYCDn3eCjicfp/SpyEuBGEu4kcNR9X/TeoxOjnxXNviIpMngi5B
6uI7CAlZ3dHmojj28ldh8iLgfgkS+s+Pjev30MtkVIajJzMCNMm2BJVrWl74qjmi
tsEs4MCu7Sv3Dj7f6s5A8FF7bGC0jnS4DI4iIbk8vNBcYHLaCzsDLVwOpzpGgZ1z
L+jTDlBQ4g9ByXHazj67E5UDkKnL0Fem+/vDPa5nRRR+g5X1HXWEi7W192MqFGMP
tMgpEVAue5jNxKASFyGQakpSPdBbF7IkzUjES5vjDeu4nOSiJvOHZUnPrw880HE1
BVukbe9oBUkO31DgCemsklu9AUyLW9gikV2LQYEacsBaDdEhNeIkPtth+xsoKOm7
Y85Qowqx3r/zGA0gEuLvziwUKhPKVD3Af0SisEnMwoUqbKhu9E1dXdEOWUoKUbiO
K60Mwhk6+uPiWfks5ji7ZXDbw4LHK8IZ+AkB+7zqdt3wu43mBIBIfA0WaLoS92QK
cszt1+uyqlSHCv6cvJRC9ELB2ubQyZHNTeUJdQT4oDGpySv8kPsqEu5Bv1SD5rm0
BeJIdySDUCzhHcS+gwS9EM/dIvyV/QBgGsLEDph6PueZft8+yUQr7TsP9o12K+fC
KduldXD7ukfcwd37W4jvEXunKcMmINpWF9104hxWac6NnQPwgXlKv2zZoK6OKkqI
Bqfy5yudJ8OedUvY1XtlGOxsAuNQKNqVaIWCDOc2UusP08ApVUVGkiduzlvhheE/
JVRdhtOfeK1CwKEpxOJViPgK0SIC5VsvYQb3fFqOHX0CaIBKCZT1XkuoUF+DsE45
OoPLm913Jxha/zw2mEUflXKrden1VZzcLeg2T67riSY88Fqa04FPrg/Z2D2/OPI6
Daw5tzJLmMAZN3J2ufqoQmz4JYDpVVZ07xR/QwwREVSCs9W1DdkcSSbo74q4/U6h
zzMamdggg5w8ysjPGEaUkNAC5lC/qrWB/6VlDwkTYXqUehcF2/45ogDmTv+YbMc4
6sFvcbvaYZNqvrSlz70VH0kiGj+pJWdvByKVjejw9cgpb7Br/ixg1m3i+LQEs8es
o1qDVFNj7IW7XqPOCWgJN1N1pdGL66U8lBeh8y/TOkcp0lfGsUq6a3JsxDUXbxX3
olfvtiUtOhUMps1hmhmUpDWUI+xNvNYlQyHpjEGGHOSaSxFH/bWfLB+A273uLDot
KlnaL6kVqZJYCypOkFI9FYEpY6qQ6cqBw2Ix/PAUdZcBoy+QigHpcEX6TyhcLLI9
X2U1VRE+AYJLhxRWU3UExzFdgHB/MDsdm96svM5k0henkNfoB70xxtpPW8isq3PO
YmkB/V+2sSH3sp4dZ6PojMM8Y142xdZRElFBmG20XMFU0ojwctpxrbHzE7mfF88+
e5MdhQIG1TLOsBgDfoC5vIPx+kdGZs0DbVL28B20t2kQ7qlLBcmjJMDHg/AldRHq
0yHn1Xyop2wVXeL8hZK5x8G7kvB3TjIGzi0RWrEHkHLFQWN2xdU9JdMwmoJJmaUl
kluKhRIyHG1xnEWNIEniek+DnvwHyJh/YqW0f5XGmcoQsC7g/GRSegRj6QuhxLYd
BEpsV8VFUbEH+EU2z/BL9iIhPJ5le5INzVR06yTDLl7qqsCWvN17beJ14l4g9oJF
aKKQV37n7ZiutJapK2oz3NcMLDS0EWm6fL6giCccVM7Y/L3JWtPxirSxEp/2Z0Xw
8EfwgpYNCxkHYPfrGOKtXFeE7YzwEC4javTo3nKJr+a2D5CE9IC0t83TcJ62E4Bi
cs8tWo2a2pe0/7HChHPMTdh08OpcHmcZNEFae4DUWmZbwlZMz9A+ewwW3mvHS8UI
nR2ta6e+hqO7krr+bLSW1EhZgp1sHVlZjHEvc0dAMyUYYQ2c9RRGBCA54d4Lc5mp
VClihhjLE2KoHL7V3XUsEm1h8lK8fWlBNHYxnqCgRAeHCbj4PxtA6N6fi+3D19Qp
7iEEJPX+8ralXbWWB7GFQIoFDGBJmzSlZmYMF6t0Ww4PhFlAkmx3knhXEw+1wxvg
q/9cq8RC8J/ZXVbWJTvjwldjz4ZohnrNlrQXe8aZDufJXdgFU4eNu0H7Al/LrUJF
CNO+kFz5ZfSrvkUu541T76KhNjPP2LKgljUVDmwBDkPbD4p8Ul+nCbfaxdtoNWbN
JnNVxJoPODLZvbBBuPnTGSKFxwDk9bFUKA7tTpKrkJ8tb1P+I7DFhCWx9teqwXat
VMYe5XG6j9UkPcfl6t/+ZEzPqHNfLYCYimEsLUGdZCIIs0TEwdAMcmtSDlxV8xHt
/5ze45or/4t0jqCoU6qfWr+ANS8aVDHfOcR7Mjddp0stpgXz7ZrxEMZFXNok1XAz
DOHI8D+CAY1Rnv+++EcgFnTpD+1J0rG0bbRp/jMMJEdmVK1dk7pAcjsD/lGiLbf9
vrGf+iTYH8M+v4KpDTBSfnq8Vu6NS1NFNCmPRJnFlGJa5QU+Jr1bIsa5iW6DWSWz
370SmekLRGRTcr0by95KYNI3vbYQs2T8YooIKzFzjluwl0vEdIZHisKZ9SxoMpoA
yaYRn0a89lt+fAkxadB9m6OVy8Nfd2llOcStkbMRtHpW4O238k5w2At1wx6jUHqs
k7HYkn0Vm9Nrbdghv05thQgQt2iZNNbpjR3Uj/0DzCD1XYy9RO/xWiObIZ+I06yb
CGa4jJEmQMIZ1T/XBY820Nfk919vIwvXgRIEcw6o7XdW+cCC72lkpi/RMrJdEKwi
6uwd07uoYh/ASdaTPRR4/t0bIWLaXsTsS6ngdiKvAtBK7tvC9JQFeL8ColC4PrQq
kgl5BKNSI/2OHjKaRNUxQykwU5g1o08ebnrfySG9vUn19SDoNyvDuxUbkB0CfPmI
6NmsK2GDmCxK+zk451tSX7u5pzXpgf1w55qlzMKtrhEP7OdHylMjmEI9gWcLngrY
2MYC9oz0o3tcaIrX6YgddPFNDpgQ0sLUydLaAQBeXjQKaFMvzszi2DRIY2c0RkNS
ces1Xt0OhsVvsfBzCPcqbn9pQYYZmrQAsszEsnzvfiwqMeOuD/+9uA0cslwbFyoT
FOpd2wBTOvgvvddWu/HqihSYGGgm7QQVQWMoNYEqu0ZyPUSVKeQ4r/imZbRLkrOZ
qr9AGTQEdFuKnCbwAB1bu0GDbG1oK6hVfVFhdqjqEIPnMRRWJALeI1JcDM2+RvwA
pZMyRxNcPqLPnWiOgTkH4mXZqHklSKd9x6hWuuocdmqGhez9GUEGC0TgUr4HOU0t
cM2ssyDKxsljCf0WPcyjwAzxahfGix6Nk+RDWS/Zr1V4BXIsemyuOgFf6VhklDpz
DLj07P5CsEgIH7fPUvUcmU8Et50D40yUqLtEXlIQAqnslpCdjEqO6kjgQm3SoYN4
Skwc8khy/ztm/8dOUpRl1cQXrhjOBec2XcwgiJco1tMumfq3rj3n4PzGtTTgsxM3
X+qUR4lpEHaoT+W3wwOiv0pVcxpY5o+C8SlnZ7BZVILoZAiheUiWuQWyCL/RfrwT
dKgXfAuDHSUl73L7TY3KivsCCoSIY2RYBPeU6VBgtcewWJiH21W0Zf47LnAJN05f
yPRze9CGjQ4b/zAlhv2IOwJRg3Fr8KkkAp2zddLOo69NUzcXrCD9zCHSH7Jg4CpV
/OvrPinBZ+sTa39Rf2Oydx/KrqXsH4bOUnM0gdSqQnwGaKcW1S1pAmLj4LoES2Op
hjQjmLIEyux3nmoBDyPgPx/1AgyDoj7C1Hub6ec/iN0+wgV3iGR8SRfICDzMESty
kUZwNAH1TKz+3ZDCl/oz93C4tfsM4jIWZA4cC3Qhj9Wuq/LVLVjCmxc8n08Lj1w7
JBn1l9qCz96amJuCrzuP/VaSuIBeZpyBtGAS9w5SKxJqcwDcbO6Ef1u8aw9/tb7T
CdCCx0Gdoe7p7IjJ8iJDC0jqDUK1XbBIw7DF8KNzNrN7W95eS+bIe7fSthJOhhOA
u4MkDs/7HYLJY5WTtO30YFt/Nk3PW8uWidNgSzHuSu277m1stQcXXJJnp03or/T1
bLyTXx8sG+PhveVRC1BqYxZxR69G7fQJy99gxN6WKmvcegceOuYu5drcOKZnnu7l
wHI8g+mdodK2Ae0E5IRFRW9ZoAkSYggloeQEEf14e5RSKHAKjEdKDFPi6Dm5uzHN
hXWc3sUa1kOPWbGPUZSike40AHlJhBbonkpz8aulhtWk+5h1R3CpfcJGLnQdEWAO
k6VyWf0ru5xu4jr0WKn5XrbvcckNE0ujWzkwdY2cM7lbnLHov4OKuVuhuau0rXUt
Y5Rp3P5xethWux6LQPSSYI11W30RORB1QdnedDZEghKnP850anBAXzricpQH2/W+
tjGg5CwcCsUX1siDVSNoO9Q8Op/A0migUUERPItuKd5XUJMICRqJLrvbTi51zM9g
PBrNa5GE7Kw0uD9ePvIqu8O/KELQ4GIsmlHSjd2biVuqBJFIN6u898cN4kkyiRvy
fjzQRKDsNTY5574vLK+KKVjVjMEKQ1tT4Jvyt+euZgr3OKZMjDj0Y8xnpHpqtFzA
9hiwTFhavAFf0eh69aYQZl3kYVJO0JAyYrhPtof7j5GMdsglCMQn6MPICw8Zudb3
rh5adBI06kALMQR7ABA5tfSQI8rd/g9W5mL6T7SmkRtw7tH5hBKktt0b1Q4jpBZy
GSVmG7h94gUJNsZaFZQ19vx3azEiFQLMwMe3BhLvoNRcs2Zqvhy7D5itz4oBD5rZ
No4HUQcL4q67xluEC6/SkAt/VMOxiipMW93uOLuZq4QECHaOf0HG/Pve2BWIaCAi
B9kTmmr6K6zrsFOb1Qvusd5+mhEI5iocAVqwLx/QXyQd6fOJmpvPyMYea7xxN7HJ
yUkzg+ZVbVqb5TEEXlJNN4TbPBwU/t2iVLAeDDHieDh2uks5pkv6sDdywXLC6Kt+
nzlr1WCGSX+Bh8PdBl4rRYxgmbbAmx71j2FA01d3zx6nWBSIUGYR1u8K+v8cCEtL
iL4pYeipQmZ+R3qirjle/iVHhl53NzrMBP9pImMnvapDvlrvY4jkij3E66xr6W3O
h7Z5vIL9TWjiCCTYH8UBUhO6/mMUQnw0KxDDoAVM7gMza0QlKkzNIO4iH0pWxEJs
DxIIEnSOAET1V3XeU/LpLM46/hzYUDd64LP6375O6yvUP0GQbqceQFKqd/3rjV6f
d6FE0xyyTttYrWnnT0sILS8jKG+l+Sc4J1xHYKDI4ES2Ug1vdvf7XYP14oBQiITx
4x0Zu/EbFLRxKII7DdL5nbnjPkRF9nutM63O1iACjm/CNxtPRWJxg7H+LXX9QLE5
hSNfyoUvv/2U48wT3XrSpj8S3SvrvfK9enbGwv9Xm+7to7NKO8DXGcfYWcH6AYmr
Y06v9cs5fqD2Jf8PDpJN9/1zsCQ2WeFCzx/MkCgXYR712D4fVQ7Ybpmck14b4XP1
pAKqh83m+ANB8AVlrZ+bw9RHz+OkGHBxXeVo2pq537EUErf+zp3/SzXy45xh/wdM
06h/feH6BdNNK8TiD1wlQzTa8/nyx5imS8Xvxr26ZfX7NyXbAqCLZ4ISFczX6GeB
0QwGVkxwNTu+YwOMS4IBYL9rPqxSIXcSfWe2LvkuZC7dNwxA4b9MZgQkhRV79ECK
7tDQQLiETXc8Gf+l4Ck0DCYOJXNvgZGxP0sGY8rBxpj0ry/DlZ5Hw5GdB2wSCktF
WgpgYavmMglQdgpOYbedZ2X1UinWWHaxNjT6Xy4ASFY1n6bj4xPyHDARxYs96ZXX
dJwjt9bK/3XCV6gClcGXkvjw/W25FD1Bj8iDJOZ98hjzw3u0Mer22AGtqoG7pWxo
iFgpQrldsRK+TZQR5XKy//RUT0AFz3r4fzFGHnTWEZFWgd6u81dzabnJZicWeu1y
SpKbiGm1c3rGOR7erj3SpLoW1N2UfoH3BnJ7Nb7zfRMvQzM7YXHfOhKHbz+QDGoG
IHvTkdyuui6FFkrgJjQzJAZe+HvWV/egZ2+3UBa8ex+BJLSNsXOjl3tdMuZMRLLS
qe2QsM2lTrw9xml5bhQLwdaQ7iro5u+vbWJmCzwyv9LAml9s3vQ+O0ts/jsmsKla
Qoy5OoQnTHlrJF2IFoExl5V2FRLfBKMXnyC8nayr1ij3E3TkZcJ2+XShq+JTBtDJ
1kpNKD7XIBXGEGodX95JZfJzvmhV+VqrfjI2P+j+iL4HavbFTne84T25m6Ci1bD3
TofXn4fdUWGNgb2J7MN6A8pbAFIDR3LTZ+tiLb2HGv8Xm/4vsuyp6FUc2Y8y1whe
ubyHKf/AIimPdjHVhIooho8rbGolpXkfJG/sdJVPkSyt0LX5bFOfaqMz59kmZj3k
kgaBkZ4pjaQ+Hfu2/4HRUTqZFktfOOaaaRj7jF2HmWSvHXj+xSZQ/rdkuu51p+0T
ogtGj7u0iSKXFyoFrMOGW/375H5XBD5QZaHrYXRrAGKdirNikqR5pZ/ksTtV8g6p
2pfriHGPcbheo5ADaZcLoWqb14UXwjdfNoOvdoB9W2rfu9b8WqCy8trkkQMrtuh8
nEbxGWtsDYq9eWHWxwciRl8WNsLtYwHElWV1fVZjWXpB4+jv5gLuBSPksKtUbv5s
I4w/R8rN0bqsMqTOKotEL/yqoAA04jX5JAmapyce8hxtUJveXXm/tPzXomRgDJO0
UWmsi0/06O+W/dN/AV+Z5a2XaO4zH5HatR0bBBQu4BWA24X57FRWL51e3KYgBHt2
7mvpLmUdxRuTuRpI0ECqXbL/OAAWk2UYePNjENYPexH2NDk4fxRfjHS3W0+GQ57j
AguIwHkP/ncn1XeNWCOJ1jIMy/rBsQZZIBgDGdh+wb5UbkHFmke7158ghvdWclF4
bVnVkJGylsf/+snZYh0O7PrdQcx3iv1n6DOjGj0UKT6E5W9uACui5t9mv7MsZmb3
Cj0+cECRN4UMLs4QLakpdwb0B/OxakPDwK7LsTGbkMi2a5773XyQ42lyP1olwSuQ
M/gPcbHoCUZxDuvAcKY6enm1adYLiMrEAGzXOOFzHiV6ah8D6JzEt5dkWDDBP+61
xFn8PiiYz/Hm/aCAYzkaLXUTblmJybQH/z5DBKP/muJoJojKy3jh0ZPwaZ2VcVyV
rC9spxzq7Dx6+KaDNw9giyUfk56rX/AzrT7Jb9RAn321HhL9RiU4Hri7QFhvDqH1
F97GCTFl0yCLEwdauJTXoFJI10WPEoKhlT2luIFiWJzp/F7zyYYPkADopmK4mZi9
RiPO/xq1U2Dq0MdakgpSnWP7puURHiLqgl3onbtul/6ScYZWxl3875c5aRcRcXRc
+E0qlmkSWyniJRA+ayWCRi3uQ3XH0ACWmzIPmSpuR5ONgMIQj6sQXH6Tjya5DJ7S
rMUn+/Ha4rs6/RUjn1BiLfpcHFcdZMsQ6vnljtYgWOifYr9ODD5SuKmo5L749ZX2
xwRa7JNOdq13FgTEK4byq5094zGk6KVpgoKZuwx6Ypu5I9u5OumEh4Bjhn5QcVga
fxERlj/Pu/rkhZ0we79qvaH4oiuisU/6f3VFxjjWDWuwQVyxT5Odck6JCTr0cwd1
MHZMa6Cm+ygfc0AqVjEPU9RbaVFpfVawHjrSN5sC3kX0cc6cpF7ZWe0ZOH2AyLVB
wIHzjEQPXJox48riJiux9NIQ/B0mZqRoxY0POppOmG0kVGR3EFV5VeAc4a25Fd1y
3nP9ZiPUc9U1jbEUN0znvmBAxZiiTvJqh3y0VuYqNBYiBI5mOUnA61GJzTpZ5eGR
GhoTh26HsdBY1IJGm+dXuqpjunhzOYWaVAxEmxpVn+Xcl4BnG1MzEQBYbyaCJ8oZ
354BpY3NfPaWJ+gOof08n8zpECUIjsjKNNubbJvhDooyVzNyr+SiHfcDd1kK8K6Z
xelyP1fEH6iXG7+joJGw/WheYWEDNgBQHpgzCJSTkQkWCa0ZLTkGF3Dl1W69PdfN
lshpwA8fzeHQBY1tmd02l6y4lFbWTKYHs179NcppvTLa8FcYMkPFh3Wfn+fPcc9H
7kU7Kjb4UturdAWu/U023lOCebZIYxt7dIyFzV8w/GTq8jI3T3AZEypyrp4/TmMW
fUt3clcBM4zV0Hv8Y31XzcFLbIpE6v/kAyuJjpfnVD4kC3lUtCoyTLAEO6ElOvn5
orDi6u69sOKxTPQHr9TD0Y6wlHBRcaw8gAlNhV33+Uo/aXSjFkjJvaNzYBXa+6y7
LZE/zjLIXX/RqRUoZjsDLbmvatGX21AwhXhWA0QXvE/oA5BINWiuFXE/ZlJr8I5c
xMXn3x+UWtH+I1x/19lzqq8U8XtVBXFN5dOZfcA88W96nZNYz2jZS0hD/cqo8LwD
Xc+crS8BJY4y5CYg9g0GV+2uEr35+KfKoXxZVmyGaLYrC8CqvH1jLV17pfKVG97j
ek384IUgGbvsWxMj22iUuT0m6pebSCc/Ibzqn51I6E5zXIGNCcX2hCk4+QWs4bIP
rwxw18N7cQrLZijjPoHW8BZnK6GFC7m15+H0wngtT4GhbCfsArd8+RxWpy61rz8p
FPNtZJ+Z1wT7BJMe95eTh/68bx6RkFm3kd+uCF5qGR6Pd+E5R+NYMz4hcCwZpR31
WpsXJGR2lshdtPhrHcShWq8kZvsXCsodfrurH5Yfev4hAdr6f9+6D7rDx8wj3Klr
VhjRCXXcII7DylxCkmeMAgneQwEHhDnHz62INuXGBjKkJjljKAqtWk3+pn/KlTbY
ebyl57wUKPKoRfgnt1XIWRSOClSNglGpKVBDa/Gupqj3d4KpN97PeAYtmTktxECv
0kR3D9dp2XmL87veMOedCoIdeuTn898k20IwqPJJOvRQe7E4yZl0ikyvvhECM2jA
zNsGpI9xN1uf3bjfZTlXwNWZ0PY2owhwpRfJ1Hr/YtUPGN+7y/UE8DbDmMlN0zOF
Ls4rER2Shm1xgHLjROZx+bbX/f+McO7Q3ge8er8hgvTYWmYDR/wWd96n+HCHIoyd
xxAbVcaPrKmgOrgZ/dgOxglXjwsBj5czm+9m+8pD4wq0qQvjnaSF4Dwuedkkqpki
+EDQpm1yAFaLCkzNOeyUXKYVa/B2jb9vtPLyO5fSDOqO+8wlm3lF4lswGKRuI0mm
yWHgRHn99ItgvpSHmySoRZTALA3vH7RsbpgWCBt3zC2RLepDw0hjXAAKIfdsEK4e
FKBfxEyHD8/rcHbWLleidg0xBQ//08KVu5vRH1+Mqa0h5tk+jm+lyYoqwqFc6r3p
S7p7apu7VUpglo2KtNWAxXgzqopNRjSEUORiasL2uPPe0q8jnLp9yW8GdN2k6jaX
tNVCRE9YKeUcuziWiu6W4PrjEjoUbin2a1bCEW1T5Fide8xpjoA/ZodJdvG5ckU7
30S4uedPgvOKkwkAAsMIx3YVWes6W3UaHpWLVlNOX9vY1exevWGUPAmgd0178KPk
32O/9Vt+RRDi5mAwYK5RhHtwjD/tn2RMdGDik+3EeYnHr+7FaXNrYphXpgJeH33A
+pgadUt88Kev7GfvS4m8w0kzoqs+DQFhsVbS+SXSDr1x819rA5YzItlUNjvCEGMZ
l/FM7vWXwOvvRGEz/CgaTAarEvg3MznCeSdocL4fJJgcqmth/EHV/981QRfuV6xu
ryhH8S9hjuHWEvqKU1gWAwFzebhwJ8wXyOkzNPlzpVajsyCHBO8THTKvmjIeulMz
YDRMb4bfG5JuQv+p6oYd09uOe/v2Zw1ipql+n4CK5WzDtVN1FfZS2HGV9XS9ZCyQ
GlMDLWC48/Xp6lqcxnuMwjIcyVP/QXYlOanKQDs9Znj5o5kSFgN8ghHt/BMhruHK
Fj4/33nJyJhDksaW8CbICMsoM7f8rKFQMwa9iHvWaDe8/5RyC4gHBaKBJLsxNY2n
3QypbAmWmiP5Cj3U4UFQhgyv8TgUCLS4ykji1+RTahXauC9HAaVrK1MtYXNF+VFS
yrSO0hX3oFPQr3aB8SptzL5EGpYXPDAEqlCHqwBU1VTR9qdgbkJGGGM72nt5XRt7
qemDNeDppfg7+5MjArtj3Fq6E6alh/JTgWkzz1qxWRB50Zm15eiildeTJ/Jq19J3
jCWCG9XLKE9PfiKAGMxRF0eitOMAmbYY2V4R/FqwPHWeaJ8+3G7hgSKJ4nAiXpDd
gwA+2RrpTzYkro2A1De/lQD5JbAWgLwWW1BXnLYJPTSFJMC45UUfoHp+VYJtua7I
e2ibP3SEP1mC6rbjV2fsXsl9hrdR7JvdzJPUTvlhH9d5RIyGNYeY/Pl2Z05Pd2zz
GvRysAQNIMQIHsWuTl2w6djqdrT3qbGw1knmWjjzEfv8M3A8p9vIJBrageAhvrpy
s/uF9CQISJgCLx8TwRaclCcqhhmaknJIXnzvLDoU8/wjkOv9ALcMEtyOSoYjtEPV
4RmoC1/gTk3/YcVGZWAwP6do9lNHR210/QdUhlbqD/DobmTrFZZsrkjldbOa46S6
K66ec1XYu5/3rvdEcgkSRqCCx5/72KezI4m9kRpaGwdM2UeuFMqRGIIip6Ezh3XX
c7PSpkzEteAy/G1Bb45N5aEcS4o/9ObR/UXJJW6RoOIwB1RWfq0+OGeLAIhKf02t
Nbx8scyrz0PxZKEB0JENc3babvQIulFw52di2clwL3GquGz4hMae9yOAhL4bKIQw
ZNXmJ21IZZaHRQVSL0OOFd2X2QmQ59h9YrxFv6T8/Rw3uE/Zi6VVmbQhq83n0Tab
df7NI6rMzsfC0V4SgEdR95kms6p/zmEXucR6Hz5NaOdeE9CvFUpZBlJBB72q1FKJ
wXuDBEG1VXcy//F0Orq7p9i0UCC5gYSmV6TSoSizUdKf3TsmF7VE6K1Al2krdCcB
1SYvN8FM8kbxNLRVNoVJmri0sypFAsCXsDhlkYJy9JcZZK6qOK0uJd3+bNoajZQZ
o2eIE1FtiK+CaXh2AKjyWY7Ux4gswLaYvTVWDkAeHkGuAqWnfDjeiFIz7Gg9hXQs
8qZZDrbztpYWrwKuxMfn+aZcK6wh2xJxyMHVLU7cucYDQHeCN/3iCtyaazn84+/J
5wr9xV6l96EX465pJmNUB8Po4PjPHXRXezxNjEduurIcL6dLpRCnamTfXh6iq+PA
BWzXX1mna0tpdQP7yV8izAt7V9rZ9JIByfouDg0FctSHTv2SHPy+sS4pEP4l6zAi
EVfmAO/W/CHwNvdmXk4s0sEvAO+BoHgtP9NYE0Ap2iILUUp8xEZ80XDrjWFIxgbE
rwzOy5yF7V5jcK4e4lTmbWiy1EAbQtC3gi7Q6pLPD/RQYfApf+AFcYMZ9wVpx5vp
fqUFhAJAJhclXZtKK00kDb91y4E9X2s8WYk3yJPNLERXtriB3jGG0FCaa6727oPE
EnI10y8KUg+tnkY9LwgjTVNY8TRkVlKEHSFnF3ztOFSsdA8oJeV189AzAuwuL4wz
gD6qVcAt8vAe9imlGW2wRVt6XVFlGsolhmTW+SHqdIFTjBJbNt0fW2RiJQy86urR
8T8axsk617T/zednTkSwRg79AFp/125GGGGFVOi+MsIPEygWGnGqcGysBSE6nIUM
YYtyiAwGnUquQa01jpYG2lgebklfgUfR1r6adOjAAm3+2aCYZqBjmMLmjLQHIXEj
1Kph7N+aW/aPpn+SGEIfQHXCSn1hxz8jdFVKBO4wtEGW4qexykLsosn7sDQnpOZJ
ufZbdc1qy5IPHLzu8JhH4xG6AkDau2ddT8qRgiW78IK7GvJT2pKTG4jzRtrPbCfF
jpDnF7IpIDQ8eCjv+JFb5oXFckd85ZOi6mD5YIxwyaXer1KruPh40OUSEJ+tMlkT
FWXmC6HKSuf88bMFsLZJhDXXSLhKVN+LThhm5cPYCK+FsLZIFpEb1nM7u9EoPCjM
unz/6vJ+17lsovcESFMCNtlbndWQOlpyfmqisYjKVBHGf2t4OksFLucheWvoqZsp
1K/UaK/jvs123kHH5i3DuHx1rCrLSaXnw4piwLnewf9iDVcIAMhvv2tHGLURNUgw
esQkSunPdhGUEZNNuOq2xXgB9A2wkuDBaghtRP8ZjGXqGjHCMyZYkNm39fAuvxwn
pUCiOBqezriUwLHTkxf+3cWoJ75/oLXuOPBy+M15HlwS4HlcqAbtXZspQmU/8gFC
hHsFgbbx2HRajcdnFdVblECXy7AUG7mwYFrXEOx09YGMbTDm1wRqwAskC5i1WhrG
YzEbcUyI1+TeJhErwMeIpXUP6nMgKUGh++PQLG17av9YXVPinOgghkHvgFoGk/Bx
wIMJ51sRrlnviKgWneq4rC3fVIIFp3cYjr3ADmSDHnpmSmmFfnshmxnKARbBlMXM
vZKNn0T7+4B+onby8hyW0CSkEn1Kg+xBsAcrcOutEGGKNYcy+J/qGVA896B5BLqx
OOg7WoWdfCSewiXw9pfJhVHx6AfY7kNIMtswtzWTH7BI3KxX79UquO7JudpjZ6kD
+8LnfWT/ZfeSOAcQfNXqy5zEAo9uqeBcd/OxAGS0Q7j2VM80oqVUb+dVTiYORmoE
5fppkKzRVHK+biFiMAkgGIrYwUiT9FUDUZKbe7hIA4TNDR26vFtYWCToWOWF6nsD
1mQUnpORv07qWhG32lLxEtoBQtzHeN3FLdgLVpEz1dfqPwpUy+rGr5Ei+7PYjBh0
Y9COpVNKNfLEnBe1HsCOGL/NsQUooKhGfPCphYnlynXObPR9nIiPsJwtfB439Ldy
YFJuETfliQoh+C89KSNyu7kBZ9U9xM1jpezDjkmwgBv6cuwxpOYNp9KZADGLOSjD
NEVsQPG1BioorzTeVYBmnv+UDteCfmbDd757q52p6iegnsNk1Pp+ImR8LXwePez1
P4XxkHkU+0ojSWrqI/axiHTgDBtGiMMiqEf/yt6AC4SSqIQYxK+mIujcuz7j4eUd
3kLPQTGGYOB9yZlnqvSX0xjrCFONTxeVkY1dSjMJAspaufMaVNcbDqQ6pnWlI96I
oips3zc2Z3+VqScBF/cre5pJwpHVpwU9KHIkW7D3qPjXOd5kyyrq4tEJWs10q2tq
tOsRe3DM+g5BCj3cJ0zQ9YkV8WrpIQbSG5100Wyg9cY2BlbizxiUW7yyHxR8pyZR
8ocCZUZHwSOzGMPrYMgO0Z6P8blGofFnmnOxK0BEKMk6/mMUS7kd4OSekzoCrHsj
BjVLPZSgN0mWNw63TtrfD2cZTptGiJeknBW7sY+4IRJ14aFjuvtDyL86zreUOOmR
0eYL1xZnvP4Cg7Z+kqDum7NH+ChnF9KEyxZlQdRElPDs0PgUdDWHq6X4mCFNmfwb
XjplbGXBvZudIG98r0+6t7d/9OpP3vNMyWk702wuZq8bCCLxjq5dZNQp/CH7Ss+O
D0i3cKaJKQ+m6zWXLmejOuVteJtSlcIaWCtmF+szn1QmYANiLPYRbigSL+etdD5p
wy4PChOFfFkcCq/Jop/eh2MKi72C85n2USZDyoDek65FOlyzZadqq54FdMEINk7y
zG771lENYiolIex4XEbNXb9H1nhHIbo9rnrtEJFwDJrw0u8rbp+brpDsk78mOQzQ
EwWwxW9sQzCa1U8Kzpe7uoSdQT01FfgfU6NDmF8GDv0ywrjeueRwRV78iLFwJMqR
yveP43DOW2rmOKtlLhWEi8hZeEo9P3zfK527eQ+iBSKNZKpfkxWJgVnbzodKLXao
wWNTXb70375b95KcUbM8Oc+g8qCju0VFPf28aIVeafK6yfbVXwzyPIbHfxpaEc+l
z2v9ovyYRrEyYJr+D4pZMD3ZNrfTOv70Hbas5q7kQXPVUOXDFKEKvaVpp+ECfIfL
UxvscpLEIBZOOSQ0M/5zfd/tIbLJ8qf8jn6liDhRG3AJyxZ5JjZoNqGqkfRdKp1f
7kauErLKHnuaXqmaXskG0xQSipC7X7Wkx7/MhsHMwnCEw9GezSxWzu5rcVqBXBHq
BhAwwiYpIbfK1tRzPRj9VfPrT2k6kUSSFwAFygHR4iRzqo/knSERdR/VL23Rmatb
PVM60FLayue10xFwdap0kBBZ9hPDJEkMp5HVysB8Gixj0oRjqF5dXIQ0+fJf6g2p
CsyHOFIkk/BixtcRMLjaqmLCLEm8Ez0rCYmp7XC//YHRBKbvTg8idq8JLwgaIzS2
p+JJTIK9cMwxgMoEe10fAvTqPMcvewhDJZmZTDl7a+ymzPoLi/f8kIuk7ROyNMpd
1L1EDNkSfZdUUHlxI3/Z/etZGHNGmwP4xmrlRct6AwS5pPftFmcleKnQEsXa2vdF
bn04oTlX6FRKweXUS1UYJrFC36OlvG5J6cKCAcE+0p+2VtFy3qpQvqVXS8hoOMKc
IWazyviOOAky5+fe5zb1lhSY65iPSTO1oasuX1W6WZmZ8L7irjTru8A12ZxmoygI
edc1Uso0+PpWA8yrXJIqs3ei+Ah1eKVEHMgx2xKHxpcXRAh2XR8pOrmFBWzmP4tJ
FAMIIrNzQiX0yAwZayO3TNbaP5v9gvpMWn9lI50kJXhhSsTiFDsBJGwjHRP2E94s
BZ4r5FtWC4Ech5aVOLCNvLFzIrxjSALjQxqME3TXLtHgV9z0RTCFnGG98MXbWwy6
5jpnF/aw6eO0CbFTsoZAgm5+S3CTDimsvlK7mSMmpEUQreFJIbJqbPu9skeFXSv7
FLuhtL2+7osLc13SMrqyKCVfdiIW4tV2h2hYzuHXl99dAR2lThrB4FLpQAYeinzq
btJkixXnIRU8vT53JOWYZCb15Fd2Pvoz3QlGbvf1zNYYiBYpp+Kc7C2i6Sj8k0lJ
q0x9JLoK11XxuUsHKSFk9ZT5X8buMIZSHia/67DFJYt7OxtfHhAWmZa2w85q2jKe
56P7kpRyuskNL5KxPlPiTLjx6IlXIVrslwjC7it/7vctEzpKmlMASosKnslbhVE2
l5kG0uC32HOjxaPDUjWYW9/J+nedzgd0oYHznyDVOeyVtUBFgzSgTI2XTnZHiIDT
13+ErhmuvWfCj8MrFQV89azrqUImyeCzYq3U3Nn/NVGboM9R26AUuUwRCWboRTUG
AZqjeD472mS5UdtdN0anw505iAhxbtqR+Skk6c9v6AiuNNEm7qMc0WTTsqnMjudY
F2SMwRsbK2Iw7HkSLMclRLfDmXAUyKtB2YY7wTk/GisXpfX3M0WcaHZhzby/qCCS
jmTCeWlWDrk0U/FLjF76E/ywFw9wbxdze6RiI0t5n5WS2WArLHCItYOkKCkaGr2W
8Ye9ptqb8SsjFb/BzpRbKl3jOwfUh52z7AXtCDYMFImnLkbDqkaCPp7oeXcXo4y6
frcAhVNXPIa9SClQddvJSJGBRlCGKG0IOlPf/PrfcHZQz5/UP2IfAqtW58uxToLF
IsZ5vn4f4jDAT8XlXJUppL1P+ZURpK4z3DVLql60EMnAl0kA3S3Oa/CQ0uTHJKsr
FyJsAE8yRSuJKfCikzCdApX/5hoGsBAJ4xu/07RpYmDiZoyJ66c5iHb2K/FB1pYq
QVy8Cl4njHzFwwLL8pfXRCG/GlX0o4yyWdPMkvF+MIpwNl5br/MChJrRp1SaX6iT
TRPn8ho2Yrbhxgrsa2P0cDN6TdNk6vVH5lRDXcEcx46fWV9LbmgzVHp6lx2o7u6E
Y7h0Klk3/7Hzj5BdE2FNrxcYxKZy8qcUULQ7B7iq0wE7ns7LSU9HM9/6UYnIHp8t
cSBUucqZfSWVNj/QmgNA/7EMZKOBzL4v0NE95dSxwDW3Dq7yPdUveNWRSqm4TQ0O
/RnLzuI9A9UqbxQh1SDix0vz0yWrO5MGPGOXpLsOZrbb6k4+Fer8OTGTnOI303DO
kMrOcXpA5jUlCq3ipVNh4IeBmz/pS4ub2PbGoCz5vXldT+1+e7MUgN5WURy/IOxu
Hqevkj9TlRAt5BWBMBG1x0FkiGA8vquzcIOz3lW67T9Jro14liij88la5yHxyIpe
eqCAvgfqlJVIIhXRQVSVrwUb7NYyNp6gbxsYLGV9H3SiWle/Vk/71F3UarTC/cDc
iLUm6q8lFEVUuisTD2gFxvqyij9FfMFkxkAl5nha/YqnGn/hrCtIBJ+wghwKv0eb
2USPcfFH5TfLnE0fCajg6/LgiN9Q2O4KzHQY1x7ahAzbW1HgywJ/4Jk56U1dYCCF
mwrVWHi6Mlyec68WJkJ+7u0QpaNHESbopHa49CX3oyMERiE9CEfWtnKCUjzj42vV
hAl0bybQMFuYXA6w8obXMU6Ibo+UU88Kzh3wX0NB3YEEVvqSI4pt8OnOJRV37gqZ
9PF5mL4g59pONDAqP0viJa2MopSEksqTP/IVuzNAUNf9BZnVY/H43J7y1YcOCXux
OAL5YMbEuaW77virySzpiVt+RV2+14o7oDSIRA8fmDqI7ZxzYaZQc1UsMRq0vQw9
JdK2IiRxsjNEyNDgyDca0w246mNBqu9Y4O4/O6QqZWE9WWodWgQ+P1nPQYLTE33H
5cPfBA5v52QVnSe+lUcjtpuu8GXUazyEM6dLyZ4f+HYb4Vk0XXEVbyNkk7wuIQjP
kgMeRaK+xJ2kzS5xbg7sn8BlbjxdmPxFYmU9mhdCgBES+oAA7z1BiB53UoP2iE3b
OgOu2Qcz5jk1iTz0Fldqo5eQC6n1tLjpzgeoZdJpubOPWyzinoi58cVRUWp6xe/X
GifdCYQeVCarDFJCinFlCepjlqvh6gq6OT7MdXr24/ukwPtwKBSb1gEfHV2c7LAk
vyqklMdsTN5oK8jKgy12ppRziVskO1A6h8MM7E5hEecEoTvVP00xvXM3BmWC/1Uj
hRzRo4D5meAmkILxpIpx7L/jcGEs4MngixdDyDPfCdhxRdHMN3ohW9oYqqdtAwT/
zfG9K4nKlkyuRSp4oxL+lYkljHqBrqWUAiWzLhjN29xOBAepUTmjd+kqtXs1knr8
675Wv4Zoy93j0jfcFrPzdtHe/Jg+txzIS80Z2wRxaX3TzrzQkQI83TKdz/MZb/Vv
+w+3KutD5fP3ZqmKvZjRSfezV1KeT63MIqJ1h/ohlzNybrp6HLrrvN0/cvCbBnEJ
/r9D9NHEgAQMYeFWrrqCyEsjBmPeCja3jxeIRr8xIQzuSIZp9lbwYOWL4YqEb5gi
wYCWRsRs/WFhCmNhXv8SMeA99RlMcHInuGFnOp4WgvgjRwbIwYdWtbA9iMz5g2gJ
aon7h8h//SepF4J79FuD4zZvMX7QitbK1n9OnJT/kU8U7iqrYiuMIqhEbhJH4DXm
XCvnCsDzwdQXk7jcoy00RXTj083fL90URK8ZRF2FYLeb17dnrJcuNpQ/XdcpF0sU
Q8llG7KMK+hDcDU+Hxk8hCJa3v77Z2dr9/70+3/BL8uO815/NWPRr12jJL9ulNps
rsegz50c7GkFjBIOCKdBV6vbCws3XdlIWcM+eSzCeP2Hm79Pqm69dyDuFJcCbY9P
dJa+nF5SubTtb3tFSp3yOMrty1CPflRLGJb2z5c1qmHcN1trFUVpR5vu087gzk4D
5ZCh71EjdkMqMIbYl9eNX2Muv00lQgiHuNVlABFPmTiLS3dppDpJakLrGpcTqZO8
P1pxWFUWuehSci6G0ZqdcHr993AeRpefGtG06rSYNZXu+aq3xjOTvF5lXkbdb+m1
fnuBdUUzqSKlHsRySTRRzwifq/V213oTZWplC1lLmDMNCswY47dXKAQWyJSUVAxY
l/pehi68OCqzIexqY2y9SBBB6xWhwP7GCz/4ravMB+AP8l0rhpdWdpdAIeGpkRB0
YSaq97G4TMvhifW+BDAUwQEqsbPZOH4YHRxg8U4QTv0QVVCNOwjcvJm80yxsA4J8
1a7wS4rBqhEHeRqaQ9uQUvrOUw/BK/SLFYvrjv2MS5JjeYA7sjBPLrA8mz3o1wiJ
rVmZLU1HLr7ZkPcZFYUkCKI9Pzy0u5/axn6zR9U9zbEW480snbNBDNyNvFiCil07
180EQsVNvuE9CKmF6MYU94hHK+NCVZd7+PgXEeXBx+RVvRnQp7A3X9Wg6xvmNlff
8qQE+D/HZg78Vjn39POivKbwTIZZGrKcaF3/XAgIRqGHeBxqBzcy0kto9Xmgj+0R
PMPEDoZRLjy6Cya+kyfF+0EF+isb7NcNpF/HcIaikprZRxmkPcDvUfcdzW1nxEmE
kU2hDqq2WcqgylapK6z74K7LdeX6W/v+hPjPXt5t4z9z572c7epvucgM9ME6bEQY
X9wpom618LneQ5O3HwB8lzVurFPCfB0F0mXCaj7jibSYfRuvLpkao3KXa2kXwMBx
w6uT2z3nzCXx5S5Ez8brskDwNfl/dU455XuGvEGynGEBgGWfJx+ua6p6fKolSHr6
Q6OsOkP9cQmayXRQS0Xyd9oA/8JiG+Kgz9ZSgsBoNQC8FfiuliNaCRazwsTeHcbH
2Lm+FhCiGa6F37ZiyBqVtRzYET3dtld7txchBNGQcqF2WzWeY5QCGJHah5/kOHXB
p8ln5i8hS4UPTaen4KBFUyA5t6sBmkfAvCURQyjsF1vM8GfQUkzOPivOeOUiX5bc
WhJjyMp0pGfQs+Kb5DZpTky5328aiosLYfYIxcxYuHb6LyzojHa/BnbQ3rBEoL3O
Yc1FYBz1xNiAXYd+xKOrqjGSPZJm88fSkvwtKBaS0o8ux9JRVemBM5o7W+z1F+fI
3FRAbiEzwRT9NqiVnotSJ/t2IaLc8fzE/KXLpztuV0w7PP8OK+8cfhCmTMz9hxVv
VCCAlfq6bZhqNizgmt5gpEN+SWjJ5iEbVcRaMwdCfRxEpXOILIvVYgjAjQ8kYgbp
GbdiKM5cadS8j0jyP66Te0QPAu02DNZGIsOTaCcII9ajgnIihwVfvS9sM/HJ5fcW
m4cWyOyMFYSGwRIx1cw24ojuC+6fbPluHA73U9Ijxv9GSL76+JrLjLJVBs9hVqcY
xcXk2qGbq7v2DIWrQlMaVZnA8aATlXvkeuK9hzJ/tnsv9sIFpFil+cn2EfRcO2az
4pr3tEhzVWBmXZlcE4EjvVSA+mhk0bEa6LrUTIsEqQ6cZ4SJMO6WYzcsVLG2yt1/
TCdZh4UQS5Hk67BrLN0TZkXc+cdIMN319TRmTrAjOgPGUSjmQOVJ6DZu8+qEYFfv
SkC6LKsx3GMDb8lTEscnqkCksEOlCS97ZRm4xIspgFYVfJLSlJQvde7eiyenWha0
LBAcuonNlkWrC+zkGri693KtaCiMbv/Dtj41o+l2DAaTrI7t5nsgDY8nS9fw/9G0
K/MuoTR8cRn+YR+Y3w+gw6IYiTYLWa6H+wi1p5v8C9n7un01DLnpWri0+TDEwKLJ
m/gsimp7dEIWuVRs6A2YnT499876UHWa4JAylwIBzE4zX3oV0xyEOK7jgZ+UT7Ui
hlc3D4866AK0tnfCe+Eal7u4Z5BMBim7QAQHyID/wvTgU+bizjh2mnllmKppr0x+
NJU1fRdWU4DwY2mgFW3ESWpBZfKQ8QRPIO3nJM8N3xOleNMoscjRkc3UnRYjEFpP
1ogv3EwNsas/N/rSnWyHuycffGS7ygjNBHEvBKTBkWYICvRjXdc3/cgOZvuYJyWC
Z9a8HONGJ78UXYeFE1+CLA2/MWyFXdi1uMoC1jGyAP8dAkf9++soDH0HPokZ6CAB
+4Oy0dQocoLj1fbokVQXWRXtC/2ULmYQy5s96r7Gy7lIUaCNVSlUzb4UYGx9uboN
iVkduzLMDTJcki3feTxxCR6xC9Z/+QT4b+kk1IocIsBcIN01evD/70duG/WTX1Wd
Z8wjSTtqqZGZoiUYogbEnSUPEyi1xmj8ciyR46vPI4kEf4Ksthx6JvciEFonQ7mq
e9TvDFFuosoJ+9wE6/XwjZTO5H00iPiGXCfdo+NgfZDo1jktN7pPwk4U1U7odA5K
shM0OcOSc+ccwz8xJW4FvMAgOFnSxwFi7DFrVmfqymS9dRR8TfSQM8X02hfFVghB
UziTA3aJ6bJLvmy095DE++SxmrKgSATt44njafS4THcFGtIttArczUkjb/JejuWp
6pO+kh92JbJvscduKFb/Y2GzYTzSe2VReysCJFwABSx+1XA/hg2ShkT/RgWFMtBn
qQXW3LRyMdvtOfVO8mm3zld7Kd0CM9pQDT2rG72vDKodyyCo8x+A/6/JXBJsL08T
gNTu9Dk0nTqxBihwdqNjt1NUZxHSscbZ6+Xqb44S+4Jdom+wf2KedFJMNMWS2uy7
OWxthPlTeRe4AP6eHlVQ+BkJXNmhIrCWDrS2EDY2J1kO/TW7ZgE8tdkyPxpSQ2a1
9zTn/lcXUk+p+FsnndRyURYArS+31F7cX8TPiZJoGx4SDEtqL+VhAxA5AVaXMUP8
Xy2qtA8UatyTIxc++GJluvgr2K8HCx/Z6eNARAhpDC1H+zXmr8IC3/wVsBLAsBlv
51PL5709uKlmYBRyE5QcA8qDsTZmrHLysIdVfqDJd4tXwwjzRe24jkEq5YVGe/Na
lS43B5alEFqztz2iklEUKGx9l89inEnC7LWbBDzhuF0Pj1timG8GfyK4krf2x0mD
h2m1VQkp5i8eJsQpX4y71Uo/LvmQUBWlWYylTsbt/9qWlJdyWlr0QJsiirvKIZZd
I/n656n+gKyeqy2y+vGFFTmvk8Ph5JQwtxB86f0LPiH0YbOUFNeQm5DlfMZeDHQQ
NyG9shr7nb8latnmEq4z/eESzKBUwDiQ3tPKtAJXK+VhuL6YzOL7L69aa4E7sNVs
HiaOo77wU6+CI81SoXpZ84Vk2VNBuCR2fG5Qj0f9/ytnMKXBEf7rxJFZWNCVlHUF
S3o/41rb79sCC30AiPY/UGyrqtW4eCcOAhDDpybjPcubbsJYD3HMtHoGjTwZxDS/
VjctqfaxLlzabS6vkVGPHbVOEZeldqgix2lW+YLGCQhMclRQVlhZ8Innllj5Po1e
dhBjfxNZd3L16qHc1//Q5cZN/G+50YYMLJiiMnL3ckUb+CLcvSgJNZoRQTtbw/C4
7z1GEOMD/rZmA29SkQEj2sZBailAIt8rd1G2SfSWI7RgI354LBIOIdDAcpjOlECQ
w06ahGBwsaVvAgvPa8/sSITR5nUefRtX8iCH9RdJChT7Gzu3rzANDZbOyI0MHa12
AjkaZVv5d9YzMCxpTs4KRL/7T9shmoF60PMkvsmSxYwIR2Mrv9m3CpqEPPFMZDi7
YJe9U7wvRIj9XLPp5rc+eT8xp9Z2p9jlt3X/v5TNSR6VzuTBgk0RBuQq+krY3cjx
eCIPvRr3wUx7FqC0ha6k8GcvJ2qR3UPAYCIUN4XubQtXOPZIU6wqDNcU0myF9ZmF
xipZxKq0VNg+Fqvknhz6cr7cg1sJkS0Gjk4KPjVko4eEtomgx0ShFqcmsRKwzFn8
LzOiQwcDfx5xJU6D7RoHJpOCaEVfVgZWr8hRSyihVJPZ7RSOZFsQ7UUyjIrYYg7z
nBFq+H+xpZJGjFFeBFYuLwxgmWzCB1X+zB6waeIJV8KjHrW/ThVqoMI2VnICfv7z
P6zfTfAM4WVyldXDzJHKwUsw/P4lUXeZwF+gebXO/ERMaOVzdS+fDDa6/E87JUPu
7fPTZ4xvLWI3GRCLUqfjJRmpXpv2UI3KL41ri/txq8dx8OcQ/1L0/q2XIjS86Wti
hPyyicAJjxDX0l3WU9cNEg4hMZRwBieaYZ9IrP0MYkmNT8G7SeID/QFUcQ2UTJqD
8uuzXb+yU8VwlWxj5ZQd+tkM4xMlmGW8ixKS+MDgKYXoxCWCVAcHMFhxyC8Z3xE+
yvmOwkGm4cEdo9qda/5rA3obncFYzQMg/O2wQS95aNZag+sEDwgDO6xWU/A8KdXz
Gy6rOX89IyW3AKzq0/mXMtHFt8sey53t2GlUhfqcblo6dWUNnA3cPHY+31u+FOAQ
cA5u5dY3vWyy03hJ4n/Zx3T+cg+rP5/A+xCK34BJEoc7m1L4tDjMSzhWdBvkzh8t
O0J90SVA0WLclmDScTwc0JgVBtPJGCCVFLa9TCWTMVwv+jYtfKHkNEPP5Z8UbjKt
oJTTCVpYNKO1rfZ2PuOzmh6jzgrHdzCbVlpK7ht6zpLcbBSJS8N15x/TwEUb/1Ix
bo1Lqj5VLDtnB1CwTQRLAFWOR7y9wUmpCumVBbaoKd/0i9cqNelwLOGQjNnzT+4V
e3zJlgTMzu7m6jhVUJa/rPj9v3VhOjoNtF29MJZxSVQROa0aO0zUbtzY+1S0OA3i
+bk8O65FaYhtKv14513Wbdbe+NLAColMoSHnp/vUtaq8EtZX/5TDEIZz1+1wuz8Y
uiBbI/5p/ka8LABk59ndtIWlb+6KWpzGDGlbrxGP0RrzRxR40KHtt9kHRljJahbs
HJgsD7arOpVapz9JvPxPKDk1UytCbvm0v4z7Gts2a3mzZQG6qM3H9hUdfIpvKbcd
A1BN5bBRZkNzj/atWe3n/QeoTrDouNNujOqzbSeNl2IrrAff22hMWGD71+8R9h8M
6yVkjtJ3qljfGvYIldVZ97cakZq+E8+WHcW/T3HATvXBGw6x1lLr2D0pz+CPthWd
sC8YG1MoMSHUFZqEN/0c88PkUXlgADfdryR+N5jsJlxSh4CJKFm5k5+F02tANqeI
0uP8ZH0/ShVdYAVewdgLyRiHnokJxHuHGMhIpzDHK2q6OsyhpAGWkbJo0c8uM1Vh
iRAAzD9CEqXpLbUtSfntpa7p36U9/Pqssl4ZkOr0RbY4/wwHVTRz+Wsy6TgwqCrn
X2F2679VrmgEZZqLCA0eBvus2kWPZTk34849L/R8+iMrxKdJ20vaVTKbdPwd2JU7
aCyDSEU3FrK2DZZ4tRCq+EsrIGtykcWIXN3M3JOKG7Y/IQIKqnxqGzhj6G3t53lW
hgDgS2K8jY2bcwg3RprmkQPcjWFwGmfz1YSf/9wnJvYVUYvcERA8iHlg6Rm1E8dC
96O0gEYNfCRm6NzPiPmVI+XOzzChvQwayatGZKtKHlQOifIyVHVBnhv6ULvJ3kgc
q0ll7EhipXow+azM1DWobNLd/wXxnEw/PlcXsxv9GO1V42/1+/NaiBSfHc+pKfwZ
Aq4TThjSusG/sH351Lwdd191XEJ84teIKj+mxPRsw7s5ki016+LCLVtun+ykT5Jf
gTh5h7KkDup0n/eKFSMIO15N/xY1m25UwFMuyhhaB0n5sAYwMO7GTrZX1eyOs9hN
y0/LsUlOkticmfv05M6d3Q52s4Ayn2MkJvJI4n0g7k0JlK3V5Ma5vx3pma4SfAqF
I2W8gQuhJYP/lhR4SW5mr2AfHoVlGYXFeBYSQztP6RBYDoFsMJPSFd7qeSswihRm
J8fO1RP19cmv/qT6Be00NfgSD7pNhCBBDvfPtqca/mbCqsq5j2XJ4vryFV44sRlB
U4nzhlnD4IVRrLlHvh3nw9N+Jsc001J8yMilDyGlFACCFKRze/qrnmBZVVeXieDj
hGo42BUL/Z/IBOU6llUeX9fETWrBQeIjHq//YjHYUnCROhS2Etu3tf21dWH9DIeK
SadJZ9AOOAE9q+lXc4lFYoxYlOzTPBw67tnucRPXcBusQ2W9I2hLLvgjG6A2z6Zw
ps+zSHHglvpfJZe4rY5GIVRm8aMO1KB+2xqO6/jpYTcS6AoziXkNLtnK7IAMU/gN
jOtQ2mDqLWxH910jwPrqXDgGXHy3PLvHJx6tJG5IaDhBC+A0ZFyWmUXug45arorw
zsuX5KgewA2Qw6drllADsBfjankx/8TbCb1/sHQAI5XWFzjrIHeNutEGzvT1TsoU
iKhgz9VSoBaKx/OFcy4JdpTkWbBXUHzUSHOU8b5s+H1bP9+nKdwptLHFKO3V9YS1
3N8L0+PVQssMVNjJkU8o7MWdliJY5epxXm2HIytulm9zX5cms5Kd2964U8Hnsrrs
Dlr0yWucxFiU8ogjVkHyp/RpzL4/6bmQDNtPnZeAanRgVpfEUZFl9uWGyhBhVE21
PE0WuSu0SmFKVMjObkzjo8MP4uiULNUnxb++q+PQX5Mz37dyn4/ebUD+2LTEW2jC
S7k7JWrz4zz+p8m5H8RC/7974swS/S+0u1GJbznyNRF1UUVNUnlV8JAjyb4zriKe
IA7Ih7LVXZ2LsxN+hfLN3rQzyRzB/+gDZU6WjLYLeO5iLYVncjoH12PH+rTdxB91
4KhHikbXx7VSP7BrrAF1xXt/O6aIQoIdA1xPLt/Q0M+0ow1lhXP4TaPDwrBf4isB
9+0K63Ca/IAizUjezn86efmKaObkacUX61fr2mZG0h4HhdNoUBukCS2g8eGhLa5y
XvMsJohTF+QfhhYBjrv/JPqRnoEB7u2gE/wWhriG9DuCsGmVbVZi8oga9XzHCKpD
uNOXat/cuvBNa1Btq2aYkNdzTs2mlffRlhGGE2tkJepZHoHibPETHWTdJ95iUpz3
0xFo352LKio/xJUMMlUIrtYYrCRTEEvQ4GQb8tGo/d4hd2ICKn0DTKrnLdUUlZRe
TsLgbneSx7ckGP8ze/F+RbuObq90uaWBW9Iym4rn3vvMqhbVFhODcSxPSJaKOtrq
S4S3MMToTpJwQTqt5nSS84TSBavr92VOPWotpRAg8OYGK9HlTj06aczztW9cXrS3
C3eEizhm86Evym0cyEpOFrmthWE5d6rfWE5KQhcJfM7MrO0fKck1nUKlmbSCecAX
cpo6ylbnsDzxwsQqeBqPXsGQxWPzqrqfx9UPL707mGu+gvXsJcMPi4Flu6TGosIN
wFfjVUKhFCvE4D2UrY0u0t+277daBkW/lDKR/YoXWEpOQ7yTPddcsjqvzcPFbRQK
/MeCCt/LSAWRaqOYTk2tCYVufUp20GSifc6T5SuaNosNBi2ttOa8igZNJMuv2b4Y
RLsgpQaFQVKQuNYLHHCtqvEBFpECL3C+RW4leCVfyUo3HQN648g/ac6azEV+DF37
yNjdAzuDocMaJb75kaIepgZyRO3yW2g/XnC1MAM0U4c4oJ7CS3lh2HDv6oIATnkD
y6ADD/B3Yq7sIvMEA9uD6s0RSs+e/ZYuvW5hLG6Ud+7Sv3kZeVG4MvVmrOZgwuxZ
DxDsBdKgXco4w3JEeFoVLXjvmcDBOmGtXcW4X9cU+R1BhqNjlDOrSLXo+AuAEom0
DE9cOSI1evtPv4x50U7fDFsl+CKQt68Lof/dh/hoi9j6lF+oQQ2C1xLTRSHyO+8Z
kqh1cAeE/2UdBi/RoOFG7qrKA2FijFWJ71B+q6Yh9RVZAlmMwXOgHfx37CC1yqK9
upNMHi2dr8jYuj+R478rXj2UZw/wZ4f0kEGp3ZACzMnVCbTutdAZmSz+0bjUoFtf
nVs0UohDeHIgH++IXKepf9vac9CSAj3DYqcwuM9dyyb9d43TjH2bieVgu0sTFjv/
jLuwKo6VK0yeZQtfgJRNt+xN2p0RkHbSqnQZ7N7tCPq27GF1C+xB8g2iw4bvuX/k
piTnpPzX3wvsZS9/nBYqrWSVADopuuXjNevH63gINxFpPElvVjCAioTT7Z/MlkfF
4wopIMSgMkGpkWGEjpOGneJsgbe36+Ehv2yCO7frPQ/E3rdiod/JBLhmCj7VoAi0
kJ0vU9qe/aJag1rfMPsjWQiAuTcNsTIbAtRTEemB4OGTK/6hVgcD0U08useMYX6/
K/gxPOfz8Dhp3L+S6j2xBnBevz+S5KaGaGob+lSRJBnb4evotIqoduYe4egdGoKI
1RFUAkMoTZWVwGF1AlrrDwwxU33e/WoUQUtys3iEzN1/jLR7v6c4JKZh7cdv5RcR
JwAGeY7jjj6AXgbO0VuZJ0lZNwqxokZLsFlEGY6l/ttokENaIzXeo700NqZrJIKI
YHaQYHwImAc9RuQaO4M1MMjmTD2h3ipSC5xEb7PaF+Ba/YjCL1BCrJiOHwTUZgHO
IyYM0G6wh3j04/XEnuqix4dGAA8tdbgGwrKcYFkcPq3IUpWM+HYz5DkKXGxAeW62
dzRENYxCKAVSCqhoHnkt+YujVJwRgwRJMtfeC83PB6ME60coSkzvGkOic1V0dEy7
XvA1JKxZ/y7R+IgRcsY9YBs0aW4UQAbw3z6mt5TKDuT9XIQkZEsQyiPrzQfLIpqR
4SkUJEfLLHz9FT6dkJktckJewWSMeyXYxqdFac4eoR7gy3xrlerMSUmfjNHIrP9K
FZG+a7Q/x0WuWzO4Zf1cz3/VL8+a8fmZnbYQhRwZj4F3rHBSwJA1/nCdhuG/QvAR
a0BO85+6OO9qKhJjFRVJhbNd1jwvrXYhHWO000wc8QVELDZxhnJKIl3+IjUiXYEg
tr33G/1Oj0GFGDV2ClqJzpqySS9+GB4Gew8LlrBNu8quyOoSFvvV3uNIj9+cAsGO
pS0Z63EnAzJo+HAFEDF2CjtD+jjX2RaucbsMz94uyeLALjqa1W+c7RVfvwiUbxJ/
2QEEFtFuFMUZCOMaxcUxO7oNQGvJBH1ZK4+X41J8DmMA7rt6If+PS7sxVQdrNwdS
dq5JHrHgT+EMKBvlC/3s8wukMp3+CSCPBY2e7g8Wv+2cgIb74DRRrxkegsvCJTQo
gfP2B90zBC8+693BJpT3winWy5ZkaAYdq79GRD3nJ5ugTXMCiqBYiv4xp1AHaHm8
ti+pbBJ9SACfIc+Nez8IpUhIRt8IrdSM3rUDqMOjHorWMebSLETqdtYekYo0oS0X
8FpYKlEA7BzIhy/YJW1+O6vpI2lsYNOGrUDPAg3TMsDEUWOjKPaoZ6sf8Sl3zR4C
NDzJ6Ys5Jww+6BXkE+yAdBgfbu5JDlHJp0V2X3Dx7GtDNPwsHikO8vJOT7xpA/eY
5UAetk752zbwYmoJRdJAWoCg+Ssa0Xf9AAlIuF/4v6C28ji2cBr5M8k9VB0a+HAs
05WTSRtS66rtesRWnfTUHF0VCwROFucK8mfFW+qiGFQUCCM5PNDaadgbPiVMcQbk
RDpq+f2dATdlKRGrBwwKoABMXwSNu9/Jvg05iF5NLIFWHgeLD24cnx9VViqQhg7m
TJOoSZP0LxcikybtGrgYnkytaX631zNevVmDhrlm08kCQVk6lWOWr6w7FYuWuyNr
ChO09Mu0/+nnsvjn9plYa5pB4OgfKzVh6oF3YZ0bTts3v2Fm+mzX9y39Oe7p4Uwj
D+mtpqtDhd1lMGGbUtPUzA+y5RL4MdzG3wm/O3pmx4XU24b5dfM0GLK48Tg5tovH
ep74cBRmNom0B9HC5DjcckMEqr8QjfUscAyzc1GOAmFQpO6iOVEdUdVtacioCIt0
KnSueFEiRqae1uH8F8NVo45nvIu2WFTJ7UVTA6Avxhk6wVatH4t9PLZ1EGyUNC8z
ZSimIvzEXaDJHMpQcrXNKzlgnGLsEteveRnWb/Q5dFLq0OV+d/6e1aeXLgJQbUAU
/9MyJ91RWwv7yf4yUyXMg7Iok9FZhs3Yuhxq+YxutyYYS54rr9shvlwoKqoRznrK
fPOSIdRhZbff8dvDKDANGN83eaIkomsQWqvaot9amJewyWK1zENWpWeheQoJf9Td
I69FdyHKdblz56tQV+NaUY9cwOuMcSdagWtIwE+bGNB52s5oZLPy+iNxRwFj/x+2
7ztGAPmtgpQbl8EMHtkrwul5Fr2vc80GlrabigoItauzsaRtC+MwU5eOu8DF8Voc
i2A4obwdb7oBT6qCJNqiwiTb2jFJEGaTIgh/VzZniXo4RD8yX0kCEfUmjVAhG036
/heN3e7exXvAeqNdrogEbwwzp9OZLr+2ZCR3NLaVEFPylIGKOvgyLwvQ7KkSDMZ1
z8XjVaOFqqB1v1W7SkzSiUVtFV3hZMVjCyye2mCL57Vt20olFGyyLbwox8U1xll8
nIUt6GOVE9n+z7lsdCKYpJUAfhihs43QRlqVSA2fiO1x2YzgAvSyFuEY5eeQDOJW
i5R+UBIw7nYh+EpJuOf74vJ0LEMscekMZjGfBdyHrZwAIdoGEGhkGYtOez/bYYiY
hIE4DlVkvuP2UY9GHCORb3iwA4UPIVggR8EP0ebIP21A+JSsEWkPN9QUuxt1S2ob
phUjS+8JwwyKcyHDHq/LiRGBqASmPG54OatYSQG/oVB8384uHf/fnENoZcdMZ9fT
e6zZOn4YpqGaAZqcwTeT5XjGW9JRS60Ll9jwUseQ4dxe3Tin88zCc84LFJn6Qmmj
Ma21F0nCsZ1Vf7wlAPs6LsFuOp1KCkMpgu5WfHELa72PkC6wWjPRkJfpPEon+wd3
wvGa2X3PF+0w5T5cWK6CkSXYq1iQzpRP7no132//Uc5Z4chdPRsUtOPfM31VDM+B
/Sp+u3Rdj64j04h50wk2w8XBvSDwKa1V7XQrZfR+LfR2rc2iWlqWPnkbxvjkMm13
2r6M/5RUREE9R+hJ2YzMqsSX6W34BN4R+fziemhZqS42BEV8T0pOBrJF0wHz66iH
zP5WnZV8emPAepnq/c3sS7exo6WJ4mJMe77/e9HOiL7YgnZg7EUhKUHbt9OnbRQh
pynWzs/joZ/Gurk+IxhhBLVbt+fz9lRe6cVCK5hYi5b2wYeBJSjApuRlyny1hW9E
HfATzhaAuqBcy7T+qKOFbxP3uoIsqb8DRm9aSuJb343PQg8zr0KCrf9eYgncFHxJ
KZkvd2ubIlhx2CpvsoIb+E80s+mwEVTlkg7aZwMKPOSIE3IXpRQ7lIL/Zd8j/mAl
YS0t10XwMrM5Z1N0DCvKGWKQL4LJA4ct8HBwIvoHCI2psblCkmmbPEbDzKKzzL95
p60n01SjrHxA5/CQJILW3yYIY5quW3VNUZHESOZta/Jidv/mOr505l8SlIExGh+F
2Gw7x+U7WuD0WMdtHYn5oOHOV3Q2/o3MQ2Glyi5pV9JcvYuU9bskpfJsWAyrFnsv
eSJdI0s26D9aL+UrJXZ15+BxW4jo+qpe8r1Qt5lg8Oj341dPzLeF5nAHYJ0Jr3Jg
mEF7dAEhmV1fhTCTRiZntrbf1tLkScwNWdvqsUH9w6SVmMYeHj/HgWCKjMau3KQg
WdXpvhy3ts6wRmvu7/jADHSwN8fb1F7eCkEqOg6uCx9dmpKvtzjBv4BAFtK7wL7C
6K6ko7+Js14qQ3vONzpwbMVHItrtAFlrERY3wkaAmPK14WRAJ5qH5LNyXCZdlNzz
RvPuqlqoc0DnFiHy3vGV9iBzxqRbkdp5NSSnMjMf9WeqaVvR84jc+ctyg3bAfo8C
abCEx5Dds23PhY2XeJXRZ6BYJq55PAA/iG/Iy3/rQ6FzMtdyaZ01NmcRLAgu+BQx
DnK5TFuvyeV3SEaQxo84mVvIRWZBrSMDasoAQ08b9lCMQ1FebgkQBRyDDrg1y++p
F+uoVn3o7dixBGYvulHg5iL6zF9g8MvV3NmcRZiwphrC6Nmh1yyVWkKZElWGJt9r
XwxOAd9hJ7jIzGqSNyg9WAruj0Hh7Q7Of3rayAgLrqnBwna4UCUZUuO9sWWcMVfI
KViu5EIGGH+dQtjhbb1CmyUn4sMraakc+vOI3z+YUJ5owo2nnAT4lfNjBwRFPzOF
/fwoJ4gITMdRqTTY11Thodx9LzOH9b7H+I1t84KF92bPnB6QvHNzU5NB2kY4k52c
ojxffwpoAhUcuI8ZXXR58KWfDSUyYsLyeNSDrUG7oa65USuddkBZcY0b/o5TVwnz
sqcg4Jut8ms90HXCFGSxYJNZp/FsKFgxIvJ484823BR2rCBjs/1HJ6BEzMdhz9na
HdPUP+Z4mkPEovEGTWmnhrK7/w807jseijSU0jFAIkLRssnM/LQBvESlHVhnVwxk
AdrbymzycfiGna7wA4uS1CTEi9KGHFb8ArdMqgr+9iLmk7FzUVXP6ORBo6JQ1hn2
38vyntUoMN5lyRs5B811PaQz6nFO3MbuVoA0pMdJRPTUZ6p7pCzNki1N63znOymn
kH7/S8K/F39PnL2/xXlivcCcSeCnBOElTzVdW/Yc4iQ3WCVS5wGq9Hf3sbfmCe8I
xdIB2TYyOadJBWiTTcyc2gRty51VdXyFpGGU6Qvi3my458yutmno9qz6WP/R6LZI
NWPLzYD4Fj5Odh93yhPoVxTfAj2+90Ch3SacYMG7O9LMbx3QXyQ8CLcvFtNQseeJ
BmOf2LmM5gG9btQ7p4chrSnbQ4OlSoAE8G/lklyWq2drxbwXYp7rqCv4cD3Ug6x6
pCAxJM0xkaRLA7Iy9QY1Ytyhb5f/uQneoqEEdIsd/7dU2BJOXGQYYaQgu6F9YbHJ
CZiXhlr14t6ogGV1hYzkg9MNNFiZsB3FR+dWSkPQWvKHj300ONANyBKSWb6TML/L
GkZ09KfVEROm4uxO7iSqiKVgoviUyQyLwqJPMqExFwo4cmYYjEcyYK2Hz/C9vEGK
l3bMf0rI1BcdSddyegh3+/aPpEqzfrWirJ1uST1gcdvWzZBHGXWwWCCMbh8DTVBP
wyUreNPHqdEI/M4ujMmTfCQVFkjuK9MyTCuiN3YDtnp11v73r0iroyiohAnc3dMV
ZvJfb8EmdZXcrgwm6PiBTN0k079UFWpWUQtmJuQauH+Ysnxnlo3IrwAPu5OTVS86
nScAGu4inxPwxRFD1jxO5Hsah2nBInXnC1JDdYvhxOoYL5qROqkoiLS1xKuP8Uh9
OHG3byTRA7sE4N/jOGDwYkT4GtyMHjGsscgwrfDF890mgGPMDBAuqcTJV3r6YiFE
9UM21nPJA4A0f/DN+EHhWSlJ/q1MMtLr7MhWHNRdaJZumb903L7TBx5G1frkAxqF
9mxeugLbIprks/wp+VA7uQ1yj2x2BD1XaarrPwjRQMh8VD8J3mnlOaAks3sMbxoy
Kr0NdBjRYWf91dHqre6DHXL5bd3XWKWgBzDg47MlS93V6Rdyx35/tIgctqlzhdTo
bo/zhsmLsF4zgD5Y6+60s3IbH4gylS37TYbF2Q+cr1NVGwoZfz+Hff1edB2Rsqm3
VW5pnMQib7bpavjkkMUiRL6dGXmd1X/aHl3LD3L8+DPzFTDApxiEh7VAYwskQ/U1
mD57VDIYlt13zeH5ax7ZXuN3+CUpv6yUv3Q8Z+ktOIvHHZ+vl8w/RNPYOB84DRvk
MpBztH6WoupauJjSHkCEBKpuyICtssgKVSIu1Sszg/2+TlabrfF6J2QEpeRuN3Kn
HKUVQOEWW6Dg3niBEC6BSVAIPGPBkccVEt++q+8f/r7o+Fr4nbjJiIePgNP/uw7j
GfjFbuRbMKr35I1js0a7wL65+oIxbSYcEJifgQCvEVSAv/SOXR8ELFSIEEYgXcYW
0O0NFa0gNptiIO4qsJwRuMfE7TW6dEki6IYdYx6TtawdNGcNiKrlTL/k1/pR/rXj
tQKXzOVKrwAmWLqy1ycxwu1NqR/6waqAUBpNZE5hQhRJPm8QpqCkWOXxRH/jClzF
sx65GjzOqbO8wTgccAexC28BZajUVfSzQ4d98uOhQp0vh0MXRGJxFE3JXKs5GlFK
2KswYQY1VFdlzEKoQSud6uDxSIaPGrhB5jBUOxR8dTQwkQ+FUyLXIOjkYK5Y+w/C
ZQlUIrE8g0BvVrx0cEGBN3Ldbwx90GdVKBzLrThjrEnLGtTbqvYMSxH+DmgApQy7
FjROFpMQ77wgycDLTaim4iM6ZBSGGEZKmrpQRS+O5Q7yxsPxxjtZf2KgC8v6eTfp
OxkZXPEUFKalUMCwTwn7MxWi8p8buYdEJWLZQw3sPlrk7yYXxdIFVEP/QARXdjny
jzG8Rq3Bm1XDXRVfO20B7Nui2lfk2tFQYwrSm8IO5xamNr+EzFOM6bFVST9K/zfE
IJWn62Hzc3//XJIAHvOz8zDIe+s6Ar3/omcGk6tdSfrdYOzODHAubl2intgKXeVy
D7GSmikdpFVEmUTfUP9KxokXu2rkoKZzT99jblNDvzsaxheO01GfAmWP0UnM9+MH
thtLIXEG7LA6LEhcRjfhwpwu79NyqjThg+lMoYbRemaE+J2R6oXdpQY8X7M3q6TI
GJ8O7DbovE8CH91IrATcNGm7II6oreJKk+Yz6gX15XZ/6MAAyLTjnDgZHMA77oSl
a2nrHcKy8Jwq3UmIDmjVtWz1t/7mVVmc0202cmQobl2qSD0xsXAxSH35mxQOmnbW
vEayY3jR3VX+19Qqv5+oRdw8VlI2/p6Odu/vmUByz8xJdg5b9nOJ+GW16iXPZxGL
jx5fmVbtD5ftBaSWPH+DYWlXJ0WVehay0nZw9dCfdxBlR8+KWcm6OgoY6L90mAIK
QLYLZeROeWv7UvV8ngZmBa4SM3ai8Y0lQk7BHrELYVmKW3TKzt/wdgsQw7mD7YMb
f6KQnbH8z1dh/KFOFB2Tnk/G6wrYX3c5+gKjDzmYcFhe3lt0W6O4MISww9yT9WlS
HpXZS5UDTfKI4l4GNeRYNV1aG3NicqledHapfqO316CRdqLOT69F4xN6j+BFp4C1
bL1x6ANA9xD3eq31dcnUA2Jul24Ax5Cadj8lgsQFZ/hRosPAykv+CVuPJXRGOHan
5XRFGzmx5Tv5YHjodV/EyBGkxuQCcDWMlBUbbqyujmFX/kdYiX7auOT+BdGlu4rW
ei1v/FK7WASY8yn/Zt0lv0S7vGAizgp9qZlp6GxoPi58ly2xbfZVuISNesUI2cGr
Up5UeIO84+Rx1impI0AI87qK8lMXHkx7y5YCrNMpWvs7221kdo9x/DUrpylD+WXK
ltOAJ+m5bS7D9ZOA1hbJJiGjOIX/pbeonR2Y4mX0Be8Po1xYGo13tGmFGBXBbu9c
GTH1oVJIAszk74kyL0ZisCmOq5Gj2MAzRMy5uEvumvEXNABGPYANHH5bkG9vQKUE
teyqDKtcQw3ymWM2rraLA9iz9VEciKmlf+E+nLNwXHNm8dCx9xQKsymbYKCiOZdk
g2r0qDpC5zZ8Qw2F1HvV026hxG0Is0MPLDdCUzeRHqagM8ETCWihzVxXXD7/L8Kz
9rNOUGISJ1sJtswU201oRIWrlno0hbZ2HzUuwZfZsmnB6+VqDjVjZhvDl3Ci/1jp
6T2rDt7npMEInq3OOoANoD5XC0GsnVQYgoMGupAme8QkFgG0mCOk8V6GFImBQSde
bYreqxhoUcSIaLpd4QpyBZ4TqfkiqXsP5GHHuhWN2jduzvSa16/PgN3FdvMrzgdT
o+BsdPacsSAOoBOKuzwFubzgpVChUGECzOVsZjL0BN8CY0F282Xywyw4TahPLG3k
Q7m4n5MR0iEc3RlMl9Y1bUINQ78mwV0SrOwuUSxPf+ZLDkW9z4EBpEVHm8x2uE6Y
ebD532/ZM92hiOHULEd69Vjf5aMBrnl02S+/+l2EqvkinnUrrIEaCl6RziW9uuas
3J0MM4G/81EZM1z32aJiK+6EQbrkCK2EabJvYkK9KEkfoa9BtYfhPJPlc3c/CTeb
dTmSgtr5XwlrLWj+W7RGcaYcabxL3Jc3wRe3c8Pfv5MCAjddaYXJ1u5o6I8prIP6
PpAkqNnT+UYBeVMfvdU3Tmh4xPv+QXfvGDIpADxihVQhUpmL0isJCaX20doirgy/
yU/IZf7d6L3MK1qrW7P+DNY/IFjrxRa4n7pB9XqRDLblDjga/c0BPmefO2kZitOB
vrDDVCEw5932podnqKttCfavtnQvJOVFwv8K9GrV0soOV7zhIYcWIycTwu66yoG4
Cr/YzbB3P+netf2xGyp24/UupwLTIWskMM5si2llXdX15Jvq6NACRB+mIFwob83w
gEPxmD6a0UdgMY9TFfAKh0aK5feNelsfQKQdBNg/KLiWJLwIBn4EjQ45kBr8Yqn3
z9rQc4cjZ6K2vsdbBRnTIRD/0cxdIt8cxEdsGjvn48UR9qJLog+rE/gjgSu3PHsd
By1mYBrekUbdTWzvN9hTK8iqJmnNXNrWgMOtyrPybmw9GWqtWzltKyZd9RcrXpH+
Kgda8hwQ80yo1NVM8S4WRyHozFIiaoiy5ldRvMqXbLFAGe14Gczyr35ml6j+gtCN
SBQsaUVr/NCp05JT6eYXkg9BOGXzmKCxbqi3GIj+smdqJlFcxpCOmrcLJtgabasQ
qU6Kkti+xroRDdaI54hULXPt51doF70aKmuDov+e51MVgBU8kjbj97Gvl4C2E7KC
G99WHaxDiGH5YbnNaUvvTt6pDbuaOdRa817V7PpgVNd8bwjpbhVMN9pgTqeD69go
rvGrVg6Vw3Ro43rOzuVHTr09woBURe/6S1FDzMIYHsutvv73gIsZD3mWJUf/aO59
qtmjomGIiqjYv7Q+j55JtICOy1kh69IF5UwE1fLe7dyVDlzTWVncJ51AFDAEfekF
s65+7ebGoOZRKDE7Th76FdEXCK09EXJtenwCfF819D7X4gWb8RcmWTq4O/Zu0sZU
jn8oR2hsbch8mdMrqj3h1BhgPkZOV5tvN1vm48eQ8FKDp1u1A3Mh+JWeCyzy0+Os
Dc++TrdEPypxrs4SZ+dzMe/keJxLD3caV+ka7lvXs2yFCB1gsgc/dC1CVosYNeYr
XZlV1s1MOOH2xTctmuVUbrg5a4dX4b3AiEo1+Asnexh+KMZD4a6hG4D+6dNobH7P
dbppTlNGeN5APvj+PjFuK5t4K+vQzpARYIX7bJ7HKlrFH5hVFm+0Usl002jjkrFU
cWORi4oscNK0OynY1BTKeoNJ0IC8xRjgUSk0W2W+M/oRAoQEbTbPPoLIIsxBAeIi
qO/QWffjOuSVp4wIMj5af/xAMWAQNauC9vUbCZP6KPzh0r9EhQk/cHyZJ+pPmxKV
4/ebnW9AsGc/suhd5ccFJTbuuirtZvlbNyWpHKsKMkWNJDK0U5dWr8sFqw2is+BB
JvytRuYPXMJsoLflJCn9pPQK8d/rYWOou/eG7T5/+FZjcmJMFZyMul3/DH1vbQ0s
ovHNv4Hl6eBHcXqAto3Q33yJ+Tso51cvBF+H8HQNunPo1rURyi3RX90DVR8z578m
UknMZzeYuD3Nift/xicKLeFw6o5JRVDbfF+Z+or2GVhbmgBlzx9thuhj+rd95w7/
A7lUGXGjwSXq2MPtaROnmra0AZFUQVlpFR331pKKi7sKtdTydxLJL6cWZ/dnXvps
VG+ypQ0OpGQHmmq2Wv0c0yMW6FxZn+RCAFWj/dKZTJ6Q4tFVRWQm4v33vOn5AFfn
nUFsyDzoCiLxc8mNAvTiLGVhd9fM/DdkqcmqfhChRtW1uamoV8amdr2WyBnGFF8I
rlapq4i7X5rlNrACs75vEDBkPjcDdpvglZTwaFS0spT6UhmFloOxgUl60BpNxCxz
HMS9nvoEo1MCqyz1/z2ICfsdYl9N8P7JgaM95Xz3w0Qog8m/sOeZrTgJKt5J8CVB
tdLULCUNqKx1VzCgvYRJ3MN0QBuPHJpFSMxV5lbNG7mlG9WeInmuvA1aS/OYMhXf
2APWrCXD/D37bHWQuVsrjNFaiCFg1aw2ONf/yKsXy2l/aob1p1X1ro+tGi1duxZh
ATmK1YBOW2zUkOl73xhrVlmaQcjcOG2D6uaX+AsLktchYUVDCCASlriS73xIHYxy
rI3mRJPN4pl76Q3rRTbtQBQEa+lgXGJpbKGtzNZNUPzTc2MuZTsAdSRvSBi/ssZI
Nt1tTDo66D09ZCsv34XGyNWRIXRcSX+6Hl/ICkb9WcDdv7VZbmNT2TThOjA5VH3e
qTXQrn6IYhTewHVUuE61+3W3Z/vhIzixMG7f2NRcqEI+TD08dLiDTFOqWKuwKTWc
vUQK4U/E9HlyOSehygfNaTge6GoHEZVLg5vuwcvHYKDlCsdLQmlSAtM2QX2lRhuR
iHUBrkKSGk/+DM8hzU13YDvTU3zV2r0g64FXMuzciTvF9DEJARjcvcsWGaezqhlb
PHNIv6YuyOFn8Xp3JpiN14+b9WexSqobqnHD/lJDuHhd4WOMpAMI5NNrQYarTFRb
C1t3Ve1C0QAuXzh9MjoIt6U24SQmURQeiwR97+dnINIwDzQuJqw0qxtvjRFOncux
umcfAnECcUJ+x1eTuX0XiTVNvj0Tu33Ce58rXfN+bfZEr6Qxahceyb2eiElCUxVf
AqF5b6b3Hfo+muHPU6dO7OZjNTxHAAQi4hr9h8LBnqlRKw2bGkSDoAOPCSqfQyXN
GOdNUp104+mOZzwuGEoOZAPdwwnjDx6Bh/f27wAnZvauomRZ6NK1P3L6/cj1XwBK
FBjSe4o+uZd0BdmqWQ/CDeTTbNBhCnDIndqh96obgxqRxyct1BspEtQDnWXpZpJY
fIVPnMjvxWPHvg34DQNMeLJvXnCVhzhZt7fjkN74LzC9GO7MuYLgyWvI6en/+bFK
G/fLvS2getm6YtmjBvaq560pWgRiFUiKpUBUoJjUn7+US6RfkqAg4Mqg48vzOJTO
3jtZ/Fg+D1f5f8jaoGHPuBp84o8p43iRa2DLES6retY1mC7N40GJwQXoc54AA6Lu
3wth4beAa0Eo9DpH0H5AnRTiTJu93Gulefj8n8BQq/xsDMSl/pUjHKvqXebWZcmM
dFc4LJkJcWabuIiEUpsKRPKNGK72Dabfylt9ylJrkxgOAAzG4yx0A6L4FJuMl/k/
/2lsBWq8KZJFUbAHDljYCfnsQtNF+ytiGYPoJRIh47u56MWpy0+MKOBQzU41lHcB
LT4DiBOHUQ+ZfnaQRmKTKc3Z+n4skbBcxF97ztX5ehjwopiQHykBbTQGj7ZpJBhO
4WdTGbVbR6LJVgxQ9DkhAOGDY4brSV29AVik+hHOBIIq1r0d2c+vCBeJyNAAINzY
iIq5sGqxmuiE5ArUPuaghpXL2FEbC7ZUHfjyvwEwWz/79kawfmotw+reriOuSrAe
GelDZsm32kiQ4boq4+LYWbPFf9o9wM/y62Gs5Ka5pTM60+WoLfoxJvItXK8sLO8z
Qorel5UO9cydcCPa18i5xLAKJjYcQxsS8dhw/v0bmf5A8LfPW34qRudcrYkv9zzi
Wd2r5JiCHwjIIPVrEnIs3rXX8JsgYK5Z3t4d8CSET6XJcsNLGU0DX00Qvc7ey973
2JUpvGtTcSqxMGCEJWRTsddj2zcuNFnnGfxAgxlU+0YHwybpQza4MlOQmc1L3ITB
Eb8XTjYmyemhIxJ9fbByUKJrj5R8tPKGATxb6+axBAb6gLGraKeIKONqV8LBjXuY
YZcmVeJJE2OGMemwPigf60f76fO1NPc9somHubWCiZESrRlqP7mAQCDeE1Ry2elz
EFuGM597wHfNxEZomiZ4+DrK2hkwtsh8UVoUktYkEwV1fUBV7WV5hn5uVLdCyWq/
NF3yml8MDZXCXq8zrOPLrME4WDjQ1pGmMFTndx4mQVy12IuDKNc2Tz69vEwwxauS
cg5Nakh8zrg6Nejfpk9ALUEMl56WORcN7YYgzq+45AqwZpI3w9ye6TzHN3FSuMpv
AHg7QtZCaOUc9mdw3/vnOi3sNuClUtQ8u5JRNLPrrBK+c/ekKAKv4arMhw2+/KF6
9fAlycXkS3eyeiAzuOGmkgdktN9suXBhZ6cn6Oxq3qRdh23rWUpHsSYah2F8WcpU
rmAjH3QUBRhJyk3Tvnfq8KgV2rCEQlLytrUm1n5XEGq8gHEvvb1vswOz8IqHRuGU
NDwEdXmaLGKFPbxrgsqw/HlRdpuvL1AJ4wfPHyNMB468SJiAO2FhTCDece1KyOLF
Gtes0NYWY253kjAdTHPIiFaQHSQVmf+CoFrKosP8uT2HJWNoYodxiz7Zd5AUtTus
jlYQssrVtQpohR7R2o9Aan9/FJiLirqSO5NZZebyBVA5EvFMYnBIwJRLHl05D2vL
1D8nn91pDp962JszfHwGhxg02qGzQeH26fhyGDCz825WPRuN7xzrzaC/QzbmXQGA
tDUMKUC0/doaR1mt1Sh0LpoQQg14ddtmXRbiCsMpngFWTmtZKUv+ZX/9Ltwp70Yx
d05kBjrBz/Anqubj2Ikcg4+8vrvRcVR7QrKuCHWHmxGg4oE6yFsMgseSulkRjwWu
kCxlxSGe3wLpaqakyQp8QbrCD7IhGyY6lrqvxxzO6LHpbmjfbRBD+4s3DMo8/JO5
vK3JQo/HbFoPBIHd3H9dLMJmLYGkDVfhjqgTcaHDF57dcxJnDbr1g6LiMFtZwZo2
k6P5Ab7tlVoC6zUQJfNXTF3FYDOR+a5S6Y40WQUxaqmrABxuA3F4g9toxHYp60gE
4zzSMyEPH0xqOZXBiHjFGucLmQtyB2hhQ926GSmfYyJ4YtnBJu0XDS9nmEPTMH+B
171vvZCZe/SD0mK4GV/SQ/i+h3yeLmN/oO9vsBpklQrxxzIPgdWKbz3TdcTqoan1
P4P1U4+S7048Pei5hw7lIM6N1ZSCg2NoLcQXmjEfelPvwheR7kAa/m1ycdxyTcb2
Mtaq2LBckhRBqD5JFHnIHZ9OLk9xOrbYqJUNz4Zx1417K2hW46iANK7t11yCqxAP
XcAPcnqxg8PHQL2NEHiSlgunFCc752vRCK95PqLVWRGSrVLYGv4LLc+tCYkUKY4k
+NHW+IUFNHWo7Sx0JOazuHlpvujrHwZ0wpsAzxqp8ZH8wHNxPwf8WITJjy9klfS9
oyBOuh4Mh9bQYVaxnhw0D+eZvnk9yVpFRBue0BI/MWI7u4f88Pr7Sr7sjic+Ly1W
TfcqGtvXYIENR7tPAxHKVldHbErZiN6qRTo+PgExDZ9FDKGVa097dhC1tB1vMEIb
MAl15p4LeqQ0eVJ9Raojar0amNEIF/Ryu9EmejOqGdtOVmuHnrwTveRG1QZdekKw
++U4I6M4TFsXijV90u131Eqh7YcGl+jyKErEsqZrzw3wc4Eeyv9It9FAr6Ylw9pa
sppd2qdssykNNutmss2NxwO9H0BrhG8lJrkrP8sw/fstFnqQLwjQwNdo+1bnJAYW
HfVY7gwjDJJdiAsWMese6NJI+TeWv8TUncGlZvn9Bnb3vjn5MI9CjF6ET9l0OPhV
Lmhalfbs67x+v1aI92X72ylXVWnA2XAijUVvUu5zH7iLQFUV//Ggm8y6LJrBLfJ5
8YLq3sjnXXuQJ+cqZTZa2ELycd46RHKtIITqWMAhfZCENYJrq1Ys26DbzVvnNuAk
MRts4PVZZ5Za0xvPvgtg548QQ7yZc7xFCeJQEU4zssGQAdgxmRyWpkkMbOvM2qB8
Je40xV9ZHvjhEz3mp5d9Bcdlm7cjKWhDTUK/xUbGvGQCmQYRzvVxbz1yXAh8bWCm
hUgk8cLawG6XPNdywu5/ZAkEfNb3X6btQDhIKUGL8SUzm/4vg8cAAyDFjZgXYeN1
7cx+GJAbf2m8iUy2IMaYgoXBsldg8iiZ8Rjj/sJ7QElVkDPC9rK/kShwFXoyQZKN
nudb/Vqm+y5d/3IIdaW4C3u5x/rsiuMb96GiaEaFEz6FYiv7lgSnmTKFwB3cwalz
nUR0fr3+xTpZCEDGVXLSKP3slNduX7AvoAkkLg3KzabN55H4adCMCEGIAg6Vuafg
lPKSBHnvrff8BEu8ZpeqIRf4b25OhV9pA9i0aV7XrBAK3sNu9fx0gqLa0T8TJBzy
cOBgX97dnU3tW46I6JFq+ippx+EECFqoRPQ2fwUHMUGEA1M6WpPrCI0O6Za0A4Gz
s0XgmLi2Ffptfk21nxsl6qlkOtDfYpQIPYa7qCgVq+akmnCAuuskY87rYtfv0y1U
BRvTR1bZql2RChr0dp3xQCiYzUMuggE1OAdyRbHqDH1adXVZ3Ybc13E5FKonWyeu
f7MgHX5Azhn8ZAKERQyB1wAvXO2mNiTd3ZyGXPtGiD1yx4/YtqQfJWzGynCyciup
Ob/PVcZ2nBiwqCsCsNypTrs9msndgcSfO4rP93gfuKflt/sEgeoyXmmi6yKexkCB
sqOPbin6t15x7KuqOO/27ZVwCvmavBDkfwSToJfyzaB7uSaGGVbAQw5GeoWlaDyt
Qd3SAy3o73VYBbHDaFeIR4/tMxFp78Iom9zTgGFzAh5V8aIYe6T2X6bshHo6qyuv
KMJz/2/STv9cDiPSHSak8lPIJJqSXaWV+tWzRkG5FKRbxfNA0V99FzVXR267kZBP
9hbN5eak0f2KFR+c4bFl89+O+BmDixZjdV+RRM0cXN6WqiRedM/AWsi8FByxoBzD
CUHArEQ37YqLXvqYbP2Rg6JahJT7Y9MFvlmo5w3cBAG34tU1E5qkbrtjDQi9R5k/
gmkw5f9j3fOUrZ+Urfb4QnDVidhItIx6j+qZ4e380rrXLK+b8iKvO1zEORxqHxLz
wMIUOEAJ3NRXT23f6Qudrn4asLOoaA/xEsrHHUukkbDbM0b9pHtwsd0Mr/m8i87U
VH2DkTuM43RHWdYaejLX7eTthxpBkLqeriyp8mInqlrILYgiNocgGk+DJRH1BXcO
dlF5wlKhBWRf8Ef5qSEPCmafzKG94KR9q/vfhckLEvsqop9aggIHfVfQmzWE3o6k
+W30iT57mil+ZFwyvJh4ywrV0vjIuFof/HR+Lr5Ed/2tR8P4biOJY36lyRfuPCBT
ymQn75YzxbY7WveDqQCj8VJOmnLcLCJz+Pajdfy+YDPCrqAz+leeOAk+TLugq63o
z7gDEJlE48z+DZRsu9q7EgwOWFiD5Oc93IyOC++5WPrRshjAPFZxqTJcrs59U85g
cyaVDeD/zeiqZVvTR1k/HwKNRi250VybI8NcB3tMobcAuaXXmSjIH8RQEtMWG6UZ
w5nCXc8Vv/llnNTwjMfH/TxB3MRuS5e70WFwQU2R36KugMHYgfg4SxaxCYNgqJ6y
18EQV2+zvzG8dqbp24KgVXmZKVLKahT3P9dG0oNb2vlU6h5ClqtX5ypRLpkmynqW
tee9kWnBF71WQSWCre+bry5YzDf7MS22DCFpRc3EY7hQXDxBydRc14ixxN/71yNU
OSj03hi0uDqTjX+yDukmN+uBsmTlypUsh02tAF2J+SA2XH8X3IQKI1vmWA+XaDO/
3oi4iooayJ2PNUYhjvmUth6jF/Q0nY3GvXZCg+v16BSHaH5GkHt5UP24aobSDflw
m2c1TV6lBL6jLxcBkZ07oz7f7vt+cxAg/Ibz8HHQe7Fu5Yo+SP1DcfiSZHDL3XQs
7USy4/7S7geDQ5GPrD5naE0j8SBd+RZLelu8RxtldO904ZgXSxvEi0vKHQVdtfg3
Ss3wCuWbuJ8lx3FlFun4nBDqYhtzrtRZq9QDYm9dN3mJ82b2wdRNij1Telw1Nsm+
y5Cq0SP/LR0Fm2BKl/8euOWjokJGahlaoXWymFSDE8VWfZ6LF63kWhq2il+cTojS
y9ccpUgk79afR1/nEYcKY1Qr7QvZDNXGO6LEAyaxGk6vquCCeb2T1cii3sntehMA
u5M0pZmlkn5g9VHCt3C8o5lrqIqqcADuaC3nCpJI3Vx6VQkiJUlnb+/xLmMnYxVn
3tm/bpk2h8ZoM7uT0MsE1QELhXj9F3dZhM4LUjXjeEWovZLZhz+8EJzOonRLnbb9
IBV/wGDXrtHc3JTMQZ540emYG/Hchc4kdWOlzyeg2XQLaIQdBazIV+wM0oWs+tBr
WVgU6Q1thhWpQAABezxuUZPh+k7fO8LWnvQInpeZwhggL1jprFiFm+N+3rpQXllQ
7xo6/f2T1sjGxUMIfAqejIJQanMBLPsc/RY6SIDyuS25PKpOlzFtrQ5/zQ5UmIyi
7AcyDX8tKzWfOE/5WEDiwoqoj5eQamf+VEEXPUiutBaAxjnnufqHUPl0qTY8uKUZ
/Y5ZDhYR6mUQcr3P0loqP2m3yyGBsWSjGd7SUmjYwDrfjPMce6TBhzsxBZ2tuX4H
s4y1BWb3Ej26z2qfpp8SZphV/ioklM9tC8KFzTxD66RDgF4vUw65wblJbaODd0LT
HdSFWs0HJ6I3Mr8PRMwwDKRqBlYQpt+TzVrHRmEw8BvruAPYWSNtdFzdVa8DtSjK
JAwilluovPF/0+sxBHz14fUFaktTsXAFFyI5ZIW1rHTKd51tfv/fuUZWnlAV3/OY
qNMFuQ3yqKPwyzD8EmDC0/pTB6qa3N7j8GdD2lSrUu+gQhJiTmKAodd4GwNDtDTT
iBQHCldYyHRgX8xgrttbWPURG2VjJ4dkH3fZ8VNiBcTu+caEskZzHQ4KAO3cPApv
ELilW56g+W44KXaQkcP240yNlMHl6cL1mJbIIxMLwDEhljwgqo/+DIU8efHIRe2E
TRFo6LyeWbX5PY30/EI3rNq1FcIFlpwkppMMeH5kwK/ZLmoVZwpdi+5VexpUk+bM
tNvUE9mruo2OqRbo2uHYd3qpfbS8lc29gfdiXOYkWBU1SXS5gZ9w0wMc5YmiUvkU
X1VdiolYQOIqG+NGj9Vyh6LaZw8j9x64Wf2FWL8uelVGLEabQ4q11dGqwx8viQdh
x8KNwM0pbyRmew3EaKzeldUjtYB/7I+pxEiPCSnfrwc+e2fSsIEoHkDgb9iFybsF
qCDwN6uQQl5VPk5BxHf6PADgTr4caI/Tu85PB/0NFdBa6t+w87KaEzZ5ayVfVzHb
StD0VRvW/UnEyjTvWWiMgU6GIMwlBACbuvhHdSGvr5yiMpdIQNLzcjaK+mPWlksz
MgrUM6tu4qwSuDgHzNq4maRL5vx3Jd73TSJ2jJLC5gOopokzFumhfRBdR/dwyYct
gmB57AXlB6AOADiIXQQwNptd4bl92YKBezJ1Czo8QaF2cDO5u8NQuVqNM6yyNaka
B1pzErqM7sTloRzbrNkCQkJcJAukyljBaTu9KS079owJpExmcvv6HrjqKNaGFJsB
/sWFzVKJ5ARA7LctQUoqEjE+Nuov2ir9rUExJpsf2HeJN2rZfsNe43WRe/aVi3iK
5qRF/jndrsgdIohN3dcNIqJsxdOIlH99319O/awXBUGURCF8yNRxfMMoL59oAE67
/kGATTCOq9r95C3z2mZABZeyNtMAxE8oNuevfVnOSkbZsIJ1pjRXnBPWLn+5sWqK
3IrdkZu6TeGjIzG4NAN4iwbrv2b4Fp2PYW2p6Z3oXBu5iJ4jkdcrudl1jzOM0IOO
uzNfl1M7LG+P/pnnR/JTKmlOuUTZ6H4+YKvlv+duJ2VtETrtX4mdFVz8bY2XVRQv
VcZWmnxqPT8qO+Bt7XcaSyrU7wyXuzP1jNk8k88TmXm6p+1hZXR2aouUt6onm1eS
5MD5a8xDYBNTB8T4zmkMmulbkiuPW2BG5bDIalQ1YEqS84x+GEkqAeRTTnyIWDPI
pC2zVI064c+cDpbVjAeboRAcYUwPYso2E1D6K4YFrOkxSdV0cYwfvcUNgkOkq8DT
3P6iq5JSr9/Dbn/KveoB3AO8Q6hjZnSnwgIg+LNtyFWKs7+BPemMceuBdKPAvAFJ
9Xk1BGXQ4iFoRLJkxKN7MhK6iGDN0ql0a/HDtHEYbDlAuaf+AlMd9AQ1TBDzoNfe
gzFSLqnff85StF15SqvR/tAhLcpuDwn5Qbb/FoUfhdtZo/KEJiKK48cs69chmZY6
reF7PUq6wM1ccbvbX8xbl5PzuGid7DmrBBy/iu5Wz8Ao2ZEMh608cZPFeB+m+Yj2
fvo6tS4WjiFyqh8tQr0gJjQwzWYWuOOLvXplMdt2bamrHz9jHn8vzHRmffQTfx2p
EnjfL15z6Rv+VDZUNDsJEOfTMHtEENJa5I2VrOSr5LFyWm4Xcpt8QK3+3RAjFJ2d
E0X4+K64y5WOE7SxeLo/Rq3WzoBmgu8g43VKb/+stycm3Zu0HqvzpqwQRkOFwAGa
eHRSyubKKuHI7K4kT5afbNpVR4swYosu8aPFhf9a2QfRb573gVoQc2ZevLN/Lz7K
eKlbTcbaA7NDlgQlI2QirV0EWgNGo2DHbZjnLQsRzm32Exo7VJmUEtY2vwUOsKi1
EqYLtazhUb0js3i1E3rpsoUaRSYqKzLfpzby0cGiek+kurF+xmko/bBLSMKT+6qX
REyxsCKxMTb17UljesEWQFEyo66UqlQPz1kyY3gQR6ipeO8Vb2QXLvTpu2EV7xt+
uAciAkbnOoGSSnVG+UmjV/VQld+VdScoaaLWCSw4XtfIruhuWdGnjbTsWnpPvd8Z
EYcjGdvYQ2W+9yNHGdBSwIwy706hnJtHHittEoTHp0ZE9mcenu0s1oMyHTb+oQQM
Zv6zJRUM4aPTAcSFd5HTXjtijKGNBe8Le1E+2Q8ryp7Yh+/W4vp/PodRQ7TddFHj
YCp2KivByzhp9MSsaSK04DH7RYMLqipGTnpNKTQ83Q0W/GpEazBkSr6zvW5Scw6K
sVvzqV2YoviaHb368vKs2qSOA39h6jXgNSAaSU0N1XC11oGKLi217U6A6BZHGDal
UICh7zizrVqTKKhvUEd4i+A/PgkeZwneGTs1L5Ws5zN3bXy3y22qxisxUMCImzz9
Lm+KHEkQ4Zj/THEJVBH5jSwPJ2L0nkBgY8ZEVWfJ6REH8+YL74mH/sK69Dpd7nNE
AQocSDKP39T2RZ1FFT6pnN7wRUm7tRby65sRvTpg75gj+RrN53AnpDD5+nejoapG
kfy1d0iRhmi7kRZfgnvPVBcndMs05xe9jxIa4HSXvQokUcre++ahk0IYb+ezRZj2
swFclDa8GSt0nFeGDNsTtJ9wshJ71LoJNdN2AIU1FXAZdp7UcPJQzrAzX3bc7Icj
eEeom5KudcZEtcIqNN4dG0r8i57d2/itFAfCzYEsZE26GS6ZKJTCkUh4kjIZUuHt
vIIh6twxBB0pOqNSWO+vMQx9jEFiVQXGbuSCvkx2UB89R8ab7W6uPK0FV9OtmSAF
9bRr7IuUTU07XKajppK4FL/w8BKrgxwEIhITmDe7Mukfbe+L6zZs3dAX5JPTn59n
a11gMdysPlyGrCzs+jiKb8bcUsn9ovdCIxAcv8PXG9rC8UjSiy39gNuY2zin59m5
HEvdxMVriOnvF7xrDbyWN2sxnVvPdb+X9UjymGpVNZ8xd8qZahtHuHh8lSEtwelT
rDAoJ6WC6y02J63mneeJe4jDzSMZyeh5WNE4MuGNhMQA0IjkZHFyYB/FltRAEs+d
SsOkKRrnvxf6+tUh5vSvyA+1EocC9nRxhzxAZvZdIlR5D5F5+U8YcRP8BS+x4K39
UuWXCzLm34+9iK34hGTqXW+gmE4vWg2pf4eNSP/7v0G5SgkP0REpeV/a2xfVl8QY
PtibFX/gqsJZYksrV2JPWibCZ9eBrPhzExuQr9S9usW/Hc1S3+VkPDmtHNnO+ehf
UNBlUw1qARafeabponUg53FkRyJA6IyuOJYD7Aak7EwP1rxb4FbDHY4MExMDor3R
FYAUZVQsuX/k+xSVmxF2sOjq8Ho/a75xi5SnABzATGNalNywWqPtRlrwT1KbHF1s
T17b39VPyljwZOf8k54ES9EDWK+lDHm1pH5qxh9T30Ta55VIGAup7xQ1uwHF0OZS
4HpcpjHXhdbiAfrDLuUVpptAQ/tiDoibOmx0jp9oR3alV5eyDBWsGowe8Wkhuq90
wj1LGzmHY3vrTqO61YVljeZlvu4Q5HL7fi5RMBZTgU4HDeXv3o8vBpEVB6cHgAJH
F9uuLaZGIrQ69WpIXxI7ILyWvRW7HG7ZSnS6G/pWeclEy8gc2n6gZK2dFkECLUfc
tUNf0bN+e0XII7AQxr1nyedgYlYgMauMEruCeVgkq4gd5VhDGFQaTgMIyo2Xe22f
a3od1vpNt18nvehLGPk3BDHNL4Wpwb70i9SeLNktc7+yFudz4bJcmWnvrpSIgmd4
uL3YVoZqcmdTFhau4mpoo6r9N3p/epWr+zyOvA2wQNyJdchbvLMNm/9y4UdlOfyO
/VG3EBGXApc807slda63iEbyOViPyHNIGNzYs81sDcOvOLrvw+4h+GF5OScvBLgn
Ke/TQOw5Zy/b8yFrXZa74UQ+xHA+nJtZQ13/zG9pGDr38146EExP035IZQk0hq+c
WNMkzN88Qb+Q2boE6J1SJuctssd6AupIYlvmnwk9BI7lYJiVTAQBof67O/VG7eEM
jjGAniHTmuUM1VjeBiqtSqynWWmViG4hcaIieAIkXNIkA9ix4hW7Ca57n8seL6m7
X0oOfxWzAXVMZFnY3qsCHuyfvsFmRyQaSt4UopN3CH7nsff8BKvAn7PG6S74AS6Q
kjeRto8Zq4/MN+2h6MBnHhOcgcopSsV+zDCEX5HG8uMxv8gnmXlK40YFkHKZtDBs
7ST0rT6pm6pQCmGLBxtV9dFqj5f3pZIlf9RrcACajSVKDpkMxDfdVmWeOOLYMJpa
fEFM4JcQxL1xJjqAQd8TsnsP5X7ErrjuY5kmggoFZSr7birqEaC8GsMImlCC/TB/
CD40KhUtv6wvYyupLgLARIVwvYfHVxnDaEAdmduBrysf0g1AyFCPYZoAWJ6zRKVK
i+p+7AXWxgizYKPciDxS6LYMwE3VltWjohlk0IgYczPUz1aCAkKUZkDoQur7NGP6
GZy3boohdEj2r3puUsCHS+lJQpXN97ynlQdw3kJuorj4sVPzQhM3VOKegh8L3pgw
Iiz05xmrYfIFDtOZ13+bTWuWRPiRIS2MPMZKBErCJBor03unldgaG5J7/jjTpriL
qQ78QbUKgauO62RwgrhpvbbKtTUhqb8S/NX53tlQh+sldpwLa3B2cF86bA318iFP
ebYIVc0IVE3V7zJq0sKSppBPjgN08gGTEkQNfQPlQpEsEqpLDOODaok9MQWD9f6W
2NSfvpHEIn4CJtsTHkMae8C3aeH1iaUpZdqs3PJtFUnL4jh94eo9SsFSBggcTAsE
et1mh6lTOI1ZXRQNH7fRUkH4gjvnml4q1ZGgT8sSKoPkgHKTtY5xbQzUaNp1VrNr
7t+s+wXby3SIro+/UzaE9S25yPgwr4gYx0dC5HkL5Clk9+fhUBgoAZfD99dmrMu2
RxcgULyD3m9Wn7/V9NF7WL+AODajdTVOH2r8gObmS7d83gk7CN/iI5c6RWabP76b
sszoVty15Zc7PBOdQ6P0JbUoOrOLlfKUU+9xpkmZHcZulDJUmsA+yyeyCAl91YFZ
1YZbuIj+tgm4gBLsZ9Yxbw0I2LWwQRS73LaEysT/CcbaezfCpP/0hfeNZ9In+Uvu
1y8YbeRQ339uhQueoyz7DnEX1Ms1R/Rx4Ir+0CvU8IP34+Uanza/m75H73NFuWrg
pYAwR9BWIHrRYDLe2F3wt/ITg55BFcLdkqsH4f4jYo7fVQbexsJf7qjryTi9Epea
fFhsuNu823zK+o8Gfv3Ws5HxxXPFvY3sPwPTpsCnU+zrIIgNmZsGBDG9ThGnsW0g
i4PoqvhdzwD3M9nRkhn1lrngSAgUGlUeg7UphrSXaI9njgwb61aGjqAQnGO/c9eZ
84zkcdyo/pYfaA3SCUgRaP10WIlnvE7HVfjpX5MNg7WVsaiqBwJPbCTVry7W2lTZ
orwCfOSNyBq1g1pURcfzl4F8hDPkfp5L5GYmeoPlIR7bT1j5TtvRCTOrWWkSNY+7
ANYeTpV18+gJanVApRbbz0e4KRNLhWG/vY4fdyDSp003gjLZ1vw/KETa8E4bE+2e
ZPBkTxWJupYJEN0s4rvLbHjfdcgU4trTtzkXjqtUAgrkGjHwa8olVjAl+Ga700JN
4Wa9RPqfEe0HDIQcJ6h4693Dh9Gj6lQ0IGi7fdU14JzEeIDEnHy5BBJFDkBMMIIj
I86YmpLIDJlFsQq1pvqoEiiOnOLBbB6t2mLcqKFN0f2juzXRTFTbGi6YW83WHnNS
3ZjRLMWRyVYW24Iqt1Hv7NBL1r7QGGPj08EtqXYrJ/snI5eLu20A7muiT024iP1o
gkNB9nSfJti9X8x7gNDwMGyEDm5Dt/LJQWEDt7mjxR67TW5MKvHxZLBZQ63HilMR
EjCXGNRrKAIvElIZSiVaoakmF53ggZBv7XHkHaQlgPuDhmBWpiGmLW2AAMK4+bc6
H1dM6FPo62UEnxlNvJYhw4/b4LlUrN7jXrRA3ei7tG9N9qSuieiLgoq44RfP9ljv
6q72RjYCdY+qLCsfg9qopR56cssgRpZuJdMyyWGbLW6J6E5bEiAtwNY5X+R6C6Jc
E4hsatXxXafBXQoY76KRgQf3wqV2JjVPrSzQOk+EKREGNh/oZ3/og6ZZpU6+SY0Z
AGT7Vbj5LEWhCJ7QLC5Md4GTWPw/YRrLxVfei7PiSzSk7PmFIgwyFydQEnXldRV2
DfNvCV3WTnWfNZ7bHXdAD8jUEiAM/vHZClE58kKNXDnnWZpY8ZnwDlKlPi1yORYw
uNMIKrCCXLb1CnKVr3rPezbtE7x7hBu1sbH+9X1G7wA71b1NNy3FmRkdRxbR7h9Q
tqg9jP/iwtmpOhXgysNWcDxh1lWq3WSBmdDWDPrGVk0nEt4YCWPkbgzi3skbok1f
SBPtdaPmRkRaxkCUoNnbhXCq78JXfmNU5lA1egusigPsnLWLUmxA5lNkbhbfDrQR
G6YIU0V6qCJUKAhwWZ1HjKYDbwQUEi7JZyHkqSiAm1284RO/T6hc0LcnuU2lnxbw
XJ+S7IlRtfxQfv5AsCq9PVeUWnZtsHc8ynkebOpn/UjRNb/cA86wGLH7UVofTijM
JhyYvvgda+UFadDr3e/k4DgR3GlhvBkKfu0ZHQbc8AAR467rVyN9m/aTGXu3VvO+
z7lfbZs/cjp1k4HK5is+O25AWRGPY0eoUwFQbvbTd54Y8OarexsafjPm3f4KkFdU
Aa9WjZCMIbd49F0SX5WeoPJQz8l/Gjc2H1wGTTcNnrFivWSv0hpv9OonXSJ2ElVh
GySgvjxw2P+06QruRwzgBxX9S8eV+MxLoND47/qvzX4Vo0PBbN3LNIhdE4MDdTRY
KQ/HAeL8X2wsnmUDLOdMRUOBjqj9X2WcTrH4DU28qms1CZTjtSHHCkdZlLBvoPjT
RmLao3oqNMAHGuXehj5n9m/gTd5CxIgNQPkYk2CLfzi9/+dcLqKgWiPwkUFTPJR4
5JGP51Lk+m+tKnzVOZq7ssArzf0p9RufHC9ysZWZSeYd1MA9lWI+zh3VdiSsgKZM
Zj5Hvmpo0RuiyPoORQoW/2Y/WeKTC9G3PXXH5ALClr46RL4QUaBqy/QIjN+5lIPA
78Vx8od/BBeygTMYU3GFTURd860zILVgK+Q5PLalFtaj5o6k/u7a5OFLVVrad3E/
p2RXiW75LjN+JHcgZFmnfRY1xir+wW7LdlK1BhhJpSOBaJwyavKhrJPsca3ZV1ZN
LMMOXE2xnbdFeelbGDVgHFCiHdXhnL2RzO2tAIti0188k70aifOJCGxy03PeoXLy
zD6PIPKLGISos/JZinfVNUFNiPReJeHQIs2C1EEH94ce26UCW4dUSs14BtCDlk7J
Pc8tcwT5Ska875wzx62GFMIRHar1FOGskjCGLb74HSkx2uimA/+DVLgXKzGBjxIO
hOdiE9zRS1PgRWZFVOlLfkz1i8oW8dFQcRJ4OQF3XzBkQhJYMEIqNDQ/Jsf+WhYB
lI93A2MSm/hBCWKdXfBpl1pyF1XN+n8f/UmuxcaOmdU70LyavXpcsQBzfao9RRQ+
zdlONWYsfcfkOSLSHAHE4MXXqk4X32jJ50FrMUL9RpSzTnCUFB5IGGgSODWG78KX
9+YD6qOUFz3kFGzRdwWMo6ln9M9cTay4uimKrAjmFCAg7Nnr2twi2giAQLa3S6SC
ImVpl27ykTq1GY5Dv1b+swm2H4M8dzscwbjg7cEGWOeNlBk5iUB4nWbd0qI+Mmgr
o9LXzPs2QAg4lYqjXuKl52RTZaIhH63+u0P+NN0kXJLzFi5Zm2pzoWGUq1mV968S
46RcSZ4Fm3/rsuTxaceMuyhYviGiOC1Qf2sGxifgivWeg9BTwDhjk22s3nz0vDEn
RT9EUGVz9VlaOH+a9VXxIhk6DgsFuZztyKwfH2NtDrOfolud5mQrZDfoEi4QcbO2
FKazttUJ8srWQKemL6KJJl7fVR3Thvj9thJMRY/7u+XXDEnIYZcReN8HT5NxWY7F
57pasevqlC5VCuy7K2Hh9hz/GdB/6jE8xD4yNd97xjaN/XpV/v/4tBxPzBqtMH23
g4jfm1zst/olb6lRBNJTiJO8PjbTn06Yl9wRwgricEc7LIF7152X8DsFFysPHY9G
46hRaYqNT9C7O7qck3LA3eaIrNGrVLgvRZ52HgsPYYV9hgombSBNCevg+Rr25WJq
93e/zzYimbSwbt5zg8TqXM3Jwvn8riCdd65j4PH6QNQHR4A8mN9Y3cdfbrz4zgzY
H0RRmGTNKcuZTIn7gcG7VEdS2GmVZJAgtFL+hGfXJlKE0N47q0omJP6okXtluk45
M6yPwSswfQcZsoHMicmPqZ869OlJ9F/eoSgl8xmMGAPtgDArV5idgFR4uls34HoY
fEdHhgfJoqmaHH94uPB+xqEsdXOa7fGqUxuiwyLjUw1Q5RA1UJx6iBp7tv+JliwH
/qVYyywpe90wkCeHUZnp2S29CYojyJOgGUVqcDbxJrjRvrXwAvoKFXbl64X9LacE
fzI1YutNF3Dzk2vE9qqF2C6pj3dEoKpOzb9SxFPKxMeP6Ys58qabQd5deWAawntF
367XJjRHSv3lDKjI86vgKLgQTfWNHCnlZ1J7PWmzozl6ikU9CXm6klYgrufh2t9K
jt3NtXCS4VepzDEKcBgVrHZLxdxyubFMPfWISXswAsH0j7Wyd5gE9NYvYm54Slwk
tAunv3WtSg4gtb68rmwXMYuCxiRlJ9DGmlAokURdeZtUWzhxAFo78OyBXnPXzn9O
92X5xs7fKL9K/PyfDQ0FNzdmPgNOaB5m7NFUvGvlO/Sg9A4UqIkI2cI99DaEst15
JkPUuCVvjt1yt/o7PIy1riMuCIgJUuODOr43219ETnhmNjLNyseJmktIW6KgKq+D
uAURhMpt4eBTFGov7Ij3EUGDzRGZIWVQ0AV/WM6GS8zYJ2kAchlGsYR2ydw+x6/D
8pXp1xM1MFmm1miXxg7XodUWEABnJt/lvSIxSAmpkWQBlCpnGdGwdCjMRhAON7Ow
I28SzEwhJZisy8A61EsCQOddOvlAQc748mQl6Zg37VcC+xzgT9o1Me4pCyRyJdom
JNZ6h5gHmf8XfqsbofJX8IhUxQW/Uu/tgS4aNUfXnIFzWUIFSnvZnydQBvwrvAtW
hRyT1wb9XwGAVIAiyN6Hx7B6FQbMWvEf59TQSlT2ofgxDhCAhPh6oEso1ACtEqQ3
fi0tQ3YW5EpXB9sV7yoZ2eEcwT+lZNFjqNoeMxJt6+89Rz22X2CvJofqhDVHiyzR
CHvr5ljb9Q+gX8b7x3WLggqvH065EF9qSykcAwBebP8umCIikjQeLfQ/7e/esM3y
iuvhkWAQpUgbOVH9dfvXxr8xHffShW5pIda1d/HF1RNWBJ+p0E+3j8BZe6rxokN9
WioHi96ROo1+1St8PhThXmW/kniep/bPk9eOcAD0I3LbvMQM14dvjN9oT6AUtPUT
8KrJGPGM9MDCeFbhxwzHHjEuk3Yf9BdxTyX0rsTBhVhbvIIeyW1Tl39J8DFfEf2H
hFHM1uBt421Cys3jkiCbI6D8HFIic+RrvSdzpEW6aaUFbbfmYfxEf9ISnhuyc5Z8
GKwkkQEzLlDPcictRz1wUGX4QL5HMvaCPGJwZC5vScrm3QZTNuLxY696oWZAnlrT
qkFftYKy8NwxrHLt5galmjOLzgJUc66f1Jr3sTBHAMrF4EoSN7TXyRgTd9KL9mCt
6wbCxfn5SU68fMOvAHLJgnMpiWGK+oivT1GyFVBymC4cfUZGNYJPd3cO+s2tC/Ph
4GRRYl4jKM8yPNjsYCmfu2Wz7FkAuscB0B/fsGJFbeZ5IhcqrZy3kPX+QAcvlxWK
JAz6uDNbMX8M6p8BUV4mG1jfaiZWuuqvCyAN8dizyZn6Il+YmQiUqNbj5DUHAG9p
OCObNHGWXWgsHqym6/7uR/UlyXO9HjhowJyDCjGd17w30jbzk8I+uFA52q9QCncz
BqvnxMv5vg7ELWg8kKW+O6J4fiU7FLpidEdSLnAPaXNC2sppq4CmT9IdBYJxV+OZ
EfdicG5UFKkQihquJVE1+tGbyYK95rpxLD86ozpbP7RA3s7LkfjGhh7g68Bx7WGZ
o876CjRta9Nxasb4E0kch1hF3msAQ8ob7E9MgCixcLzGIQJOjoZBvdOzX3GD3oxn
m9MSifba++CxFW2/YyIZ7VbrikC5BMrvJdhyy80YeSFM4SWtyTNkTk7nwpqH6z/K
vWo41gPvNgrLpQIGfF09ttgnglmG3xt9p1Lm1BgWJ2PfgcrTiXUr2P/1T0M6iY68
MajlW2WT6KPiKuyYSX2N4jAulpB33CNQ/V3mIU+HBeJPeBbuthi+zX9RbI9PzYb3
YcsCOendUMiMfq3hAQ87WiEoLbLySDvEW7e5GmAM/jKZLtmTUX3IaCFAuuUSZqcd
4NYfd3UVz+OltwqaM2gM6yCdbP+OsSskilZD44xAJQKWzA4GcWFsRIDJdUcjvByy
liLEkPdhYI4RDhqzJsR3ofaIzPhvtd90yvLWjcb2fvJBcGCm5T61/oYyt+bjwWIs
/TMRESVlBhymZA7B8unKBybdT9WqymmMUv9sjIy7f00MU+Z1eQuz91s1mQGtuSZ0
bfgfTl0rsfNuelp+OdDhRdRGJ82SAI+O40Clj3XjWjSb8GCe9Y0fDWI9auHib7m/
NbHacSlmsDbd/mUEJkbl+Xy5eH3C1piSff6s1jqO+hCDv7dGCG0TrebHWy9E50hW
hU/0aX8WKUI5uH/Ve18gu6x/t0+1VYAakEvjVckM+sx+SumPirx1PsRkXRrEs3IM
44VehEncUCj3B5jaZ3M4gAmBEod1bG0tXu/JD+gVZUKQirC0+/bFfwtBEKHCgoCV
obr6MawkcMKXkXFE715rdEKXM3f2u2rS377BDFiCDBJ0g3lxLgzDL/smFrzf7Hux
r1mCDJCyFL9f2ASfJozyY1DaGufDjUIkkzDSMqo9bCHCGe+hUXlWwYhwo6qFHxM/
ikengBOForBItOWZBftCNitm10rvLqc9JxqhDqV1zclsrv3DyU91zJ9gL0DbgK3D
hv1eDnCgvjOfKgSJqs3OZ5Qav83BXYhfg7z6PYBAvCWGdJJzUImH1vEkWmYrO+XS
qSqbdR37C5HfY61L4dfNm0rn3PrYYEhjq0/CloqsgIbI8YpjvgfcpnO/GjfAM+oO
jfVfO3la3S9ZCYku+yIRTnWREETtXIPMqhCeNNHNBQZmTR1A/dITeWcV8ZvZcQxI
QJJQdC3KFvO8r1G1MQh8O+Wuplj7qlQbBydtVKh/2SnbnfEPBoWc18+4lUlERp4E
Yd9Y4Y1zL235b9fs6x+Ebvv6PI2tk7qIoA1hGWqmpNvPcN/Y9MXQHPZ0r+MMElqT
aSHcBylqiBLpJko7B3eL62lFbxteDcJqRQ+BJheAgnbGtcWw3z21f9+/qM657dfp
qpwnlc4fR2y6uvmU7qx7/3UYAiRtfJHgHHyFBUXiwSUTF9Yz00g2XA5IiTwUFEgq
V1Ws+b0eFK6VADmnDFh0Nifg5ZiZHfq31GuH4n3UagVp5/Lch1SezJ7Xnbng+CEY
eP0llGhNDvBiVm+w31UKXh1S4yPAHSwDwK2NU0K33GoQAY4DGGpRPTyFElnvmgXT
KFmOUjET0geqUO6X6FaqT3WWm3+ydrfIs1YA/EjDhbIcXVHv+ZhHaUelwHE/Si2Z
eRn6kMa9tmA+fhrXh+TGYNXVODvB7LoJAAxiP8IL/6KeMP/kKQmefvM4sLr+xljG
tnzAOKjid9e7qvIreotTuH23iFc64xHfDwS7tR5UN2gFp4FE/yFkbBVwdhB8+nWg
5pe9vzfzdHrFPdK3+TMDJbcVzJ9a8HT2eT8mawwXcFOL03s7Df+KPx8YBJWbJuUX
bTl5yFzK4hO+k+Nff9LmelF84mlu81YZ6bjXKFMh4P7lbjZLVCCoGotl82FnGTe4
Ik/b27+fEv1meOZXR3Z7/2RyaTbBKdkbRu4SxpOR0uUFGcGf07JUbvYbNwhR6A8s
PaCxEPYZXUALJfPdaPPJqBpfJ2VsXD3D0HBN857sBZ2IiXCrzLzIz5fPJoELkQCK
GZNEm0zAyN4tNKrQuZEm1ZKKOcqgWRmz2u50RKD5mkHpqvQtGSSKPH+vfbjHtIjx
RCdZkNhWMuL0YPZWNc5t6gAbz7rWLgL1wvFI5EXQ9PPvJIbtYF4MOy6rBCYYec1t
S3XiUupVplBVzoGh8tnZo+yjdkEkfxY+CbxGCcZ6BzH2adx0rxP1vNA73uEsG/nK
LWOdE+Zc3N76rB0TvHJ2z4LIIq+HTq6OBaggzDsAlbHFYz8o47aJNrnllvgiwO/b
hVv+r/0o4nUC3vDzZUyDJmyM+rV1wfCs1X1EvrWH5pnNH8wmgk3Ycq4dblgds6Tp
2DkMhxDYJUUdNg0nJgU1YmOYO8J79xDHKowPY3zPYKKlDRhslnChchSM2fVRE4iN
wA9DwO0yvZvGpBKwA1oXUakaMtei1cn+xhwRP7xMa5tRtl31Hjh+pXvaqiA+qNoR
j1NRO8srprBbgM3eRfEuLe0IaXp+RJTBMks8aPsAs9ZAbnfMa+Q5nnw6mxmOyY6E
x8n/C4b3PgtC26C2s+UKO8Q6CmN1kjWB6QFUoI/uaPFspRpp2JVuqFRnEwIDC2iw
mL9lSjz0RebIkon2QJ2aJDHe4MXWGoaXitAfvAAfLp6LnCUfzYhyw/J62QbRiSQ7
M7nR7yp3S+TY6AsBMXrvSxcCwofCvtwaxUuM/qTaVzPym0tQk1/Et5kdYc5whhHb
roGK66sIC7ZxdyGz0zX4CjAqF62ss72R8bb12QZMNwLTrE5mh0PI5F2tk74Mz+xu
DYFXQijshNZa1e7oxCYqwZjRLndXXx6qz848dQ067TtXW3KPxj1jOlcHQU3fCAmJ
pQLTVM9TVNgpyw/WlZpgZg1tTR1qOnPHEvHSMw4SNINOKCi2L029o7NzU35Q/BDG
lqXDlpPR27LvY80qHF1kgxxZGVTwDrF7HmjBvBTO8+AG27pM63dxfdNNuCmkf1rV
liqOPKrME8R+L2fzPfdUTdD+uwWB6QcgoykmQuEo+h7AbxDt7b4YPwc6GmZFmt1g
EqObWb77QUeTCKHWgh3QU0GhNtOyPTPp3CFeKyAFzknn9kn9V0WamGXcTRDkQ5JC
mHHtjd4IQ0UKi2Hx8q0rQWBN9azhLGcSjqzzgGBicql3okwTKhcjN5DPRA7HhU2c
qIFHfPIxuQk3m33gWduvls4zKyAopFEbXiwcvPi1Kc0lboPWGi0NWbj3GJkyuzVu
PoZYg8Jtbeskev8BqDH3rxSiQZCXurOyyEyInR1WgL+uom6Yd0X+XbLZmFem0/0b
92nx5U5tmSmh8e63H8LYITUo3T3YttNZunQTTTWzz5kDhvcUg3YFiu86LFZKnLea
YZ0C1brwg/l4cJgITdqhBKUs6E80edz+N1PLC1g68LJ9aZ/19iBGC6turKkAdZrW
pxyNVAk5ArLdtbBdhrdkIMonnCL8GXUsRVdVRTp58e2T66pSzZU00KEMnz64WpjP
W+ksmP8ISDZKKiWz2dOOFgjHl3DhpwtlhfTCWs/SeBfUFnoakUsjAsn7N0Ceffa7
RBy2/ms4PJnhUuzxXPENgs8Giu3tEP/MHxAf5hkLiEoYbPlGUyeVVqp/0go4KTdh
Xb6F92htXZkhm4ZoYAnQf263zXjGroUthBKRxWngNhB+Mwe8WTllSKp0dLpg8Hf6
gDXHtSgX4o+Tm41WHr9YNF3nL7bT2a3dShLvu8Qk0QFufipuB31fo7bImOjxrRkB
hkqX+JQVSPLqHY/gIzPMtmLWhhACPEWPBCR/CqPnm+CdSMvUdbhrIrKmMM7SgNA9
8XFIkyGzzBL0fsEkPovhU8BMrClD7yLTN7bgiXUsuOWv/QAmGdjuhSnI/QMfkajJ
gR4Opp1rmg+4AlLC3B3pTQuFONAEelpgNLY3oWVA/sBauZe0iZeCjQ0U89PiXJoK
MAkBgBB5CsgJvnkw7+NDocgEsguTw8bTuFDrAJNH53o2tt1mHqF4SQ/hqkpfFwFb
RVKnkZN6zzO5o+cEFAgzZIUiP2S856DYI+RoWcco77cgfyerkDtyEFs+NHtMEm+q
nWAI/R/BfR8fCggrnbxU2NiyYHsozxk+bl4hT2xF+a/1O2vUyv6OCGGaNNnBZAP2
aE1T2qzMjddgaVw/16cf552g38s/TOfgwEbJI/Y4SXzRmQt4IPGR+bO2EsNqz1v3
PP4WZbASbc+8QXnnHyJrYigD4kbIaDG0fCV9gncFOy6q2eAizg6Iodu4vYBE3Aa9
5y0ToYfQMoCCIGujsjpX0InHtRhKFcirI2txhuanN6Jmr4YWysv1RDQP+GcNWct9
uXzPM/7CDrJRHYQcClu6FZVHVyaesX7U7ACe7g+eCoHN7cmGIfWp4lz8ynSJPUEq
kzBhiJWG0bxHejoPT7uevhp+xwxJRI9a2XBGODPETbu8u4ghTTOc04mZPYVDxObh
fd8vCpmuGo169o/C6ZJl1K4LeB/Q6Jjh0OUtLf1dtEdE8aTQ2fvB9FbR9pmG++T2
GjQAGVy3IcWiher804iuf6ddceGkm1PBLYm6q03c6GT1l/wvQ1UdmVBT/+FtOzXz
7RvSozMFvV5u2LLPeHp1722+0v2lfPJ7xaPweXx6gGcNKFRyrVCQRNumYIMJ0h7x
chYy+QGFnIPZr3Fft0QzjHiA8KzmCPri1mcpC+DIbm41JC8ATxlMZbkKA8243x8C
9LGtD3QHzfjGb/0WPkZygwA5jzbKTtrAIhbZ+6RmDys51L1L4u5eTacfagl7lVbg
P3QBTZilO2IREoxoUPR1SIyUNTtuVkDK+DOeGrtbjNAA4GWJDw2Ck6UrRaNB+N4U
hGYarLSXVaqyI0lIOxmoZ1DEop3/sRSCZly+/Jr6XmUkr6IQ79vG2lSd/oVnoI1E
RsOCwBDfUnH/+2x+O0Ak8DfoMSZZUB8wsoz8qUDavmS8cv/l4mQr9yBigOPoYNWI
z2G6bySy9jiHCiQqR7NoqCSwFJV4Rfgm/K7lRaarWPBUm1wtEj0cQtyYRrFPnE/3
p5XEtYd6ZJvSZCFdZNo5AWt+AyUuJgM0VI7DYsNFZ0rhbWZJUo2pE3VNP5y1rmoV
9DxkIj0EUsFCE1tufnAzTRGj7CbRvAZCF0PBuvj19/F7/F9l9UW7abYJqyJFwpzj
U0OgWJvQR2/SnxY03gReSQg2tqkTygKE/em8eM5R6BC2A7vmBTrGQuADAeiYu0iS
Hfu0J0MPrKH4kY6UocRBhy15eDaLSAPezUCza1UWqku6F+Hi84RJEM0KRKTYQM00
vLLPU5QvezTgbSsTAEZ9LHuwHq/sL4mKsof4/MTt05cPZpZ2U+cyyt1umN0vgxyG
6+j2uKm7uAldnY1Pj4YeIdSFW3HdEgZpdkhglbCrtHAnByt3LAaebXenq1gIyV8x
gE8sjoNps8i/r+kBuRiB8EZQ+URzfaTn0muX9OZMT5R67t4AYG2YT2OKFtYaZeG6
smNbUIOsFD+j3voHL3NaFzCPasuwaXaopZwo/7F1jBbJ+L2B355ocNNz9K52aEbT
VH8Yj4kURvruzOYOCUiYnngOqJ4InqIuv0TyyJhBwiP2RWH0ujEQ2DHsG7x97b34
OWJjLNuEwf5cN8wFTwyadZaocy3ls2w1v7ONVge1UHSJVPIFldnmb9oIL4iTrzKJ
8NpTXdt8pItmDl+oeB3c8trw5kvbHNlrvXQJUvl7G9GwRueBza4OWsQG/KgWtWMN
s6xyRBdvYwWoPoJFTovEexWXz3HjSj+mURurUb8/LINI4UwA3gPF12h7jYjHiDeI
uO+h3Q//IE4ypJXtRJ4AChmvRwkRZR50ertM1mMPFQDMOzFgkukb/ul+/EfHXITn
PviwYwgW1NXnKVzflA9dhYq/AunHGZeyDI19T0pGUqwKEF5WffOe15jqkgMLscf/
6nyFTDDbsc2l1ruCYsokuL6LwVEoWeKDsklYraCCAcXfDiztJsSYuEBYUtY6jOes
ZV7rM6Bk0O1ZSF2ClC8y+CawXsHSt3tGycYOfdTZrwUJ+uCnfQ2TPjKojdWIt6UW
MnU5sB4+NLtfJWY+ZrW+0MBwl/K7arn2piUXKOO31z+9Jt8eioWWKhxnUxZYzoRT
y9FfPn1cTO0vrW5/MDZXKLSByszlkleu3yqoOSogL6uhQVRB30TGQOGxUXseUOK2
RvYjSot5IaVJZZzzT2ffRowTr93T35kY0pOe4w+CNSYars3YkIo/f+IL3sHfX/kz
ts3y/jGsCphe/0FLju6yE2A20iLYNs55zUCZ3W3ZYYRZ8l72nazhuiMWfM74ryrg
And02BNOiKBSsbEJCfC1eBRZrt593lupboaaqnd44Qfok9ZbIOCbLahyZOAESEOX
of4/rg3uaDj0zogKnvuzgd78DZRLBCLicRxWEaY5i5Odk3M5YrFdRb/nmjJczx4T
xMtWg8XFPNDzRatzyN43tkZcmIwbGe6viPfooR3NxFUJlRFkI19MmxAIyxqonrn2
pq+BUKMCmMXHn4GbhTSqWDCVy/v6gAVgFg6OOSz70cWEw51AZBMvkuRosLzfmO4i
PiB6+veqAzjJuT4Xe+7pEYJPgeraCYwD/p0LE3HqJpxtGianna3f2N5Bed5xnM7R
a0x4/cN6SR40vuNfHNPgoXXX3Sg6L7o+36HcmpT6g8QIDn99s4p/K27DRjWMIsMQ
JKqdZbRRNWCbVYNkofm91vhCZlPuf3rXgmysFsB3akljtVqt478htpPlxKVjHqhr
Q6bjN2Wp5Rnmt+1+7hawwGTcqNBFfdikDGcmeGYwAJLTktFxp+P6sORRHaV+uK29
wy6sr8xQWiaRaE5/Fw+prVyHdSDoeKmnnlEEzJYa+WwxyWcJHmsedSAhXMRL4Abd
VcYeCm/5smr+DA0rODAlGJuvjEDbOyN/WFzKW9CHgqAL7/NjMEpRrbIgL2aKhbLX
aQlKAMF5WjWlmIc6AuFA0t5Tl3VjUf6sDxF+e9VTuxsz3mJ/+rNWL74kECw2E6bD
Z+/ALXr9h6lvkoz9K6eLK3OcVSyt0l1Vf9bXVmc5YLQka++9m351VFaMSHsxxPe/
hMdQwqjmD2+Ma5rBQv03IRZs5uGV07W8R+xaf+zW1mb0uiSeF/ozxNQruSNDiTdX
uEazrcNCXmlk2mSTMpn6paKkvaDVWhCmrfTudNuN1lcfHZBwmz9AeiVa/t1B+v7a
jGe5IihdNB6ibrPHOnqO0NhMJljHD2wetHNtPJ/NZP9HeBKuz3Sdy/06EuMtsloy
Iwdj+4qGY75nqQM0tpgGsCk4OO35rr8l06MdoIL4Phv2Hf2P7h1DDqiblHZlp+kj
kYyWCuVxLw5/49xaIXEU7pgKBXjhMMiXcnTJqE8yHkwRa+HZaqdyafvzW5LYy4UM
3y5K6+gL+C7gBR45J2E0A9ufiyBWOXnNrLrWpU0OmmnDgvHT/ioA8ZWP5EZzOAV1
Eimad52XGhx9z6W667HPlEVt7WLaEDKOWpsFiLNg6UI2Cc0TN3eMxWWU5mr0RPOI
gjxoNaihRfzguJfhk6AK/BwLZ0WZM0ZuTwK2bYSovJl8G5fYg9vo4L232bKxh53V
yFFSCFxnnVQCioL/wZhLFOzU3KITDDGAJ4/XLzVuWn40jmJVvlsLI3IP/fN1rM9m
0lGtE7WUEsEEbQM0RbgrFlEHrSkhYlOjhcVf7E5IsN0wbY/sv8xgK5PQbmcKewY7
va0d45jyXzHOE3xJDXd6qvanGuDEb8VWu23QYKkkSwgJBRmE9ZokTEOnEWxBFft4
pyNIfR0wO9j5VaoJveIBZAUOUuczugQKmwLTwMm5TyBZ+Y900HrZhfViEC0v8gHV
y9oOXeNIA08zYjHNBmIBZvO1yGbFCvbTs73vKkWv1zJMcqbjwrGR9TzOZPrK6WsM
dFzDhKXENMBYLRj+hoqSPK897Ww/qvLWssRXhuhWyIaokw/sB6kb0gkXUWgZMGsU
KSxU2NHQkzX/z68ibAKRnwA1cYcLeFacMRdnns1GYarNk/CL3qNfSQ0YRXYRzCua
kKdikj176T/foTbaJLF0VTfvb2lZaS7MGIfpTNxbpB5vwsVHQxJXVpNDDpPLrOCM
vgG0c0ghVJbowCsazy8ux0L8MYoXFHV5ML8kLinb4odJn+KGyg2gfHj7v7/8JGo8
nSUKhOnIoIP4gwwY0nnlwpUTijrW3hot8zxqs5bwhCNSC/JBs0TdJ0o17ODW04UF
2RlswxdEEZc3taKpKuvqtCmO2w30SO5BKovDMX2WC5qlguk0fb4m6UKGxRs8tT5d
NrEuC0ihYzlr5rzF8LXww3+FrcWS1hl1Bw9dHC++Y1e5pQaELTQk7TalCMwUxIOJ
xKaAMybN7iUXy1gA08jNkrfJSMo9BbzCYa9jKh/Cm8joHQvTLgTySL2420/8XcX0
QSx0umauVLKwLYf1FS7QPddIXRMmKI4XMbco7/wiRfiHfh42s39upPuZqcAvRAvP
4GQJVvgfkGTW63g7j/HzT9SeO++/u/tjhPYXiFrCWGH20vWZurpp7x8W/rV7pFRC
6w8dzh2b3/a0GB66JGANcxbzVQXNuyYThv5EwtuRkwbI5qmc7/aX9lWrMlVLBUwD
cz5DTiZWvqZcCPqFaXExVLv1k8Z5Nbw0Lj6FCc9hq8mv1wbZ2oPuS9WgwxCt7av4
ORm81yDAXJ96cK4NDQtoN2f+CZR4446sKYwxdC3dFHCEvkof4p5LcFZwJ8guuc72
WrPa3ib81fh47GejdYEV8icwgalQhLgpY0CTgyTBAdOIvBiLodo43E/b/4nLDy4d
ZOAyEkr3Soj3DGlR2BBntqXmasUs3Bo9tReOmJo8kQl+xiT9CH15ttkFJnfcDIqF
bkYwMJRo9sWLS+EOnSSfJ1MLrkj+cWQuXn+dUKTf0kdTs8D5+DIhABDHbov5OzOn
n0cuhNjM3aNvkLAtIYrrCflEIMbstEs+0BEWVWd49ql3IJHAX+KhSNSM+j/eh/TQ
p5N8A0lFQD/eWSRc+FHZLUm+qPMSJicwTX3hZai4AXmkZXBvIeRP/tv4ndnC5kpK
0q63tPcUde/x+3wQCpiFmGvU0PCkrtuGNSlP7bpxtiH9tA9HKWh0Mn2mKiOBxnzX
Ec0FL2EnEKZ4RHu75UltAIu2kLlk2sA/N8Yu0KBamISliw9f0ZJzx858dsfcWhAh
Ss+1k9JCWNP/jYtgB6jstWO2/ftrkLMwV5noxgkPJpQb0S/2uA97FyBnrG2xhpuS
BUZdak1q9KY/VebspQMQe5qPTZD836ZU+RXBSSGmUzVxBgBZeZ5OwHrYlN/RRBrE
9TrARBFrOg2EMXjhRjdgGpVd+tBou9b7Z0tuwDGZWwrSJIt2UXeeh2Zv9ANdhK2M
SnDREzYcTK7JHtkRyJ+n/2K17wWV9WFr8CtX2mWaMSYV8R+MmvFkMkdek+Ypj1Nw
QN6ZiwkrjWLZ8z2JLg/bpP+X4gFLzDPs+m7QZpggOI/Btbfi3/d88QNn9Pm/g26G
nCPODwQLqFZa0jix+HhYgGOGb94drquOFAVoqPfeTvW+s4tATdt0A9GZJq/s56kf
v9HgD+obGJP4sfhrZGaVEH4xEh6O60fK7nVyNjKjQoapL1JRMB30a7ZawRaLG/ox
LG2tTvO+BOH0xNabuuMkHkvn1FtrBevloYcmqY1rOePQzkAblHmVMjxtgbpJBW4G
EYUP7Un0o9hMgx7rKGb34E4MlB/7OYuc2oe3rQc/GhlgLMVaguIaPv4vjj3eXLow
Z2WsbeJdAEYkxoeRC7FjLGnALonbhTfmq+HdzEcXUw3ILLDe6GDaSMivP2GVmW9R
t7gLfldh9JK17NrVhYkD/n6oE44b5Kk5lKMk5/xvvbtqzjdsx8bKa1nm9UEM7PAP
Fbs9bP3LnDskP81SgJ+g0Cd2KFWXIlypXLu8emLy6HY8GmNvZisLMh2NZDgUWvnd
UtmDd2xZRokhczs3NvgNebZVoUGLJLxJZeqaFn19N2ZNpBQo++AD0XcfALjoOgH7
C0yYmnskgbEvX0lRj7pDM2KpqnscFvLetRWFlsaElsBJW6F9Pi1YX7VyxqxEsaYq
WlQ3ylTwO6enXmY+R525Bf3JNG80lR7y8yTRH7a/YLxKMITsp8CLCi19n+sgI1mx
hcgb/JETCjzacbohg/SNXIIJqRO9SvQElLvuY2rqckIMrcb3XobPPgPwNw2Z80Kw
Ox0LWH6zXxS+zilUhL/BtyrbkKc21B4IDs9sBgqK30f0UrLWvKjWtQWdNANE+U0v
j+zpmiqJ1QQItYmD7pHG077rCllcqsAAg7pOplEO0upKLjYf+2L4+RWymVXjMoW9
Yqhb3CscXvRl6cXPJFyUkVuK5vsdYzlvGnH5MvJfPLlNSXUKSzryq0jueDa3cfP6
36GxDzF8qzG4eDinh+MB7URsSWBvJdc3gNqYEG/SjLB2ggSHrPVywOmj80IR3Kob
AIHRIzCCRPspJ4QfKxS28k54+EqrFudSuurGBgi3pp40iYmibYRg9DPlOoT8xDwz
36Df1J+RwPDp4AT2lP0zFhySHZk4WC+Evm8dBPUok+ob3zh8iz5JHAPPCyAdPnnj
1xyYkyTdJSgZ2uhZ1QgZI7tdV913sOYsraG1duNVXQ7l9GjnQrjpc4egt4nFEvNq
hoSgYcRg/tbKGVSmdkY5OXW0YnCYbauD7b0blt9MeEXehDyQwX7pEnNyeUzdDwRh
R031j//KLLvBpZ07mCvMKaWUDfk6E+QjhEbUl75mKcq/rDSEfvvKlLHFlvGFi/bF
JvlLXf/dnKMaX8HXVITKUlR+sRspzvkpcD7hnI/axUL4ChSssAhDh3EdIlGLKOn+
AW17dfKQjAOo4edBjEJJoVgTDy/kf+ofSFQ6C81k7KHHZAxc+lsh6xINgcRzMVAx
epDcX4CQ9r49yDanX6kuoRQXSFBPh5HT12Oc87wUZBySqzDEQAq8My2Fo44Ik8YT
TKDDf8xIFE+yDaa5d69n1PlbTFjThrCYKADf0naPJqlY35zLejHgFRu7pBHjJ2Ku
E56Ht73xHy0LWN9aPbe3hlN6WDg53PTLNRqC5xrt1WMk+cDa0VJD3vKRDVum4Zfk
BB6SKW3T/he+UNxcsiQavMFW5YoeMmWhNmHhAYqrBJFvi11HCKiv/0djBgkdO1jh
ojDuvU+WTB4JKtW2tQXogghV6EY1JJby1b7/qWb5ftA0spmZv/crYvpqrwzegYsc
5GNDUfSsJRsl9iHtuvHnPJuukmK6k/SD9UgrXwLNuEOQ73RqYv9hT2GzGGe+rLRt
wbrRYKeUjZ69pJDjzhrSBZQuP8lgSdrOh3dpo9wa29CCOUhmks/hOno77hIlMhxc
2rJHTCugzYn9KnIsFFrB7LFBKhrGl9IFkUrdVuGma3EObiHYVfbWnabU+/JjpZRl
sBiYVfFlfdUklCFaC5EypVhL2H+yZyzyc25qiI4VutKU5Ute7Y9oj4zuCmYiLFhN
6+EWVznHEefbx0qDj7Z5MXuIw1Ii1tQyIc7VDO/d2/Yat/gXs3YeNL93bBqU1tgx
1IWsfnHB6eIyJSgnPnoGNnkPIb5lXhWf360bEGZl7Zt9uLnZy7Ao++gwev7pbYO9
mqlVs9q/OjkDE9rGMgmfBaHSeNdLaDtX7pw/kJ691n2UxpwqWyx2n3bm1YunN3tU
NurxITApM/dQiEPE5+CmxSjbSU+MTtgDRvQsYO+Yg3xLQuR+sbzuwAsmEv/Wyn6j
ClTtAakH6mjcRcjgwzbboUhZUbvB8dnz6QqDZoUxm5we5N3kxrndogV7wXu8ou9X
mf9bPwtoh6qkc+nZ36UdckOaKbAkJxch1oyiBKx8v16izQvDS3WKR/HP8TgHWoif
jDQMHEiwNiMAF+kWIfuDMCqxrktsMlnDD0dFJnHL218kKdLMbTCrtJ2gOhJpaJBk
ivj4lr/TEBEEfg1xoNMs/ZpRdmg5ePynm5u9TvKKqcuQ6CV/e5D5L86juwQAbvsF
Z0mS9S+YE0I0CdajK7vJrtPTRrFZfuNRXMx3gvVstQSEvO66H27/ehAAj3NqXH95
AodmpgZrfI1+h5AwgS8IlfUFYMEgCrPk4B+NxL7jCPIwgvzTP9ylZjZHmHRYZpTw
v+t73HIPSJsfp1VMmyXLZEzCx+fcy50zkUxU+NMhS0BYoAIRh9S81M5hDc+9I8ca
cAspQI4pVTSojCc5OtEM+YC/C2idLuTc71n++d0qmxdpsE0voZd/Gd9HGk18DyAG
e+LK2n6MUja4XopQcjYwb3G4XqiXp+P3aZS1p9zmSmqAkyHFQB5EaRcmtB4i9wJH
ZdKiCxY7q5pzwlXfbSyHD0PCY1fvhl0rpv9+Z0lQHZeOjgxAoTx5ngPYN2US7fsr
YZHRtoOAO0H610sDNWSRas6Jt9ykNzfK0Omq4NLyq4fkj/D5q0Sc9SYAxNc+vidM
ewiRbKnUGHehPnRzD0ioQlFtoOGtm1ouq3lYAOFT3Dz97qwTTpte4uAbbGfhcPm+
NiavtWjPldYjRVos+OtB8jcFtex1S9NAKQSctSspjY0Pt2D6aehj28ZYH9PEjwYV
/qgrZhZCW4g3Tzi6+ODZ3hUpDMOgShVVx+uwY7RhJ0twEZIfwEaevHztLAU+7A1Z
TOm+a1TfaoO6Y2fmaBPMw2nIJTHrg1uviBwgjPcSWO3yIAcw++J3PeCm335od32n
FEFPuGkveaa84mdFl0RAORHjuKiZGb8Bx56Saj6jcFB5Oy5DQgNs2SSHDqrA5RjY
+2guc+8C705oOYhYX6hPrcQ9PTgeeKf7CqH5i/24/f2hfhq0LnmbC9tKbZ08jkrE
3hRrxxOiUVpzCp4gdO+HVSBtUguzjocvchpnP0qPR9M5rGYI4z3yE17SVBj+NUmy
OELiil7kGiV48gmjX2OUrdWIGFoiOZn/W14Ll2bvF4HZxlGbACQe7Hfw9HtJq69Y
C9ufdgKmGD6CwWtKFODcgmT2z1w0oaK7HIEOadoFDZIewHBgl+nhQ0dZajnr+P6z
/kmICtBCDGoqJCwq+VRMm9tNa14EguolZMWpx5r5/ER3R8vmUKvwyGFWbfHhWIVR
UyMUjHRf3FHGceQ3fzQ6OuETf6txjiYKipIzeUZBitwEQHFvRn6tAmrhpgrVcL8G
Ld564JMPxqQg/BIW/w4YQtyBSKoTcTR3Y7t69oFD1D6LsTiZbUYLLBtZXhVc7nI3
RVIBAEYQTJ8u4dJvQm8V4ExlQir+L/5haHsjzDCDxBqgGFQ5+H8keMzolhzGFpWT
s4QzxDfmQFs+1hWyVCV1k5qkn1lUE9fkGHAvLcl3tnSAgSkLauf6FGWqK9kvya9F
eZYjrc2n+rvAOQLnzvIV1P2kTgfE5625WAtU9h//f++nTgov2rUxqfeVkUXn2skB
wcgh4bRTiWFvvnwXRna9rvp5is1Yj3Sq98AsUdsW+OdCAT6nkJStAzhT0RTuAI2g
yynC7qVzDNizuHRVnhIVocASIuzWfymj2Qhsi275DVnTwVXH/zpi/eQFX+Dc5V+m
O+fHEr7HdZzDhCin1G/+pabN7hGAZGcjF/C9LscwPbYbhsEcaiyRMnmkldv0ab7i
Ndp/UDEjQnSkzKVHtmfAUFGtUZj1tQJOGF27f8Fv7QOFK6AuxFhUArqJMCZgu7w1
ue+a4FdgC5NW3TqwgpHy3tHaq/fmV2bQl4xEdkVghpWlyo7zDg9PDlgrTQZLN/b0
VzloxEga/iTFp4BLyDGVp0XWzPu86+E/ayJkxmjO8ULcEQX/wBDDerdBNvhWeyu7
99pXj2M3v/peDrY8qeAQZHO2dlJuOq7TpYEWgFdKrW4eeXHBfLdn6x/07YyaKbTX
y5pceuCOT3oQ4GbqhUhRMHphiOwIA3hhjFyNWmmb4md1OObkrEubgs+uud84zpJG
Giu9VvZl4vMtGu5FpyZ7xiAzzh0r84kLPnFXLPz4jfw+U3MF1D3WyWyANSLqgOIy
BwYLDlNS7ignmuOlvWLh/s9J86B7TVs8Z6+CEf75CT3swCmnJyJ3qUPdgGCchWYf
yEGnNKpJ0iRqg3Rr3sAQ2caFeX51YhzzfnVtW8LL4UOOovZD9zYNgHOgiy4k+pw3
zYazxVRGEm4PTiwRi/DJXPsZH5mBqlufxspmw0E3qkZZVmio5dCLTXvxQKAqbzN8
bO55JVBxoiKHdASxsSsJpntwCG0iNlrnl/s/lo7dwRU53maJV3siQp6YpbRCZQo6
bp5fmBfyNrf73ZZnnhJyLC5v+TVn5SkMbHNt2BvWaBMbLFt1IotawMt4VKAVNwkn
E3J3QrGV1XrCf7xQKej9ZnBsGBVRXImGjztHf13OJTF4Fv9LJILDnD7eKLElYBtZ
WRbjANF4NDhxksUAR/BXDUuIs9mg4XWYAZhDvWnunYi1nogmvPfZ+gRxX62l1nU7
XTfBXeOz7oxeQK9ZVPj7qXmwzQ8+pdjAF2PTSjgYEIvMEroOmO4xjXEIwRNy977v
SYeL6WuTrE5JtSA4VFOJnJc0Hdb/A4a7YNySLmGIc1+QfrJfIMF4J8pxYLSoJNhl
FHCjg1qLf0o0F1+CIXYzrRojArpNMhraaVdeJtOc8sxWHMJvKS/p7Sc2bPzsNjTM
E2IkQgQp1qxqzj3Js8gsRpmci/kATFoWd1MW2XR+khMIX2PRBPSLwljvjWm8Xtoi
BsTVv51P3SYK2CeYkII79SebztF6vXv4Qok4p6FBCfcm701lfVx9MrpMBC9sZ3gI
KuQ7NFlnxeabbH89nBifmkoyoabl/T3RYXmoG0MBSWi0m2jOXSEx1dLbxe36hTxt
cqYTRzMqxlxHpYKuo3FJUXIkuqoJKNWoL1kMw/HeO3Rawu1elK6i2bzHlGbsS866
96FHrUz3UWGv7VywrjDA9crf9VZf8xYH1h+z+FP2NMX8SGZhGdDR9rzPEYJX0CGJ
mm/x/zh/Xi7b4l7/3JxzCtIYy57NSJI/u57TSzyfChy778avqAa0kS6gmC9U2qf/
5AoNjmEwTcytAaMDp3xCQM0qncoBR4j8pgh3f1eRzUCrM6p4+oahOkKY9+rNcER1
D/hOv7d1y1MyBYhD/SirtRIuB7oRq/hy5Ko1dNP1YHsrMo9rCR4E2m1m8t5fbeEl
ZvmJACt808TAa4kc6+YECB2k8Z6lKQP2z6PhPO1Cv+SoLMAL+MZvcAA9fi/8Pi9v
EyNRhfRqRT/gMC3SMxZ98b7YpoISJ62zUQEr6wP4Oc9qz8vH3ZbZteO8/U4Q4KQS
KFkGgSaLNCLmCe7MHAzxzQFUfNEGKtuuNJ2/HaSAkbmm7IgjEWB5r4seZ0priQda
538gSq4I6ZOxUllSko1KBRbQtZT/ogLZ71h/Xc/YvL1mKHnOKBiHoxHYwAtnR3e/
NW5aAZdW+yesmK1VS+HnjcPhYwnU0lCqjeP1qGCwzKMi0qhfrgMfUkCGiRv1j1G4
zkX6Vc2R+nvYuGSLNIN9F1qgsjSSoJIOostdNpa3XgALTB8y6wUUEcSK7Culq4XJ
T1CF/Za34pi9d99tfPpm2OFT7DkSpu19NYkcAQjibdpc/p21IDEK6WE1Y5ze2Rbn
ugNRMvhP1tlXBPFjysoaL7/HtfD09qotqfui0QR3z4pptAUApNyWcw4Kb7E7vTJV
chuH5KqKWMYm+1tII87MqAd8DvH0yRs4JA7X78e8MfKWX/h5NrZ8GT54QDW63l2d
rgOxpV8Mfw62O6WyStTQE+Q4Q2c4Qd7GaNKLcOK+Um4H83fdnfHnJ2EwsfPjug4T
iJCDLoqAj1ZmYtKj4kZpzl6HPXYaUhxz0jeQJVCrZ2urguGwoJYNjH1AeEvoE93R
7olcOBKdZSLB+BkJ8cawtTWD6Sv/2EuZYOR11Mhn0MNzHfe+Gb3FdBy5niNGh9v0
97c4KNdZGpIWR/AbPGojUYB+DZIt/z93oYvCfWkN8D93ulZQjYxUdDEbs5rgDlTw
k7/y8Gwt2Zy720/DMTlZgyWHTEEe1cf3KjE3H6Cqk63dmNkkQ36Uju9iluXUv9vN
IqdTgjxXhcrT6S9mplBHDJK5Tm5vIxKXqpjLrxH5Wb54xylTX7eFp2Wl+NtMTqVS
+59nQuRCvlFmTAy5mhF/0E7Qm+YPPAkUZOORhci9fZQRmdeM0EbCb73Ps/pFlRvV
0/sXoDcSKiR7efxqBcUB+0qXoAdph29t5hiFsOyZdsXzi6WYo5zxWwxk5S8mtpV2
Z5AmydCh6alzpQhAbsVuxGbDWuBBdWhuBE813UmjX+MTqWaj05Ft0bcjwQTMigym
SVPg1fP1qe74qWJ4KklCSsGMWQOFnwhJqJaCX2tvdKSsw7V3SepJyOvGby0W28kK
UZrdIfaUaD9vXPy7u95IR2OqhkgLZLAkrf5ECIOdaudZTSW44jRbUiqvsaY02/Wb
EOeeVOZcFbbMDZenZ0VcaqpYA+MDtzx0AgX8LnA7QgCdtvwajwnFbt06JFJ8UZxH
wRLGpp3rPXIFP3rpOHktOs5XVS39tI3GH/Vn4OYUNvPLO0M+vt2WWWKtnFGQqwnr
LnUn2JWO9Iqj3AywMoGF3oEwUzcF7gTDHbaSZFDfX6f14Fw6Vy84K7EcdesFK/uO
TkYXsLpS2bpR45roLjSAwRNu7eZNnIzx865+LY5deA9GmEr8h51cucg4Ow0H0kUP
skCm2vLOj/ekn21qoiWy64j3J9OQfFhCXBpSY34nsDp8JocArf10UeT2n1s8/J47
og6JhcCVy4XCd1ZDpTqHAQnfZytGQS5M/zAehj0qPht8/FWmzsoyCn++Ib9RmtAr
aNgjqSwdKC4clBijqmOdyRv91uO1zFlNoZdaurCfPpzWvx7v4K+93iGJ97bR5dkZ
pk2lb7cpZVa97wEzEK8FDWwv9ZbAQ0Vj6EkMCnqgBatu3G780vTXiOCddWudDPbV
agvKg8nkyAydFcfSscaGoAjMvZsPppovRk0I4JV/oiDNdifo3L9m0XtBqjhR7aEX
R0AXlNyZKfnhDBgfihipqp0ATjbvTzYbaoXsvW8hbzyDV8nCIKV1PiUcjyC1bwhn
2HKy+S7Ve5u5fAuVNEQFP6b/XAWP5FiaKzC4mn0BJrdHpa/GtZoguT2GbZPVkwAd
mdVFmH0LnlD6OboLfAR+agBG7/3TaUG8NPHezFl3XdKGDLSDOmkPuYooxnd8mpFz
tK7pC4locXJUpLGElVbkI1IPdKbh4gNrBPXAMCwyzBnmdWFFMKu+3aizhxVBgWvA
mAT77lU9fWPTZwe5nUnKa+GE8lFDqVGIKPnWZFuWq1/Af4gMLt7eVIGUzd9+WIBL
c6S2qmHh6NZOm2cWCHNVxOYH1qnLRFX3XvywfC//RBmNIUJRdc0MEZGu8DIdaMjz
Uywi1RAvYXxTNCO4ctPM0IWe2C3f4RDT6v0ZZJdkzhlBX+UWXRGvZHKA2Nf309iP
NWMiG/TbHWPe5aGpmcxKWU+yO86ZLnfN+ppeMM1vJnfHkXGn/onTqaObIPDGNeC/
+W/rwvmdQ57y9aOj3CuekyLIYsk2PZ3YZwAS2spNP3Ddm0TWUW40coVtH5YLM3aW
9c7y0oS7Mtsk47Ltvf/0MDJ7dCm4DysQO0zTKF6/nk0Q16QfvQOEj0ilBRzKEx0Y
91m4YbTQ/4IQNxKYU3k9bdjehMCGfycgidCQM3zFKRG1VOHw6mGXh1i25AWlKoUt
HhNGXwJ+iAUVJxZZKE7e849CMiieTe6ZtdIafsJrDCS0vPHXH+lqdEjBpdO8mwQH
ldL5KCzevfzeOXXmcUzgFBP/FpA7FhgrEhUBXZQE1xaR19srIkoGUUejtb8uduP1
Q0Op4n3QEMVxm6hTAm3/IAO4r57dMeFRW5WVCBow3uUVrnJbvxBZoKGlYW9t+FNx
o3wWzwVawLcu5WwblsTQRgE9GeLLD/GAoeuNHXAq79+hpn4ZUe3we4X9HZTC3GJv
1k6CQzquyFmkmyoGdAiwbYBMAti/EP+dTuhP25/Y/LsKoFQBLqeFcAe7Jd00e/Eh
NiscVdaLtqq0DqVXuqDPFz44RWmLYWMKDGNp00K9Tf5bYQjwITyaNwszoEe+urry
umiasp7b5va/ZU27jfaiDR79rrQBSqhkAuSFfra5ikmp0jXetg7l63dGfxzyAFAu
ydygii9ZY08c5BpOaczqz6xutVJBjkc7BBUIwvNFRezxJ2pkkOgvnN1A/JtM1Whi
Hm0dInDVx1BqDTlU4hX8uxgSAiMH8OBh9eDTonxYxy6u7sm3hjIbgBuuPE+SDRDc
MRoI/k7fftBwRPMCm3MlEOoFExtI8zsRZB6AM41ZcwV1trMnt5nu9tta6zaYCVsW
KFeQvLBM3Rtby4VwWMXkcWxXNZ8PpWOY0qPw7N2o2ZBGUcoCWjuAoyV3PH8HZoPq
Etcyi+ElT0rGGcL6to9D2EDjwwoWgl3wWZOFCFmEWMyTO2qajmGukJxMEPx1jNwh
XxArqXDZXqLlYN4lStFYViRrSACCpfwXhbRoHF59fNWQ426uNIDlW9WWPYAXSP7H
U8NY4Txt2vidDcB/XLzLw4Q17leKsmXclli78brWJSLgGYpqOSgAQx6khrgLE2TW
VBkPLem5cA9KkwcHRgcdxqgBzlO7Z2n5OUNwqiQpKQqRLqu/hWuk+NdGshbhmltW
n6e6ccHf6A1X15B/WLEWM30rjqhRCf2fKhueT0K+vYkAnGGSxDQ1rS0P5N/zfo0Y
1zQLehieofmozKcJVFwqqsdA7WcCUqyZfSf7oyVk7eKrhbUXaWJVpgqWhkFzk9S2
HW+NFGGnIOLb2oSO7GsdW03GEkzHXnLg3xekO5OpaNqQmaktbcROQBDCXxKv7n01
T7G9hkLOYaCBfRCzEf2MjjhMXKHczZG/VJES1rYNBfkDOlNQp0k9wlE6MrjoJHOZ
CJC4y0fsi9Lia18GlbglG2YQDAdawrSHUsnIklIg8wbvzqnorDZuVi8qAdEPDczr
iTnm8y21K9XyqKPbskFOld8qsOJ5wHGwx0m9buLxGO+wNhWLcZykxxb+RyIgjH0Q
fBYR4EUogPQshnQXpn5W8XGdbI/iu83rhdtjcRcrFKD2SxOj7UHv5FpQR7JK4rct
2i19wOlxIRq+vrQBvhyegqbXjwbyla9XhcFPry9+tPsGoObep1bkuv4i7yuDUk/m
RUikFqROI91STsRDt2Pq1luSmdYtz3oj092Kh3DMvxf6TjuVt4VJbpmwVt6N2LQp
pTmr/hz2IlPcUtWQw8l22J3jLHvxJnGJAbIJK1TzO/HcoZwqq7XwYcisX4sfzLRz
/XXhhpTIhT5twfnBX7JzkxgPFeHIi3TGghD7mXCNcK9C7eiGTAmCG5Xrn4/7iPCx
4FX1FSTBAsVZ2zyh1K/lb3SHbyymV0bC1FH8cMzDZg2E9RApTnrluUPtzIN0MDvD
NVk4DiFYhIa2wsxJ5WDOGDYfXVAi9GLvNna9HDkcBsoMX4cCEV4YSNBTccqLmpEi
ekArKicSaVfEVQuJfQLEKuxDiShOi2YMQhdnuyu99+BOQE23/016oZkAWtMUptM4
wQ7XKEUR0HzzsBbq7NSvjnqVLB3IpvCLgCjsuluQ34NWeuDWJIMiMBPOH3xjllVC
Cic5l2+eCnB6YdK5Fu2Z5884flZK2aXeJ5d7zRdMzvNmWd+jdmCTK6EArjHJHmEd
xPwmLvV55ESQ0I49qkJ4fpbQvbIavSPn9D4lUoWCEF/tF5OctRky5dR4WDoc6iLZ
wvNNfHN9WngKtc45ACMFLWL7ClUfn6W0dw0mOPA5QNa0Ze7dj4nqUggNf2kIMgCf
mRvz79+OsB5sPGqzHoaY3OmWSBYiWJO0pND829kwdJ7419zLlm7rgfpyg2tYSdnl
vPGges6ekqtwUcInS26oXI7cX/9IwrUlWNsi1YShRbd1UnuDIx1yKG+WirrwftpR
3cO23fSaMgp9JmZtCRfx0loBDJDZsA2llWPPPXm+Mq5cne/9KPG/eWy7MicbaLcy
owanwRhWgU5C8gYiyfiATC9C4gXHJdNVjOfsVQM7CH2n8EUS9c2y40LjTpyELBqn
hF15YpWLh2b3QK8r5lJpJGD6YJcIpQOlZgs4nTGumG9AOc/MAWj34EhC7/WuCP4g
dbONnqa++LwchjVvrhPYIRuxI53YndBBprfetlDXdRDjhniRAUknL0vJEsty0QDY
YpevmoI/zB4nmFNrxwxVuv2w84qC2R5No15WH0/Ql5FMR6vrY6B/sPY7xG3Q8Ku6
2v7tYA81dX0uvTdFzYKturuM31PBYOonD8Z2TDCl7luDVLmP45TuR38XuzwasAnM
lQ4JaqwsjKRfJOc6CdHZMzgcNPERFOB2MVidiz+Ex6ahqWHfeMflmVyXkJd8jnGe
Xm7pc9uaaFXZ2FSrJSBkfZvb+g+uXkUNtQrvCASNkGzCEHBfTFVM3Vw3cIjHPE6d
8aqtm8gVQw8sqaigEvNKABGDDSbZm3etjj01AZ+tYPvH6lMppBOF9a/99YPi2bMF
XS9lPjz3O67/SlDfm6eZ+M7cupG29JKQz/6UxN+7Fzj1rMjA2WiWirjdJcHosM4E
9UkKrpS7VIgGeLqoQA62rJk+5m6dhan7ENkTpJki8xPxveMQaHXxynuNqV9jYN92
J5USG4GMXsdg9AS/eJc2yIQacIbodJ0PVoFsg/5Nwz2dIciJ8Eiuyof/b4CV3abw
WfTU/xCflwBSyHPsxe8y8/b5/zDjlbUL1bwjhyoPQuwnBi5GIDoceE2MAxyYksuf
tmTYHsSLQ1OY4yX/9iNPvDN69iuAzu6V3HyF5Fz0j1bzhVOm2EfrNgqflasTUvy6
XF8C5k9eB26OGseWCZIXZBRA1f5Ya+VgMP3iHuimzKsjhmkaStT81oY1rzhrN5eN
MVW92u8egS0z3QwOWrCEf1GCivBCpXseiOjGF5J8FKMoSDM7oXFhNMnj2cjpqsFl
k6FPeW2fhutkeyRy/qiNk/zDS1BOz6Mcc2wJq6AHGIm2DkFs0omAJf91Djrey4Be
Ffu5ej5TTvMLlVa0cHcB9ThK+ioOSgVyV9D6ygcHrtI2r9cf9M2JYa51W/OmwUqu
e5+3XKNWIRIRQ/KHXWfW0lq2KrCN8b9qMtyhh8HiJMnwOmiRkb8+OKBw5VBYGUuM
wC7M91wQRSp/kTqkxSO0hLwi94gRxpjVe2h/n4+cfLjEwOjuZwZZC+b7iqlbKNC7
yGhYUHfgi8fwMtCoAbVxw3pOfPD/BQIMm6HyzzxKsD8G2Tv5lhscqdiH3SFi+iwJ
xWhuo4gRbPFmOLSJdlv8yx8bnV1r59efeQAc34gZXrePgYOQ87Xtbciu1EuA9DbH
PzSoiWH9oJURsScRF/iHMnbHXcwxtDG0l3TZsArZpoBZl6mCG3mwdUcXD5ElM2tT
918+KzFkSlILfMEkXxa6dZU1kfuldzD1V+UOoAwOCimIPiVdsja+76lfvV894p9Z
DLV2OhhfiNBbvhw44XrrgTZ5RIdvgHAv3HuKFlwHe6WUP5bKNrXeHh6so9VGO4fl
xfpv49dnIDmIl0jSI6gjG9OD37Ea24roGVgdxMZfPV0to2t4aItYI78tomgwS8t+
ivnL+vTizS8p3FFvU2CGvQuJiFLNsvyMDs4eH/x6wUhzmAZaRHQBQKpxqTKu4sxO
WPEGtWpe1hXyhcccD9u/3muTOXXFIdoBN2UBtNhijtuQbVehDvREFNKZnQkVTA1e
XVrEnWP3LjKEmYu6BnZDsVqEPJx3vvvUNtoqKVLLEbLeu344ESfrjlpUJGYINKse
do6SH15HbaMtNP96890aAmFzKMOfX4ajzz3z75niwXgu570IM9wHi88AXPfkSCqF
BT2aBU67depbIHNroK9JTPfNlOVLbDONXyiX0wBuenGH1afsBlgMIhjpWASoCNPD
jH8u2ZrlFGrxYSRbrX+5aMJBD/ykXjvjUrp7JC0pmeykmJdw0ZxfDcvFoxKEQewG
xajXjcQcvQ7Gu8x6lJGz19ID21I0Mu1sY/i6FbJDC57QM7hjGuf1B6SpaHMKzo+k
qHTe4h138wP1ufGgK6A/r37FZuL6stjxNu8AzuHVXhB0/Jely4A5RopkQZa2x9mD
wwqavedUpDyShdOKjve9yN9q2aeWWpgOZIAkvR+kMmjMKbDC/QRpi5gSNRWcrnq3
Fxt3VlUN12NLfqGZtLNq5MFOaptItbbGrDBaGLi3eMqtNCcN92nMhlxLvFCFEwp+
ZceoCNMJyeJ0M37QNRHhGPg1jw+J3ZKOklM25YtLUe6rOzpWg7JjaJDV1V5Jw+rr
QiSfJIs5UdYjqmizxRBxSrZf6uZv+Q42zDOLMlGI3WPyF4phsliMzL9OdQ70OV7g
XubUTWGzWPcruIzeN/eUAa+Y3zx1B8iXhRP1/+Kd4h9O2H3qusDu59tIBtffExr7
wKOIgGMGjM77Tq1MRkLgKeVS2AqKTAmtmXwUfDZ3f4yZN8t2Utcb3l31ubxtMziG
g7ai2YOGwpHP/pmHeyrWnVecPQygbH1twgoF1a1n4Q4kvS5MD/TDHOs9r/HWTTq1
jg3XXSSyk6+LP+mIBkxhJ5uyN0ZC8w/VgBX8xd1jr+baMO1EJ2s4QZv3l2jUIHwM
QwZnV0KqQBIdLCU3OoV63ommLSs7mfJNVWbQRTvCosngd6G65zpRmk/LLZpz701m
Ezd6ULEz4/e6NNoXwxcTWqjAiVpy186tjqgeckTdfq0PDBigH5PVywM0XZ3sy9Wo
3BKwlQYCWjqteaZTqgZhL1J0rtinuk4o8zW0lxtLlwiS+2ZjqOmji7PqA3LHfv8g
iHCKtduOZi6i8rGVLW8Bo5kfKrk0Zu00j3WYOXtiJWDkDkWB7HxTmtE+jNPJjshb
yAPcEBgoIYLhZ40EuUteKjLL37T1lmakXEbnif8eLpbTEDjpITXjvEeyldF3YwwY
E1wuYbGrt3I/IB5jQv+xBjXu6NIpJ1Trf5rk9XuFji6/+dSNnI/BMXpfyhRx6RQw
WzcJ1eUQolHUwiPIBOlBjyvoS2IF4sfyZHyn5NQwlYeFSJhRa28tpw3SDx/m34gb
DWATatiIcolqxfsURa3YtmIfIurHNE/bvI9vAwOwTncXgeZV6GVB05tEr4I3u9E3
mEnVxCT7SZafdfXpM+mgd//UxVD25/kknMXtW3OtHbdpkJQ4bdmd+ydSQo+sP3+K
oZ8wpz4Nu3JR1dEvmQ6oTSUFGwfR4WJK7XTxHokxOUyqaoWvMhIykAUoRYeIAJiu
kPK26n1/Bmt01lG3LrSOkT8zTKWg+9jAE6xg+tqulTvDlMCqSqVpDw99F4WwJxdn
XcEvn4Yw8dvxWNfPeMM+jTLP0xUZtvuKZuPoUb7Jrmt5uGo1N/v/gnLYGkC6wo+N
Ndo1HTKRHYzoIDJ2RM+RFF3ovaxmxOG8rXv2KTVITderaJyvhOd0UJrXawZYVBql
9/jh6+gPaL0P80Fk2J6JqREmoVf6CSj19gnfmNGdg8imjcMKFAZxm1jxNL5QruGL
2BdP3Y68b+r6KO6WE3E55JXs/gc6P/oHjzn4sWBZpCaNXC1ERjgMXaS2XUdy4zwQ
bLTHMTyNtpomxRjTZbkEdKDlcWssEQPLNcpOSInl3Kd6llm/V+ujc+poANACQkAd
ANCWSKWwlHfNGsuTk3of/UI7jZTL/SEb0jJqeSeGx3eSdCVWxomSpJFI0p7wbQWW
wM8JXpOW7tYMDKmPCAHCcX2afg3pnvJD0RXDFSTpIkihrvd8AE/l9zFkr+eTc1VA
gGxleh5Mi1cEWTfde7QCBfBoQDSwLOxsJ3JmNIZFCayBEEY2WIzRs2XCdDC5rDuF
tmjAXfMwE01Txd3vmerRE60tGmw/wu8oxAydsMl2MBTpXFNYO9NWYqHVXHMaQLCx
lHZ9Ais20UzL6BxZQ9Knl437OhglLj9i4kU4PCD17Crewwr0Vs6f4UsYss+R5xth
9RsfGSGN7xgym2xHAJX6Z90BpkSg+w7IHOHah8wheDfzbVAtjTX0MGHoYytXvD5Z
AUsEVY7YcDnAmgkEgBrvunCNMbVptmBtoULk5OUZ62brX5K08wPTIyaOKpRtK4ic
NU0a3gFpivQaQlgQTHo+YxhQNhRghNK6ywxJSFHG578rRLBoJFeL893qXExZWWGz
Tw97VkBHtLi3LTOhltReLWGIkrbDHui1irfMd0jNaPf3W/AkaA8Qy2lln0qxXYdh
2hAA6I83JCAQlKD8yfQh0yw7lXsH7a1+y0EBPeQj30MNS4sfJ98ytcAzx3mgopgu
LS3tFcmDCZYvRn1/C991zvDRpFF8iE8TyO+LU+mO6nb62S6++zwjdra53+hwux6w
WTioRb3fNEwiqtIC2m9BcJEkarHf0eA+y49jPm2cPqvpjgnP8SotEAQ6cOIjrQkO
fKY3/FdeffeY1QOZy4mQbZhuXAIdBGtcS7tvDzgEhc1fIlZWijCiRXGwr3FJHYuE
wx3KMLIr3ClRKpJ2UqOIg+/KDXiCAeM3KOJZmMew0A3W98iZva/JoGMoumJUn5er
C91o5Egs7Fb7QYQ7CecosMzl3QlKuin22+UlmWNEMGCQ5647eU608ujPrHBU1+Hu
slPK04KOU2j7g7+NHuWXtJ2CufdNxBr1AIvO3e2Q1pBO8MkB9pqfvRtdEJChxpLX
EFefwBGsQvGH/WZA9C5c+aPKDF69DAd20AhUcVzv0dIH9WG03OeuiVJd74ZgdaFh
boFCGNZhf8IK71P4DyWSTq6rg5zJmXGxbl26bEXXS8RYdZe1F9hJep/k0Pd7mRr1
M7X1oRH0hCvIlatFitLkOiIXiQH9mHRXcqsf4GMuMI9I+fO7dv6wuyIG381KDFXS
yELpDsYOzy33/9OBqQX5jCDO3jAeZzJiJyyyyBJ0ZYjjJjFfbUwX657MfRpO57eC
vBj0s5+mZShY6DpryjFK/MrA4opD9VEJ3xPmURcyAxUbjbROG9mYI/EVDrd3+Qif
1ocebz9/QgUVo/tDc/71wZdr1xHxaZEkrcEnpHCdCIHu5HTz2N9ll1zJDVrwu113
Ho9NXI942EI+owlMgOl9ISyL+rpy55XyNcRt5Mz2IZc2A9RUZCHMToB7s8arFaaS
AIR+L/ktyyIspCldClkoL+shSnmAUdSNCwtvHhmsXg/yRg2IcMTwc/lubxGUyHqp
WTMBSHY6QuIiTtqsHV/bqJW6CvqTQ+HSSVwJ85MLNp2mH3AxhOdrWSM6f2H1+4f4
ofcHYeNvjR1ExP4sE9+dQPGD6gj4g+fr7IXUCWHvtDayub9utl9URO32VVEk5S+l
mbGKn+SxrPzE1CgJWln1JULi+IbvQt/hO2YY+ZaOUACsONYpzdJz6dGUL0zsge3q
UbP3Pk27WMjxufu9WiwCPXvyKgLHm0zfxIVMMk2HcDMK6otXl+umgfMrWvUvVLZ+
DBNl/zKfip+EIW0zPpGRN9hDCsC/9Wbl22tXvzp3g4TINdcgScvIgF9ecVEQMbOn
IAm0FBZEev5iriRwyq3UsYZ/kje6NQZ37nl7NZbKg9CjrKq9kOFEc4PI75br1PUr
LvLGAibRBFUk/qG7ZtjzI7wMJnWX0HLSIykIOf59v/7BT+sFzufRlmzqbSEfuLd5
bS1h+tjiRuG6mY1sZNoVHzYgsAsPQXCaOD5u1JmjC0o8ryjsv6MqVBYDIV7sITrO
LzW6zDrSYvx5qzFkmekX7LhZD5z+wUKTeBgrizDoOcYdlirWK/tU1ezCcf+mbGgo
z58K197cjqyjl5XAeTB9IHSy3gyixyVpP896gQ9LHPRdSiZIBcSUXYG9PJS67a9g
vj9uZU7ocYmGnjzDL4sfN4lQnEkOHTAj5iJU2FS0EksEJtxIRi3hlVKy/jzk5wy2
Bfp6RTa8qjin/VTUyI7hX7oYybnICi2SdcKoq+X6DuS4wsqvO98f1LRdHmAgwPsT
44eG4vjwLWh76v7mjLW7YX3383iwJSfpleqQELiu+b8iJpkD3TejNtS9abwSIUsg
YGQpi8K5AHZp6evncPundLH6uBojL16CEYg5CKxe7jDAcgiWLHyNQF9RTuExUvVk
DpERpfi8Ax/aYsfvVxbSvnPR7fFqGi3si5pT/XL6b1jEvbtOQAaRMD2O779cz2Fc
GJUpdPkRAEnw+HmNoM4cE5gbHnNCu54J0qfJeGgjmd6p/RxV1WMVkBRgpw770dKL
RDEU0/7fztPfaQ0pMvsxZpz+mffC/icHIFeVLpNmlNmiI+6mu1QStYKc9+XMhux9
Ra5PiyZijxvDhg/aiPY06G99NMCQj3JW+JdQMEa1MkAclUC2ackqX5wHK1PFFceM
tvJtM4kKl/2UcNF8Rkg+3i4DXaAC5pR2GG6FQsR29B+C0BXuNZUvO3jAmMpEigSa
vU9lgDbYpwHOCqOSyo5M8ELPYIJpopNudB56Ica2Ss7MSUwciVmxVQBuEOPlGPPr
VlkGB2v0JAdGhvWNkRnSjNGDkRXMH0di6bonIimlmjfBK/i7KoUIj8xGOGQgB1NR
DSw1AQa8Ge41VRlzgHuLJ0XVXRFBD8yXN0pJS0IeZUozdvDr8SRZT2+pZwyYD27I
ItUtj0yDFBlazwyfBZdB+CKM2SFc5d9yj/YlW0YAa9pyAbdb3cd8UYx0iSkm26XX
TW7v9iiFdvThSM33BNpwV9uE5d/smMZZ0ZZD7LZF/791zoUrazjnnDTp8iWnCIJs
rdSaMcDFVsb2JSoro6oTqlEW2fbxeDwkVMgdro1vr/i8copIiI66YhlLhJUEXHJB
Ekhv1sR2LJrkG1EgmPmctudF1UKpwOmLseXhvI5+O0ndy25+NGJqw+6xWsCOJ3qF
684IlbKG46vpk5UP6/FwpeCVnnzN0gdBauKWLARpzAvBc8mSBG0zKzqrNa1/5zm9
7wQo2gOg+tX9uClAY4KzqEBM4VxNP6309U3GtO+Ji+3KlH+Na3WTBjteMcJ/OnmE
hdqnahHr6LdtBazNH2JkGED5XqPR7NQokfeOxonMOyDbzsn+02yYPxrthdzqfxtp
pKsq0l80Ol9jEhHFLWSkX2ScZ1O1DVNwGs8X33akdC4SwTe3bdzvyZMdcvlpZssp
+TAgbLeGXmjlMGf1FKa7QsLE1aIYIkkUL/LUT10b42e49hXUvsuM+FLKPdTjrwrN
d/FP1Y66vrtU83ldiYj/mcFf+vEixkr0W/J1YrNBh2Qxn1W+JrfNoeWkfj+bPaaT
eoi2CljX3mZT5wSxF9QTVXbZeS/0Tosl/YG9H7yACQKDo4PN9kfwNFTrHlsfS9f0
6Q4p649RIyC2BrNFZ1BOku0I0LoykaSCGXQotAInzVHMDXA/T1cFvCLF0wcnwIxy
coYgW9+UOAYSMZDDIcwReuBNb+gMomxjhQhy+0HEBFWZeLRV2PfiJlVpTzrUPGCU
ApPkuLSUc0YbaXxwkqBjHv/D/qDn7jMQBoUSXSnFHo9TdAk084O1U3OQwQhYCgww
jQ91q5lNnp7XIA/wQ2/DBxN11rzIK5wKT5o8+vjrESH8B4vtHN9qafmrR0tXvZ+m
ObeiBXmRETJP5GqRWwocUwzAnH6FnsLBx7aAM66plJi1ZIYksbqPLBxvrj2oA17j
vZ1FQWuEpIaMhrGPkvM9Z97OgLUvGkO2MzXBruP35OINZy3C/+G547dkbIZaSSUb
H6+UNi1GIMTT5R98rHaAHLP5/vDxMjt5fpg0lK7zKFJUOK7U+eCQ1mGDp3BS0l8+
xeWJ8QZY+ilh94E4c7Mi+dXv93Bw9g43N6dX8pp4fFKOMu6m0Z7Q7gagMBb7pmg0
5NizP1rEIQEFJMFX8wWSGfJLLOBG8+SWIIMQ7mqnT/2UN8d90gBt3ooOMFhjWAFM
ZoJxNpUZqUIISGoAYY1Gy0f4cdpoB26BN6bzHRKvGgAidJk1lkWM78OEyHPQje1M
8RPiAFxvgYmZqZdeEKdEw4oV95JFb2kLVmb6DC7X1iCjyc/RZvWxbUta0pDvqtbt
AfSu8/Nt7ULY+xJVFPLJ+kcVCnBd/Uo1k6860nDMjyU2MvSRBn2CluFThBiypTY3
a6YFcsAuAwADxlv+4rAuaUfRhQshWnDw807xRQ//Z+EocOv4JAjGkDizEx5EoKso
eSZjkHrH5aUo6Cot0vvTKRnI3FiobBwrKGt7fW/CeUjJSHhe3gv/+3akt3DCAjaT
UM+aTGCNIvF0/5W72rKXtTDe5s9C2eYtjkJ25Gn9JBve/RuvD6GrT+61Bnznh16T
ZIOVxzsAt+VkdhRR2Tby/EcJ3xfms8r1LgwdVlAFQ1A2jb3I7fXywOVZco5d+Vd+
dnZGl0R7R6K/ExLdAyeTrnvUTkPpdKbUifY1qIBRo7rRZ/Ryj6/Nf2PUjIucakhv
Akhkv28wwR9X8x/JlS/pieMzJofc9WviawM6HAklkp9al/QXqyrVX0XEKt3cB0GP
SQDsjJrTsEBUsPOcj6Yb7BaWoM+0InCwltA3KU/Lp9HkVX/DS/6tobn5P+TuwmTP
1EIUecghACjcQevCOzg2DlHkx4nfhnDIq0az7pwQyBPGzzgPOFhCGV2MtV04IllM
qjxn8my6qibRvNRdYGCN66hnP0qJt4a7ZnJhXAHOLGcov2RQplmYQv68HmywlzX0
SOv18nO4oU8wild/2L6Tsd214+JP0wcMQFZ0Kc0l20Y51y5QckK8fnID3rkHIz+t
m0yYv9PnrG+OX944Pk59o7MoGXPDGHAd0YI4SqFrI6ZQjlicjXAontMuPGZ9HHp4
Kzyqg6fkDepJTjjIIn81OIAw3JKWYI+6/f3kHTwRLsUUW0Qi0zhnr6nj4Te8PwIE
t2GiMs3bHhwcZLe0xpaghudg7nUrtupcczqCfguzsqmIESdcQgRxr3yAqoTCdI7J
F2zVg7J9Tj95EpIU/Wn4q6OT8D4PYXdTOxz5Rb3I/y9sTF89f3QWItxhRtxdCpcy
7uqt9fXtTQF5pCeUxsc1HGEUNCtFKOtIkcrgwZiCYldbf2lW9sBGLPnhNGfnTGra
MUzFHy/slZmpCnxrG2pbspaPW83/eU0sB5dVxWHEoV0hRZpnrYlPhejh5gWZjjvj
EgGFCNbPTentOeoVtYzMf0WcZoNYG5bxwM2bZ8pq9VV3sSPuLMXMh1NXN1FiT05i
euRb7rQ5EE4juPsGayAK/GMgGCyFx0YohmuT/j0OFTACOACQaYtXHXiQV/mqsC0k
5RS/lQDnTNiW6lLajk5b0yEeSxTbeTvxwy0CgK5DUIqiR9wU0s9noNSBgvZbrcbV
/xT3wH3gRu2h7uBVx95Iikj3OVInx9ym6aUIksCxiGZ3wpcCNxs2KD4k+manOuGT
UaON5acaVW+PTu08nAACDiBHE86kvZ1e9HDRtR0lG5eAhgFO5wfWccSmOXfZWuX2
ntanQknrgobOPna0gfb2g6UDswlhS9Sd5kkkmfbSZFB+yVr4R3cmahOAxYV2Qghe
oWGSUEJ9RQlCtcwNLihocpSPsqJnHtLKzP3az66sW5Ji1uZEfg01ZzWYVOzpoXmD
dY5feIPWCfRzP9oybbXOneWJ1AGA47TwrbRCN8kvBS2LdW7FdQvHRkqD3jZJm0UC
A6rLJhIILI3XCin6TqObbdZmUeKi+BOFXc2l8CTbCWjlSXVl27NEcVl/8TfEGig5
yzwhInGjC8wQf8pyQkdTnbJPNNjgOzxl/QD5EfW/BxZ34CC3mav7gKbzXXS2EFVP
zI2vVm3kN2nNYlTXaqrJc7hLH564AcNCel1ohh4qh90UBLdUCW3RF44l3Oi8zVoj
stM6e6f6VCohXK4adp5/QP4twxRPbYbzmcWRtOJoVOEGY2ZZZ/lEHAu0mWeAtYKN
pDVUVOX0q3pfNHQG0zmGw0HUCIjA/AsqEz8Ly9H8wpkC6TMHN35UV4AyNhKSp+Lu
HvTW5t8HwcHRRax5hFCX8nYyVnLbitD5H+Lyd3YZ4nA/tgCy2AhqIBzJB7rsPbCI
tlUCEDHw1a7CQR2rQJfk/RYHSXTAy1dRf0DjDmtKpZBZ/37D+TtlKRb1/+CIevK1
tbiibBPUORGxYxxBaZaHkBT9Qm/x5TF9sBZ/VIK+EwY6uo8xhqBbTT7VtxYQ96mk
s/aCNN1b5j47VLVqYEr74mQHkluo7YfUzp+2e/aN3uAyW8f36jLRZN1FCqf76z/d
q0oXOb0kunjtdFR9J+0BPjqS5eVDXZjISzxMZIL3DstetkF65A09V1v3Pf/EdAT/
gNeCzBEE0y40jEevaKh03QBueYs4J9xkKL4asToZQLM/48JABCLSQQfxGJ2EPRX6
N40mnZGpzqy547RaPNzV/CCIAVu71mCGP3yYO5viPzbL5wlbXxku+L1q02whigEE
a5db4G9igXk+62PunPMnlHkKmKbFxLPbChkZ/0iFC2K7e3oDhig2p6rciNIOKFtk
Hlx7twEHxZk/PAnMXe+iGSVuRi7qDmcSfFgGiRjZLuutmV88mkL+ro1JcEGLsdV2
JsOYmMeO4hObgI6ROhJXnTXI9Ul9E5I7qr9vLU8o/6Bf9Ma7FMakxZsq+vjvjlRn
SYhtbdulUMP8l6oImVtuwqLvqHEv81GAHd+tzGAvIZpuE6KqvktCziKzfdmHZTxX
gxW56iJjci4hurH7/+j/Tbwdy1Rz33cfp4jcg68R46erAE5iIwknMKqJ5JWDdxrT
Mg7nt2LtubhchGalsl6uSLOqw0/8gSXJKeG3UAvbigjOOl/xRP2p52SZ1QqIkRAx
REdpazDhMst+0c4SAFRIdEcPE7uoQIxyzalclM1g5qjnSrnzrNX/8VlFnRpABasX
SdeNMcyHwSbo4rMMAjyEWTMH6M/n5wR9JVtRZDs/rKZjDBhcJUD4zfMcOjroSFvN
2zKu1KomcjPDjz6IvI9clktus9zYKfITznYcMPBchjkRTItP6QiXg6ON+vy8Bufv
fPDuzruCQBIKsvXyvd+coIMD9NW9LOh/erUqBz9i2ZFUKXG3IzDK4Xob+soPRy9a
mUtWtYxS29UBahnjdquuZkk2LHWemsS2p8Dy+5UUYUWYRQL1Pc5NfW9+x/qyGJ4s
YNoZhFyGYB3Tg0EEoJ/mJt/QWue4jgY5w/3iuHVaLT8f1rjH7urkvP2wArjTqo/9
kKcovsSji2PmjUp8Og15YMLcNZHwDFJ8Q8SSQW23TJfd4+MrR6nvGJUTzIWLu4QH
PkTgsS4oap2Ybs7f2Z2Epjuv2DC734vbL0Zy+6c73t0cZvQtKCwzbYAz/Z9ZFwzr
ydnpP10aGr7znHgjzP3PrH8QU84d8Dcjpgg5kehgbPAU6or8MMl+e7C/Qo+XCAPR
NhKGrASh3u2//K5ISZiUGRtDMhdbB8Ed4PTTCOGbNeRBAVwa/e6Xd8XMe7+vAaa7
PGvkpUYkHdFEdVxje/fVIZh6YGhCgKv1qU8cW0+mxH4BuOZamexXmzqsMbp0SNQz
9M7ExsArRgzcJYmUlyxxBDE3vEce2iUZ5Gm0iJRPHe7QENMZbQGwH4sXjXV2w1+p
y6Wn5JvsienAYEeMeWC2K4WMeCS/nq7J/dJ6kRuaKMfj/zXXLCnDnxHr2CU+Zmob
ugDzbt52waI7q4cTQxD2S4t+bTd3eR31aifWcJmlfJuRLOOTaKD9Wb9XxzI5Wfoe
yoJtGjBaAwY1YeSErDb0LCUHajzPuGfLszXKrcLDRZK0DZHYVMxOOVCPPYcxistT
oNRWl2mazYtTuuw543X5ampj/oibJzd+X0F9LwC3Osn1sUQGMKZHjKGtZ4wpW2GY
dfjAgGAMkA9b6MU6oHedcPdUBlcO6hm4f4luQNzk/uM4xEayVgctUmrtdgHhcj93
3j2SRoFcPyB+TvvzTWzB0PthDHMSHr+zdIydBiTzRu7wcyI2zT1aY5APIupsblaL
mByXheAACVKuOBK7V15GPfZv+iN5/26j/MVZMeBi8sa/JVTAMtWCVew4gtClPhx3
yroUUwQJbMohF794jDKrJmNwkr61+GMSE23ZX0s3KDhYlLLLc2SFRRIJyM5S55zu
N29RHlwBdrqhN/HCg767Wo5qYa/l3etIjjnC5QG7pd0V35S+T0VkbhBajLPiVEtv
KrKwidZ++ESxDIeOqlQg0V/aDwEHCGN3kjZSqZr+qnfzptZGbl3wnKoATEHepHf6
uDoCtksAoLGAr9psXJVCNkJi2+FtcyQGyv3cKcwJc0dI269dtKhd3l/hgcfErhKt
3htj8qwWp41TkidH/PGR8TMG5IyXXk/580fqZ3xuaV0j3ABMOZ3JBLVAq7pHjOV0
Rbg9sj2jfITp4mYTe+1R68tNmtXcqdJkTfCbTuXPbgoqpVzvbKzYvpi/amV+fk6g
b36NpoS0GcMz+POwwdjDBjQUP3LgzG85r/izJbW/HW3/4plrQ11g2TlvwfLSAxU/
GMIWnANGa0pwkd1Ux/TkfP4FWSy5ZbqN5kvXsa6GD5XTA0yOVPaTGMI/fcNriZow
w20zKkDN+RSpkMC9/neqtKYBhnoisMAyw1V7xeJgSOVGTEW7j1XBDcr2mWwH3DfW
IRJCwCmJwlZ7PmDYmiooZrxSIE5FwcdqRYyGkdGf0f2vKqY4KJWHFiBUf0Tx2mEa
4i3RfFOigaZCsov7Fsthg/nOIsuCfnuzOfr1SSbJ1/DAr86xADcdvyiDYDUQPOsS
fbAmSBpQrIIGKiLwfhksKNn+cAi51xA3j67UIq0Uwl7bLb82JFZR49AprOpe1eha
8hr/JpFh+eY5099QMf4cei+pPMN6lDhyEJeuHh/NWQgBVW4vw3BIxpGi+bIT1Doy
IOJS1iAZBE1FRFDaurFKz85XJFLa2szeI6BZ+xT5+4oDLLy7JZqavHPANMORqRM4
0mTn2obgG0Z6BYl50j1Lx8o/1UWe55m8jd9gf5XIm9cOiJJEdUJsp4ceXFz7i0KU
Tih45eqideaMA6QP6tRsVDxh3GB0bgaVR819lvf12wUaiHeiu79wsXl+gEB0hiI8
/YibqXL1ySqo2N0fs+h6oTfW/lXjfe2DrUFMdte6Ev/XAPYaZIh/fO4UIOFBK9VN
5QCzEUMBEXJZ20fmhqroRRMUdNddIBv0HRGMg/a8Hk7+4vOePv8LtorjjhQKEh1M
YGFSDbRqb9CfQFEtXy/y88xNWwqHFodS3EqviNzczBcQdeMgi/rhr9GhHQN65/Is
SnJtYv8rYBlZqgVnJdBvLGk4OfltPLSeCDi8LSKVymFwISOCqlkITA5qTHKM/I73
Zgs/jyPL4Pxf306tiyqvyyTxjpnPTvYv6vbPaBD35I77UuULpwvoCoPecDfnx5c1
CFlk2ev4e+zFLNGX4vwsUL5lSoYOjLOaS8hmzHhAwlhnTUDqkyALnVv8IvWarGXM
DtyOIXDltHsjccoAgaPy5w7Icu8NL/+/eC5reBKkV+sJUDIh9pdI+oGRXsRH9spv
az0vUvPPgWAaxormpIFdFjH3J5rWPkdXYRRS/ERjSomeYar8mEp/AnRU12/1PMfS
nORPV+Cm2yZ4PtJ00PMGHMuvbwSbx9A2JGZurNuRYMxKTGwIDe+Cz39C7FWyZTrC
/hOCSdLCIiycCIzlbsIOJ37zYr+JNsjWCr3n3LXHXKpS6eO/MwG/1bxlsMkUap4S
/4M379Nv/mfMxme1Y3TWrCS9gxlmrAm5t0T4a+J5SuTmGB+efYBAaERQmME1LQz2
C0mll3z3LJl3Ffs4b6kgd/IZi8UQkBC+VY4PXbo+J0deapBNPlvoRU8jbimzNUuj
LIPBEnW6pwqL/0kYtrYjLAAkHBwn4USRSuIgldHwxrQMZ3agilwEDZGNN9ZAomqE
y6hvMOdGzDWrv2mEYHtTE9tSjdPGyFAj6oh6M2vlo50SNSEy4dD8fJ//KFLFC36E
`pragma protect end_protected
