// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:39:02 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
age6j7n3nc5bvFzRq6+fd4COvlENkjgKYtJynm6xU0M0dm5Nacnmw4Ik4RXw2d5k
5Exq1UmCVrO3sXWxTqEyGVGyCRHA8ksAHKj9uyCMnAPjHW1rEesrKlPl4Nue7219
IuLk1z58Nh1OETFFMkXI4EFZfQnRynHjcWNSiBkQArU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 5584)
NkqXzlWa+gKtwG31DeDb70axov25+1nAW7+l1ljgIbWdkfozQLW825xfhD18vOZB
DVsw8Zt5K+OHKkctFPdd3DkWNa8Pk9i7Q40zyMA/mcVDObZIJX4gxzwxJZU4SSJ9
SzkxMs7ZIjGHuKWzHeKERor9cSke/m+fVXch53K3cwogPzAzfNH1gbbm+GVoqMA4
yMP4wRo/xLjxsrNCQd6BNxa4YopQEVtw2rQH44+YSc0PrZ+mzCkKO/5078G3lC63
6tru86v9wWOnpX/nneTIKRQJgyqHsaUCtNdnocns5xysvJFbF5lQMc9jxHjz1f5F
Fyo5JoQ1G2acJPdLyRLmZL7ye6v66uZJLGGq+ULOkdFqH9h7daeXmceUIuuph84A
365cDCjS5vPutH6hu53paULGsZusxLQY+clZClpZ9AfUn1aaaHutjraNLzFu6IQB
UBlT5rj7Rg8WKKTJac+nqR+GR+oGFL1t/JWKBTN8iuX/KaQIXIvLuLiVoCYpqeq3
EShKc0tJKCBVMfwdkaCsM4cEH2xyy9CYGAbyLVZMWzuYCDwMG7dolOquIr5OjfYw
HRj05pzK8EtJvQOFSsbOf3oqcD+nzFCPMIdmOSati2PMozqqJalpNNU+mBIDgcbl
EGHTGIaeurWn+P7drOdZ4pVOzcAORfpPTgUCyMxzi0Ues8YHn5r5s+LCHH6Co1Rk
3BF0Zf47bR08l3TvOH/roM1gIzCfe6rtYxflN4Fwlbq7xB0+TdpgbpXNjnE7Kfc2
LcdrvdH2TQ6kGJaZoODuBEntcQE3qwjcZP4rGLwMZlHR8XUKvFdYOtK3tZflKOX+
mC2pDZT9jmfsKvlOtHFVNXq5L+TckXY41y6NUDFRampDGNmIJGtSgVM9bNqa4ux7
XIPvFHmPSxkavXgm+VcRo0qqjnL6IcMkiK7du2YYSPFzQTiQyCgtIdGa51VGWpQI
4mgau2sLZHNO5No3kGPR2RspDP+eCx9KdGLjkuqmsP735D2dJD0R8vorgkzY8q6e
8SIx2h7b+eWFuyvdAfLkOJkSx2pSiKkQ+q5nUc5angol02Nmz5STS94HWOntvo0H
LqldqxT4QN+7m/HjnbTlUNA7JmSFvXaektB6EwkFLaX8Eh/LPtrgzt/yVZkuNG9J
qRcaQWgpc507Y/AcJyJoR11LfEzM0HFJylsvLyiUPYh4RP76sEwN1s3vbhV05LsH
gRnjBd33aLoyETk6xTC5LIlz2J8jXfG9Hkiy+U/OqdSr7tR9f5AMxDqTXNfqCBlE
Vx5DkiIoVAE6R3tNCGu7N5CipW+ObelJBOS9+HTmskSvr4tGn/6glwESmc+FOeuU
TsgvSTQXuQgCRJIla4xUM734MP5INC8libhFl9/jJlTPvNUSQ5UxcUZTk9+LbDG8
krUgUu03Txw//jHz1/7GqVHhaMcHx8YYK3ZqQBt1cqfrul6ZVKASdFggD1xK2xDo
h3FiSowlUHxV6V50Yhz9VPEJEkUwvu/d7tsEKdVvbK/L9NHdskDs1dgIlMg1Sgsd
MTtOew9GCB4RBbXVsdrJ0l+hb4DIpi9OnRLV42XxUpl/j+J1YPobUJ0gVecdbBKZ
E/+bguLTBtC+uNrc9jIDF5WCk4/m7+Y9X/HjvLsgS7Io/a2xAxG8ZbCR+/ELtw7z
8ClYIWzRsLhd6HLCOieZytfvGOMA26PJhGlOe5UaPk0bmt2C37SHsJxHeBOY0duy
OPkqjltJFNII6AAAESa43zAQMZSIubbWc2JKGqlgb1GpxXreTsXmKuynnpa5Xpsf
W6OkvV0JdHspRThg0k7EjRqYXiJmVljjuSuAC3h79DrFtlllk36DEUqffgxwUrJk
KknjDEl/JWabFi1G1bxYO5ijaLJcsJNMWWt5NjlhT55xnfkbdHG/ZVi/p7RfBsu5
P8MEGoPsCP+MPQHtNhJPgXas6tlUD1uslDPI5icQf2NUG6x9BuUHeGZ4SouOBoD5
LxBoGGta7s5et9S2doYDbd/VDI7Wh7tnlks8RzmC5QL5ZfGnAN93DWmFNdtelo8m
3IfkLT3Wh1m5JCemFNlY2Y+nugai11ro13u/mjUo5aaxjUPTrg78O4J+NzxT7x9B
tAvAolpNtJctmT0yQDlJDWxFSzjwTDtf6ST5Bi6kokov4Q0k9Acs0nZgfJUCeIvr
pTxnFQyjRbGuiw5adEszMkobWM43wII1p/T8Fwv0mVT0mZI7uZ0slKLK/LLZUCCu
82zOYusIhHOSq3oynL5T3w59umM8LqIqjhi2USU3zATEZOeI1oCmAg6toS5gqvX2
pAGl0sjpKBrx4JhiNo6ExUHo7COO3bEHNrnGbn7iJme1LmvMvpF4igngczWWbi2e
+PGE6dLAwgm7us8CMVvVDS5TxBI5NxVohtMIPkGKvbnn6cSjU55YpLSWNjyo6n1a
BtrJCr0TZDuyIGfwrKI4i4qlbALAjjMAKwTSPxaJMapqMKe93DWb8QO60SuA64tQ
hJd36orGje2vnXmCk947RMOBRlCmvKwWnJEl42hkS7pCBcWna+oLqHM7KBRkkSxw
RUxyCVQ/khXh0DT6d5KkElYr/O/weOhXteZBzpB/Mj9u3ua5dL42CTcRTT7BcEXk
KGhzqInk54TF0aJmZ3oQaJJpVeOG3OoV/VDzJ00qz2yKgqzRSY33QxHuGSGUg424
GD8Yp/8AIHZump5TLklIdlfL2ryCP8ubt1EvcZqSlUnl5vmpc+A4xU5xhV5JYua3
pyiGiaRNGtjjC8yRsT++V/r3zgQFFRo6unbVac4IaeCP1qtKOTifo4AExJz2iGcK
2ZARIt7rD7aJfCY+QYGnNvNeU1pbR0BV5POFcqsP+NVGMoFIT2H1qOIWlrr3LeHL
v2Rmb4LwPTYY9DVrtUwlHa6igS6Y+NNdcFOw02DzYx0c98B5VVyAhBfX27e3OpTC
XuUUZ0NN7KOC+csghnqQmWORyP4M7Acj6XRYwZBSrMjDsb9hJMGZKEkzj+t2y+Zb
t62NwRdNWUOjTxG3OmwLPJiXFHBLRHw/FnhUgF5NKlOEWus8Unbon2/61eK/Q6jg
zK87fVtvr98jMaYZ+KCdGwR2IEQm78GTmkdm7IkirHddeODvREZ3ml3XMZe43HIR
EsBmwd5ut6l7mL13n6GDot4zz3o8/gxd5NbB82tGHhGEDTSmC+SAYC7ERsmENBt/
UegpNZ1vVDIlG106juvu8xYzsMcJuAavTITtzJdfkg3gvvMFui+8rcdY/EE4Gk8n
mNBXcUEhhnKCpMj/tA5SdP7C1CiM/mdNeW0WgmBId6oOoNdBl0lGIv3BMYgEo7pk
G0dARU7chXYiHXDapiaGAp7WZdkEaUpj32tUqmFJ2S+aNippgfYVItpxxI+72RU3
bKGaC4+/jvRoR5ekUBBI3gCMzYUzG96AB3F05Ml05zp3XqT8xUmOvCskgX4PfQox
emSHuckBgJ8obnJsYrmJku1IAs2UPi/HfHlQeb/T8zWkVfHJ8u4LhvGI0PtFXumK
iOwjC21jSHdX26I2gfeY+ZHcJT3BEXNLp5hTAyQGpkBMjA3L+UYWGim6QSsEnPiJ
HOWJ6dxBgUKySsIrx3eECKPFuSypP9oRQN/MiPnxgc1zELuIK87jCTWIZqAeS5kq
Fccy+iLJzmKnDKPxU6faaV3clZ7PAtiMbt/GEnXUBajIL23dsBoGH6UlO52z0btX
XvIRLv4JnPed4SnyrhMrqdf7ZwOFn+l6PImcbg6EUXmOjwxCDo8FzZCxskPHZ3Mz
1aW2Z/KEr0zGDrl1li3gpSubkAb8T6IahNsTC8YBN3BpqYA+Z23KsB3DhruqNgDf
71nXaaLrIUnjpXyGij2QQ+Of9XpJ53RxE5VIIykIzz69FyOGUh2n3A4Lkue20ZBO
o3d6BiJu3XYT0ez7/ggQnl8i1rYuvzXHPfViauoytvGpLfMBLeiZBxK1tkB4QGWh
8coU/zD7rd4TociU5y7+omeYT4igDmUwYbAtYQHz6hRqs3GtE2Oj/+/0/o+E3qp7
rsYCRXC3D4WeZppcgxi7G8/2YphMcL/d6TlxyzGpjHWsINn6ZqSeJ4kLguGo7ean
JhbjwzWVrV02rA7Lw39YjnHmSCPm4cklh46C4tRwSf/lhNA6cxmUXgN5/O0UpMbT
lrn2MWmbR7dOYBSjfmAl2o4ikPDjRjLoaN3+v7PV+wgnZAlB+bQKH33oXzeF90CM
sRizuc/21z6sgdfhBTPkAnhaUzgcUmjPmlRcmHl03Ccnciy2rTHuW537iWtRb0Zi
c5q2SBRDTwR7/4TY9dY0fe2scPlOR9Z3X8fZYXzHrn3rmWarB+fmCV66jgmFMO6O
yUHIlJIotx2oQBwms3om6u9lsIaesGhWg9YdKTrwR7F5F4sN5ME6+Mte1czoMAl2
ZXbpQUcsT3sy9kkD8xQzGL8ROT7PZcTl56iAEnB3hhMdTHduqTvkaw24BuQQWCeA
x5K7Gn9HGjvMTt93LJPjSZ4saScP8uAFC3b89LCFpmWNQG9p4fepGhP1qrE2VTzT
YKHVr4Ev3MfgdyrXPOC/t8rI1iAlSFwmKaiG9xmW/aO4wDXwaoJ8SZqRQq/6BgE9
lGmJja5hdQlmuVYiYCJxAUeeHqkKhQHlMisCkElxqWQk8lzoSTXgmTHqiu7p9X29
pSAEEl/xMzeHIvBOBv7zz5VzFWnLxhp1JTGe3aIQ/dY5gEGSb6OHH3w8yh40nXZc
VJsKbIx7B0EvwOSh3lv+OGUTJBwUFvIbYhH5Q/BMUsam/YlCl2nL1+IVNZHiSspv
QQbKlKSuR9R12mIh3DuvDqO1wpn1GWtAcc8nhIfo9WOirTXO0NO0nATKKtIN4ZAq
aErDMxhIvi/UMDmT5xmUVNRM2twlzK6o5cFQusPNX3Ild7xDN56s6xQVN9C24muZ
yH24NzeVG3zf+zECNXPwOJ/kEFjiuQ80HFB3jYAoAPqToCT16SCSb1weUBoPwVcY
o1hX4LsUiopDDy3LpfT5vyxi3HwCAHARY39U9qa91a0KKyoBDnyR43oRAvHn9x2b
SjVlC9QRdkWHW+zeTwHW5rB6FlSSAcTfxkmzPBX3MX8z1cE/2T4Dok/E75uGDRay
0hNlbfQlF6UM8R4OoMjgNlvBK9cbRvyv4FqWYL43KXRtDUjIcbR9ylDKBlkadjgf
HhsAeqXhBxV2EP5VP/0gZ6xp8Z3kZLX5TPInFZWqR0jYd6PaTTTzCGzvLcTWyhW2
TIZYpYaWVefTAobZ9zJEqClJ+m8uHDMGGWfiQmzwUqN3w//HJ/Vtni7cEUxcxp5V
VDKUemTHLveg/LN1ZEZWhWmiXcgLcGez3jX/AWWdS8/bkDPRiQHRasGEw1ZuOH/N
o6N9ETj0GJOzpO13nqG7EMTaQiNBrxX1pUcHSmuFV9TynfanovGyoFo7d2jafq85
dRTHDQCWNl3AgoW8uKYyJwRqvUTkaY9FJ9cQr1SPEju4va02NGdwDJFcZvoIbQhV
FJRa0ORkgE4GxVQrrnvVywkitsOJqTiVN+beSb2JP+D60uee2WbxzOwlVhQs0d93
61W6WIlVzY6hqBF6PAxbGSCoB2ve6bepvJqYp99in5msCzfx2rz+C5CsCVniatEz
dN51bt/sAgo2hOLlG9d9RX97tJjX5lp3NbzX9ramx8SS5KRA7QzAxAGrE9Hjh/KF
RO04CQVyL0t4A0ZOtKchS9UwfAj2CHAUbHa+awKeKYCWctj4jnXA4hdcmxFtS1+g
eEMEZocXrf3AqIb8xD6bjt6XqszgY7X6CU1EnqsmgsgIF8QEVjv6o7Fqe+niJ1WD
ZVm/DNnTVvi3iV4zWivtCG6yqgc8He3NR5N8SSallp9LeK8ixDAOZxUzbPaoyDSe
aZikq+p1Cso4Kee6YJfDXDMK1db/VySLkLfNgckw6oQnph7bZNH7hsnHfjLtng2C
D2Glmv+FLmCeSJWAocdPZj3Ly1L0ClHhyVy/AICB+DLCkj+WXAOSFCevpyiid30F
P3mEsycROB0S6aa9NWCQO4lUeoeESG/+CrCZkxCPN9uf5Ljt0tBziHu1APfeauD9
tEMrxZrPtvYgt7nCygQ5kbxWRJrf/KpHutW2BSlE2qw7hlOEtWasjhXMI1UWW/Mb
vv1EgCaX0bKIstWGz1r4+rv2b3r/aFxfFzPIhfYgoyiW3F3oMfXLFauSjdrslntu
E4f/Ofv0T0sIve/ki29InOtCy5zg4oqcH9HX/nJZ8LlkPI7k485I5JCzacC7g34d
/ZRPfYqf/e+Nu4WKEAGyddd+r6Urj6qb1jK2wkzsKA8WA454Lmt3gx5e2OXemYlv
pPJMMCFvUHNnqVg9S4OAjKUdaYQ6kAeH3hDieURpcq+p0kNd05t0oJ3ZIoQWvzro
31dGRfhi44z/FOYP1V0bBx3rYBiyaq74Au3CAWrq4MZiEb5c/vOQyLavYS7jTk/L
Cyck6FVrev9z9sx6OJpPuXl1G3KomYHqgO+3joLyupeX8nMZND9fINmZpD5LSm6A
U2HZcd7rIB5ScRNFX+XDtdMeFxYllmcmTyDWAwkEt3E7Teo6QvySEuHFsniglowC
AFI0OmeCfdNwZ6+I1UpUuN58rc2Kh8YN9Rxaf30xbcDuD+AtPdtlZh8lO0L7NPSZ
1qWpxQCmQp3pSuVUIvbZ8BCf1h835Qpq01dZsZq7Ntg3dSXjj1UgrNDP09MK+Up7
BZITL7pqERC7pFadEbuyh5Sm6Twf3mOsRi2G6EZHDd/SYjc+RNhEyQAsAKH3gryz
GOOMDvFbb0jVDB5mcxF4D2oWJT1pGTWdd4vxTgi47zY0wmXT9vMaP3fyolPsRzeP
7VpUkclUtdYYTvS3vIgKMxcevNoSGmOXJtlTDXfbih17pq4H4mXJMMrSjbdY0MVT
JX31qeO4TEcpdiVLK71sLQHpwja8EwfLyap4f01h54/StDF9FmlgC9kIHISr0pkn
HGqPIH028HnI8kC4THPDKOJMRxS5XMY4wT/x5EIWFTRiEYzJDOR87vblZRqql3gz
DrfQCn/ChI7uuBBbzT5aS4RBEHvFvPyzpeM/DR/z1OuC2Cc0NKaCemNpxJZjr0Si
EGrrYvFMGhloh9BjkS+U8u1wZTCCWVMn3n8VLtf3nvcZX8/WX7mJgIbdVqDmiyOF
gL2HnPm78SmGiUUHkebRvP2Ku5NBTJkG5Qzf5V0XPIXa3KQeXjMkUCNvThfVwc8O
LHKKm0GJfcbRx052A2vxbg10uk50O7svxkHgdXIYq5ZL0hWLfKXe545oQW/90MRj
PdkbpZRIfUv1sM/Gi9JQPsDrOt0vwe9vy+k8tiUbQSNt2PdjV7gE/IS0EAZ7m4V3
lG0yI43BLwoUWEIn66PqVi2wx4aQDgA05cQr69id9vdQvdgYYL//rwQozYJUw4aM
hfYYKd//3AkDa2a2RjMiaQ==
`pragma protect end_protected
