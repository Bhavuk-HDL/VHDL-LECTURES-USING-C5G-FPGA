// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:43:28 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OUgC/5gjW5FjFyInm5ocju/LdyPZ5vQAaUvJEWrOETGRWYfJsgaXwDkvz148UkAN
Ot+/EIL6gBwah2U8JUGGTMGL3uy1olqjEQjzraPE7I5aQ+9/634yVMcEmo7/J3Zh
wVrC2q7XrTcwu/VFI0f2VsbcS5cKI/5OMCccSYyKv9g=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 13840)
JwlIc2q3b3kzcJQYH67EdwtHfBg8j5EznvKUBfSdutZBwwsaZUaVn+E52cBhlWMH
TAwJr0YYJryW/3HRr4Ko2j/SAgSWVwZ61aG0o+81IMP3430iTSC24dEP+cQNjsC7
L9Eu1z7cTX7tGhx41jA++q71pRXFSJA76SKf4T/Blz7qRFkxc6s5XZ3jc5AoD/XX
7WUZVWGhgITzfV5Q+Zz3fLYDPE9EDya0AsqkVr2Z7/zpj28+NJkj7knw+p14q0np
VoXG7dlvxCfCJjN1tiTEcmOb4YD66jgpWVZS09bgHk4cIAx/pbMP79w4NlUK27Xb
XOxtVnqmU5XgxRAG7BLSp3h2Htaxx89+Zb6RGTgI/4MmPP//q0GGoq263C3k49wU
Dw1wjkwxqFR+YVX87b3s3o2xmyDCKMfGxF6cB+s1FcHZE2CKVLaIzP7vK+NirOr+
wjBF15u6xYGc6+5oKOY5K6DNJrC0+3AQlLah2ddFS4wmCpdfdzy0NAmy6qR8UHO6
+pknhfs/JecVNKQLJcBNN1CKjl9TFNGDa7razsgpk9NeTKs+aD9zesj9OtS5CUEp
Kyi2XYhgLteGbROux0tvTRbfvdN5kCI8aHgHsUylzbH5R6JgWv0YvS3eoHfwiqFO
Pj3xkKFB1oxRKOhmSWTfw68dGoj72YslS/jm7WgMfOGTBeE56GwTwTP0IGhMtENd
G2j7DY0nwCp0jMwCz6UMG3MpY4Lk2wH7v1fJ942dOekFOq3adLrk+xnaMjC5A5Ay
1QwMVuWIEvYzfb5CvsRktwBb7Do2nERkLFg2xKT+us366JZMYP4h+t35kJ/4GMXr
zQGQwfWB3B17LygMsGEAvMx4kvCTU26dKqgukM7MSiuziT0/5eOcsCdysJPqubsG
7GrCPhp50Ppj2ENlT4Mg+CuihLaZWyYx+Y8No5rl4kS6oIxRB59HJAb2WKM2LWTc
cmfi+M928pt7qAVPPC+5Wllh5r0MQjVqWVg9Vg1mE7NM0+IIAcWXDiYHDe1ehCsj
fR7PgeS4nP/Ulscr74xAaPCf+G17epYHQOMDaXcWsx59pKySvKnf6dtS/zq5HYAO
xAAX0F2ZZ0dmQMenFFQJZ+RZ2YDoEymnQzM5QIRW/pQM7y7gRF+9jd6INkmKuGhY
TUPcypQCQPDseQFznmOQ47hbDQesuFwVU2UU/fRT3EBvIVAJurSiL2ygYx0eI+DE
K+McflPZxQxzjoi0ndBRW5G+aUEGWOXLAKbLzDUnjTKrydXyCXXDVS0wXks4BkY6
YZFZ7bm2PeROnkJcmLk6Md2YsXr0y+p+z7xXm8clmq2vqyhmK2NMl59+PGSs69Gv
RBMteik4qZMfViF0P6bvAfRZaERmbo4xCKWUTewKEk+P6PtMqw8L0pNpG+s1sF+8
c3K+T1Fqsdc9zdDZqUgbz6I6au8qdNP8sjBu4o62Y/xnXR0nEya1r8c2ySLOZm+j
XpWBodJn6Z2s68laqn+zi4yv4wYrFUNBrpWiMpb1dirixWv+Z3jllzOfgU54BotQ
2F6gUzR+odA/HhZt7Airh6JAIj/Yslx0Zrb2Dp3G9hc6epVMObyw+y3ILa3ZDoPw
mkRx6lXs9v5ObFdkycgWQkSY2MwFaOV1QD8tSZVYvCd0+l8S8of5lk1iPcncNo3/
A5k9BlUU5xsLQKsJaBKuNCsYSBNPl2DaTfTfQCN0OlJKIGRiUKl5yP+6Kr7NVyo0
/jbCo9/t/ESf2T3ncolh+ca323B/+FsHHcbMDdBxWYKnq5cSkurmXs64gQ9VKJyw
PKQxI00WSGyeCxeQ1/UyLeXni7/JFKDIsxj4AfzBerhyoprVubJcGwVptARI2CX6
Sna6vV99i5TuhbTEqwnYgOVHEZHfeK3Lhp54d/isSc83ZlX0nCRA9U+oOxO3Ee+x
IWF9gcU6SJXjqINkQln6r9Zj/oiPHeUSoRJd17ueDvvOW02u0TFaEQxHTCVqbaaz
VIKsS6dVqEq9fY+0GOgdnlRy0EpHhw1cpRuOoLjMnD61IU3jAof5aSGShHx7ZWPN
3C/iFEvY/cHkWHBXgCmDh/g9Z9HaOxDSnk9Y7LTaGDCSTTeEybLeDr3FOWV8eoPa
Y/4rio7ajBS31jFp7PHBzapooIB649n2hdLzqowKmFU9RhfxuOfcucUjMWPa7uvw
cxTPYa+eC9wt1RJWmhbUpp0Aa89PyyQV9Zyc/t/AQPsZ7I0pk0X80V/1AGinD48b
iOYfWvui9lHDb9kqbFhEQBbAvRaswBAxmflrW6b9iGIFyEB9ShQyOussyz4x1QZQ
KM6wmZnAX8o2dtbKKtVD8fDsJGprBO6ihnxDXcAiZ8IBj+hqk9Pc7tzUbZ4EI4Sh
abVxu0TNJ1d/eZPbZKspvkKsdFHEHdg/RSr3wIuMTOflAw0O0Df4nbzJoMhl69bj
2aNewByiGMujiGXlbS3zjDmh6KvQXWWPw+AzBkip6IE9mUcxGcvlqL4L77iexh1F
GnwbGJbh8Ipo13aWszVk0NsqlkJfnpBG5nTIN5w3tnXLTcvT1fhZidu2+QtxWpdr
0umz2OzuX3oOBUZt/HvWbjyzZDJLlji9XXpcs29Wf2ENrmiBw1uNGc2Mox1NhXyF
qZ8oHHA1a1U2WtUXKQTxkTFdstcnAZTPqSc0mFahrqdgo4ow+WOhUBt40Qfv96fI
w4wGqInfLjUlYPgUHYRvWvY/K+JokLYWwMCQ0BEzgNakVAmVo352Ac4wnur42CU2
/RREYGSfysGx/u8TDS8NZSM+YJ3HYc7z28DpLMWPn4eTs1pyWUcUmVZa+0QIFFFj
Y0woOpQz5kUkzIz0cHRcizOy9dzNBjBs9Dprc+fsSgArSEuds10fxe1UCgY0wpxH
KnjuYuK9WiCFW19pjbZbrSMtxvzSlpFsiYgMZzCPkUDaC/dlMhelWcqx60i46TEp
Rvo61VKFZLmzBfs33J0cnV1LZDG7wv6Y/XiIzLNgC4WrBeHr6ePOtG2QMJj2UGcX
ZEaDs5SvqFWJWAJfU47NCuYM/PnSkJj9c0nBpnMYUpLVS0WV9z+Xk2RMPyCKXGe9
zTWogCiOE/uC4QlCmufTBqCkflHoEr3p7EvUc+tFk9P01OWvX8jupI06HGPtZ3M+
pmWiLqoA9vkJgC0L15xtnOvDSXAgdeVxy1bwM1pqst6fy5h3ZNezQlS1ziKg7bX4
m8/CCQilxiJbbExpP47/YNzpYDlJGo58MQhyb+TMun1Xppe+QfxGd7cACXWYpGh/
/69QPziks2gPcEVwrUlr2p9mJCl64cIl5IZJ0MPKh5uTrvF5mZp5D7Fjl6W8zYYI
vhxJ2mMnohOHFDUtqy6twPBWlx785PNbnfAA0aA4CYz+uLqIbnxx6Bt3qJIRUUZV
rqquwxb786iM0hX2cRtt5D1+oOcSOy6CCJ7bPjNYMlSAK/dPai5aik2cIFSIf8PT
XqbY5UWQv63qUC8wRHXxSPcDbnUN0G2idaglxfKyWkiqVstsAyKQt8bjwtPV471h
TVWocwiVxBx0NljMNZuJdb5Vq3Avy1hlO5HH/g8WAt4vnatFAmQH4ZtT1hLnScvO
+8KOz+G5cyEzDpS0HqpU6fLmffIRWo2BHnDi6HqYbLqnoJVdTHC3lFn1ZGzPpm7s
LabtjKqYMsIn3IRUcVCPI7xUfFwsqq/7GTOHd4W7EAwd0q0r4SWBvd2cyrFSmALl
fRbQqyQdzuNQEmBBjylxDLgbEw3HOzhOsGBA9cffFFesuzMxsKp3kX1yqSjvN4IA
VSVUn3ryXHw5Slpk7MBgR774laOGtYJjp98lq/vQkEXUKq3Pdpq97ch6DP9G8PVu
0i7K+3JOultIlf8EoZ+DUSx3zeqb1s8rHL/aJT8ivyHgT1vcDLO+IB0hKmRVVyRv
JhHWilYf2U2udPPcnhSBqP0dClZtrt4+J6KwaaiYlL6ngpdsLdcDEwaf1i6uSBDA
dBGyHofzfNWsEkt52TbzNSK+mYTUfnooR8MI+SaArEEawo75BohXYiGkqZwCL4li
6n5MqqJq13yvKolo+1ILpk8MxFExnfyNY2H8pWaB0hOMEPMX9Uouv8JQbC1viAZO
y7WnMeHDXxDJ7TVV4VINleCafbNTPODdpblxIlPtZ4uwm3970k1zFgWQl4FcLxtZ
uovK2IOulAxb/X3b8U6qb88D2ltEYGc0F1uxA0nVXTtNnAr1sb5P/BZLJtrHQNOJ
VWAmFxXKGiT8m1D+R8FUE/hI+kzbXZmvqO3oEJefanrkfkNHWouPdxd+IOPbj6JO
noxdWXOyyV+EVjXUQQct9twXPTnnlYLo3pAUHWg0hNC3JApEQApoLcxla3Fd/Qzt
Hkh0phtZ0ow+9U3uu+5U1YGyY37c1FZJiKrd+Y7Tjmv7GZnvWurCZ/LHXM4cDkXd
B3299QTz9Nw2+UtWfRYLkPVaaNH9zpq9Hbeurp0fpvVWo0xxwZtOsMoZ40GIrSqa
h5glRfxFVNhI+TS00UEV2EW0qpuuHkneujyTikfQxDj5YuOzo1l6IAHEiGA2ToJm
ybzQjpeukMk5dj0InUHhkQCT2QmmmowxVbYzyWOE6q+hRMNoGgomJOu3hZhqqHMC
LqnseHmnTtB+kM6aKEbmXEV8fof819MJKw+RVyk2pNZsKyibtd+NO8RR6VpU1GCj
pNA0Hqk/h7wFniDs5ioi55TIWuqAxGt8N7Fi4lghvZdPDsQtmEh/QqviFxIhmrvz
QklQ6AdczYnPljvPg69Si9LuG6Ve391bv2CiSEkWrOKVEWKycdt0yifG2hT6cmPY
bIvoaVdHscfjTaWTfVTBdup372z0xecMCsbhX5oiNiPKrp69GQjqcpwsc2gp444J
QUNvGbjtw+ZaZ7PokpqcYprMTYkZ+Ppw8uDLz4vh6208YOn1Gxi/XRjxAEwU3/H2
paPBtiBA3IXhknvGhfdcyp3I0d/MTpVJ3lFbtwRvKVAOYDRG4Hi7VtPeOcY1zry1
SYRbIWvwBR26rNwRcV6wYlc/uNIvqnO9OPfE2o2LEiS4ghw4SZsgJKForFL0UVAB
sNIXdycP6nlF4waXtbChFn2keaIoObPtp1cPkkWkg3av3q1i+FO84zJb7FjG91ZO
XRtHX+ZJ32m4uS3Sp5xjR86880LxVW5UJi7iC8hl2ocCtZujTlXqKCGtI8L85dlp
cDc8Z2SntUzpVsRUrvtbbmkLNFKSybjHGtz4gL8pf9uFDMMk8dFDA0p9XCESaW3q
MRjJvhl9soZdv18JCdkJ30q7/IYoHMtl8YPi9JaVq/HHNEHU8f3WULKq1QnMld+l
Hcx0B42ExvtrzBQKDv34tRJfi51jXRdnqtLhU7wpuoqjM6em8uD5UUNBXO3/CIHL
zaprKjWH1AnVX7yXZOQdPBMqarYqhT0srn+ajQIia9ZCGaUYxf4Oq70a1pM9H0dn
E1pWp8ybqoxUocDCSMSU3v3f0S1JA4mXFmyMazLSIEK+GSN7cXs4vm/NZ2JCLEoX
ZYCrRXYcaztDozI14UBABfOfRnFsYm2V26f2mjyAgsicLLghurWPv401/KVwZVeO
bHeAaPkliZtcA7Yp+n7s5mxqGIRhoimK3tpv46l1+cfcS4A5qysorfiY9NMpqIP2
uqeP/qS8MUInN2983lVJs5dTUiSFFGIqs0xH4S8HdbwH56tNqSJGiHw4NN/46rem
7hEmf+RobgmdHHZ7r4kyYrZlad6T4eExeumkvabRUwSvtGwAuizVRIOT97x7gGGH
XE0WFZAc0sn+SQkb8/vKniZBSEMYsqqvVzWESQErpEdrlOMWY85T4SLMnweGd9V2
nslDBSP01UUlpJsSMLXfr8aayF7Mnr6CzS6534cP40VuklOktfcBENmA1umBG0JL
YGrDv7i/i5PGnJpkrbGP1paj9IfVP4eBeELd0FuCQvo866uLQ0mOwAfVfg1JZN0N
gGPNRfZIXjlK3b3ywW+E18W49v63/naisIicG32j8et2hvkp+L8Xie/zgmL9CMH6
XWs2l/kuIpFad4m2Z9VhG0WC7IVOjdxCiRnzPN7eHDQBD3pTaCtuswQayEDrCOMj
w5xadUovJXWFmwtsUwOQaMzQxvuEcIQrnRUm/lUh3fo8bEH6kRHHbC6AboSRnV2Y
20FPcSma6WYZvCaJDBemg7en96WvK+shhjb2K1bJufIvrFweilCdmHtnA6f/E+yw
xgi7xcFiOqzYyFtGJ8jTFxZxbpa9lia/o6QxKrjcZ3fTdAjDCdRpJNCAxtENYE4t
RyfEjud05DiaOhF8jDLHl9wXVDAjdwl0h9dWGp9Ly51PZ6ov+xKzbDq9U/j5VlhY
tCQuXX5376hjVhW3bWBx/eTKtANAfqIRhHIw++Cg0gp1Y6wAxeYA27rDVjFrJFGy
13Zh8d21JnqzHHQX13tNhjULpF0LgaJwbeLXLymH/s5v8bxkl80JvnIpgbjarY4w
xnahDHvYNJ/yY63iZPkXHFg4BY8isGrTl8K/NSyZt7oMHy9IXJWrwCYazwyENqsB
fSqwNh7/pjCJRHZlswyh+5h99mfJA/E+WU34DX46cRhUTDLiOJ8tSAJgJePaxSec
IiSIHkzJx+0hem+JTsn107Btst360Od6LnA0uOZ9/EUXeA+enxqd6ugAw5AExCAd
pLphAxeTv6xn9B9ZRJDDqA6rSV6YyTPWfe55aKUcYKX9JUDviJd83IBqhXFPEMYB
buCOrU1/EXQcqTglrHQMosGNF0a1h8CVD9/AS7bt2uItHtL/G8/rfYXiRr3mwaDA
QiF8pg/vMlPZONbOedLfKAV3j1CbPaYLDvlAtYIHkJzO9twEMPWtQ8+PR3dH5QT6
AYhWc9I/+70bJ0/Je6gnqMK3nH26t2shXydyucJchhEMYlvL8zO9z6sfdAZ8QYgw
xLM5dyz4/eh2n701Ce6g6cBsCX4043d7X25tjCk5NYj+aKP3P0DBtJxsDvm0fWs7
mXsapMBQOfVugOWdM+EDlzgYYsehkySGQC+PhzTCP3A+o0L6/CKfaeo7kkBI7pZ0
Ygc2nKfRgpHCd1q7gICPhvGtRGutyy9lDmoUt+GNFbytHSpVI9oGbC8WsXJFJ12h
89+518WhYTmbtdki9Bb0Ob6Vns8fmDlwhhXzD3HKf5mFhm9tOX3zsN1B2SZ0tuf9
yGqq8qb8QBE7DvlydoIBEbnDMoBAHfsmtOmS6CnYF6JdahS9M2D8ehm+q3kLwDxh
62hkq7eZvSADo0+d78CLJXslXfdzRfziBkGhDTiasBgtJul9KH7pYv4Gbkxhkzs0
SDR1zQBZVamUW8//08USTrfrvDEAHoG6T2VL429uvqd2sBdby26eihYzhGLn9ElY
y9gwyKfxWGHNc88nIgJCwlv3+G7cdmQw5jH68pr1XrqnzK9RXuEKnb1402J/2J4X
gkcBqSEn+c30QSxA26mHqouli5dghO2ANsBLLGI7UzlC8PGy/paL+h09ttBv33do
us6KOixebmx4AzpRZxTYSejg71qa6sm+MQK7CQU0YIqyj29VgdwJqJOfPiAnvQGz
m9FVFyFKodgaSxLPDASAcF9T7jkq8orIrGi/D+pEroCqYVfSAEVqr3gDrhjWTaMs
F5G87gg+dcs/Irzv2J1OQ+keL71HZ23Kdw7zjuZ9w50w+WCsIy4wpAao+HK1PTie
h72ZaK7qcFv7mt5WosCbhP48wyBvcMoZ3QP6toDJrxRFMfp5lNcY5ZkkVzHjBEdR
ntUFpmvz8CN6f0ts9yeC7LorYW39+2HriR6IFWJl7GCPYDepm/51ji0CmsJLSI/7
b6Y6AzjHhzU3tg0Q/NUM3sa3WbB53awfKiIe3eQlctYgt+LT0FGMwsRYnGPAehU7
sAbsh+o6nT/PlonrL0s1NFBfs4IBbhN8AYZP94twLBoiSA/1G0BzCYL2imzar74f
RGI5Lz6/iyZgcczPV2F/fi0KzkIa6ynaJYEsRjBfp1nDbtOONgQKHr8/c9/AYYj3
kFw6dkEbeZNujh0JI3urBQ+s8ILxqa7ia0e7RMqpRe9qkQ0mlY5gpQW4LS9sB+3+
VIpfRw7Mt6fEYZAdurQtS+8BTvyRGpVExORR2pZZdqNy2oOR1XWdycIdvxDdveF4
fW0YYImHekWbBh0P3m8yfUr51bgqb7/sg5M527LkcV4gWzSPYq0YItxgdiaSMo55
RkI+M/u2ZQ427rF5p6wzKmLCfkT0rCKZP+dkpv1hAvyIqL04J6n3vVMEvn+eIHLF
9hz0YIbHz87yeZoVZ/NuMCO4XfeXm/1zkj/SaquCEZsHTPCpk/hrFewj53JEe4yY
3SLPsSURg3UJ6VJAeORei5AAAG4tKUp58HQ/vKvDAo3jDpWvO/EUuhQTq/3/lH4C
T7EG/BlraHY4JOgJ8R/ka2n9U2gWVND8ZoSzCCAUQuT2DDx6l9wpP2sglcXS6zoV
kSiepUQRT2y5CcGM6Y8Ucng1tv2URrPWGsmHP4au8PTcS9GPILApdW7Bvj8hcnF1
rra9EGy1MGmvV3hBbzQjf+C1e/rWbrNNCyMluWsH0mNOUc6A3O4/XosEPGht8PS9
RQGqF/cJ3m6Vo/VY7DjPh2WqEFm7iz72e2mKfkymzjMDgTSf+bA7DUxYlYEKtcOl
eIOKUt+tBhuwOWQgcp9Kp/rXSE2yL8QwT1z42oke5OjZIFMFZ8wu3pzOQ+JOEoeo
hxliAlqScSxe9sqs5CjZ3MNdQMP6Kupt3RTotmsc4Lmb2eBelN9Ch1EFSzG+o2lU
VSo5VaUkLhhe0I0pgaUCo5aX9OFbsdH0RpDI5QTHAz9R1MhF27zh2bnbRCQgQiM/
qw+V6b76O5/AamCzCtJMOgIQlEwtobkV/KdvvLLthQEbDK0IzTMAoh+CPsbrxfM5
5FPWFe66atLsjbUKY6eo1+lw3XVp9c+nXWpoZg2Cst4awIbl//ppjbZeV3GtPHTe
7GxATRUgB2XC+5nkcOztRfUZ/7CxHySL0arjr5uVdPO6uDUxNW8Uto/r15Q984Qg
Kg2rNqIHsN9wcxgKPkpjiZPrrcDAcRjx8E5JKvJ8MawZ+FThSbSv0/totRmRZl+F
R2EyUyTInh+AnxEkB03js6eDnPl5hyEwdWFk0+0G7tS29bn6YqNmFjeaKJTlTixn
KV3Wdk8r2jGZcHz6n6dgciJ5nxPYxDCdbFJtZahqkjfE3kxSZf+3tGf+BeethsJo
iKW9ibA6MUh3yeXZzdzDaeuaz7guoMjqtHxNrKtCFK1Vntt38Dvi5VrzmCpzE4ep
UeOiBpxtnQvE8kTvEXL4nT1/pdn7hnODbDH/eX+5qFvjwpXe9LhhqJvUPdTLd/4u
f8mi50ngoWbmhW2jGWx3KeLO574wEjYxdIF++BgBUHE2VLtYfrznuZTcwvG/pVu1
4Lyaha28zrYVSx/DvK4aPi1fWw4TctWs8WSY3l1WvE5Y7+i6h3RQDH/OWPjq3Y5j
r+xpIjPhTDkXOMKSvGwy5wZ5jghJXWdKsWfZT84IuRkVnlxgxPQqSkP5OjXdcVdx
/5bB+5v4n96pEr/Cq5eRRRiKoUtzbsY+GobWn3hklVS/NeW5dGCCcaWfjQQlqiXL
qLglGwzZJtygMv4tUpm8WmXwXAtIRDFCk7GhpIy0BvPoZDe97R/KwxFAIh5ZB7YG
8lxkt9tmrMBKCAc1mN8yCh0wBGyTpeHlYpCf83/c3sxh0QVNalx5YJaVqr/k5V62
GEW2tZ57D+taJyhJXxkaYPnzsLIsqfKbx3FW8U60gPOJn5jhb68ZntTAGAAI+raN
OuxxmRMIicNhaxKBX6Pj6fct+K/22YybMGAmTVZ9Mb5LzL+raoXT3d4mYVSAT4PY
0gg1hZZcD9lBzLFnb6tfQmHo7XSjfeG28lre133A8oeV2uflsTL9Imrxy9oV/o86
ImLwsdSL6v1tSndiHo/CgO0n1ccZqCEObEJFRioWi3zVgaMc97pty7+57OXmEmwn
UiSjzntUCDJ8LR9YIMKWV9AvLEOHCltrpnByGPVFMKvtdIBNyPpLUbM7b044PytW
X1aNbpDnjKZQjzcbnQJCY/yHSjPNYL8FCsODQDs6hm59QftZ8wjmzQE/Xr+rE4j1
Ut3z2ugUH8mC3s+c9ZfA939DN3OZhCFQQiTCCORJ04m8PiMGiKTHIPLfWS1Irygc
tHMwoMGMuHd5K6iPoJh2RVKFijvktWtQDpCQPuYFEEIHqXvMI6cIG/Q5+UOMEsLO
5QCiyKdmIq5/++/82szjxSTQXfgh11qEvdAhkI3HirNr+23DlMa/oBCgjo5Tk7le
z4s+bKBKpfqDmrQhIbqdTHFUwLG4uDd6HoCvt2hfvDm/dZDRpY4a+ebKuxxpfvs8
agEwfCDkJKJ239s1zy7mUib6ovwRyilEuiXmY1c3dI1iJpL3FPOKStPc6cfkJsPx
QSvzXolcgpeKKnYDxcg4dieF8eLu9efv78h2i303aSej4FicIPtiseMxiBTndWoP
8rJgHxf0Dv0QYJCmcJ8BgRXBfsK7dQwyxK107KIRxGv2M469j7lCe6nIXZzBK728
xDjqk23amJNPyBd5b7Rfbi/XuTHvLPl7HSiiseqoabbOmG7vQcMEoIKYP7cevoQ/
8bAE1mXKPL/H+7VZBNqrbSYkvEqtGwpmFYtaYjDRxnkKwWmJ+cMgIviEAKVlzq/T
9nhWqIANyo1LMh4ozWxaUIWTcm8ECg4hrzVlTkXImvJHbxRzjUPCb4yqQaue9UOC
IX9eNZbPiR2/lX5YDsBPmxQrMEZpjz7iCNQFO+hfSWDaLeg9dPgB42CXj+UfCs+T
kthxdQE5Ttd2s2aKJqOlQcCHNUat++SQckPKAoGnKK9npAbMhHZN2RSVohkaMxwa
j0cD3VyC1yuCYy24PZbPRMDun2AyP/H01AYH9NBR1ZkubKkJYG3U6quN7fQlzXvy
LD3riolFTYxJiZcATXVGXbBlJLHLO3lo0+tvVhpvIAeAH9F3rbNJmfsQ4Q7wdmy8
ItqKEGtXxufBT/pLJINESqUw4kUaAIfxmyaLf2nYf/IFZLlalpaiB4BtkTKWEtwW
XkQmjgb8g3wxi2V4jgQ6rYOnGglphnZjiulobvtdZJE3YFYkLoOxnJtCcfSveucE
fAwxi6ktp02Rw/3WWYgIVWhbJtlrkDbC2oUKgE3M6zTuoJyzUglMlk2+FfAfK6Yg
+arTBChIrbXzghVZmLNC5qjg/cpggp5dsk0lCEls9j/damHYuo7bzE4/TcLKVxjF
Mdp199pqnUs29m0wxLopeSuM6WIavmjlDC3UxcZmf9FkYE+oQQ1YG7fpWeM7HtdR
oNjypPKi+UrdpXfevmsBrkw8iyMZmP/SsYbEhzG4/yj3usnzTVJeULKtwP1ySBkP
jJ90HTGh9X5fdDKtCJGHj4+o8CRB6TpYG/yGhHMXpr0X4D/LHmxnovhvR1Yj8jBY
VqRlNjBE8OhRnpTupi3iN+pHpcX1quD1aWTjUSKiPXuPf5K+fgohYeW9DTqat4ht
5oAxuXTXJSP37qhdG1FwXHyGs2ZvL0BguTw0TSlLlAu+pB8ZCtHuWwDPLQnk0DM4
p2m2ekYLaTM4VYeLmR1tEWRDxvX/eW2gLUVLUfq+OqmJXxY+fcq6T3JwiowbKaaZ
nYDUwM4TzqeDV7QLA/hrSFiU7B3sKJIr/ErsWWyjQBRGxTcSzlSmtxFPDElV79n8
oMkzcNVgpCDVCr8viRbM6iD+eJnSDfHEDwN8FoWsyhUb6qE3qBo2nbMp537wy25/
6ISjOgh6gUCy+GNtgvWyn773iqKWdZtvlveeTmocI/1nL17CGxRfLlq93qEpxY8V
5oZbhRNjDjTUedkHZ7HtWw714gR0HcDvGVzYdltebc/BZDDc/c3tJ1MX2Vutgcaj
/4N/Z5lJjKuSzkASwk7oau/HqjuCr9q4Nt937ixugOnpZXf73PsaqAri26uHDzB0
rJJ0jEgi8Eu4/BfyAahWhNWUDj3R3zyrL/WvI7DlJP40mQ0QinSh8qat3HZvPDKU
HXlQDYWMB0YqE9CGCei1sljwmQ6K2GxwgUpCVcxEgR7XxDzrrnNVNLYPZnlX+5vT
3BTC+3/wBUqVZhvwyfCDGKedSbN2nJQI3TBzuEJZzSdP9Cz32rSdcOR2j/UqMwdo
PFe06eRNjjcR89cuiv0pk1PgRlHDJror6nHtihApK2p0gmQrmZXy6TJi0hsOTfcV
RGrEnayYZ012zMp+I0ONMVcjt3pJjWin4+himsZrWJSOilpb9/i9Dq4+BHMX/IfX
7hXZf+R3yq66Ec2zgJGEWRDYL3OhFbADUouXiWS7tOkcZU2fF2P/mGa06WEGQVLS
stIc9dvAMq+3BmFObjpz9hmjMivmgleejQFDCKto2m10LEupB49tXpacP5eB2hja
xYpSm4mb+gB2g6tB3/ufjt2U+OLvr+PdB1dkHk0mcPfYkDWSsaUANvN5AE6hrFYo
Qhmx5sNvRd3pseOXqaulXSPgSZYq41xQaedcZCflDcWZnKAjjSuhou9LnoqS6MmB
8m3VVZnZcXok6CncoQuaYvZoxv27wLplzB6m1iYL4gfPzqhNvJVtFkKq6QVSYwIu
sLTNbx9cONOgq+JaVJ0mUqLCoYTyM2wieypg3bmsAANey5nafc4nM8vGTMnJq7bM
FVO8zueY/+Kh9RzRM0cglBjW7ypj/PMbFIeKu0vA3eKP2zobVE5ipFD5tfZ+A2wp
5uoNItpQdyKNyzAwDT+Tty4l5dabE2QdBnUZTt6VfKN7drxJ9LKbt6wQ9RSEpM6O
RV5vJIrw0IjBhTxoolO0EgXg8fC6kYXBi49t3MviRBpkQyvLcSQpPCuBw4P+mkTW
jT3oQL6qYUcBR+rwhJ1riMnL0hNNbEN6sMRQAteybw/Pbl8s0hOa8oBmsdnOfRZ1
jObefGqFMeSNOvyZiqs0sJikx29Z/ASOmhFnGWhOIwZ/0KfqitGZzmtMS4qoeWLS
nw8rG3agTGGkgNKSj4rzVuPQoQKF7ntrMUbjwwq2gXXhNxZOf2WMD9hQO+hT/PxA
kE2nlpRaYsY95We2ovEuMFMHGgwgw0DagqrZW1DrRxZXoi5DSqxbyf2N2pRHwadB
EzgLrXVbcTMF+jySz5VykiboTqlPwSRqcheGBRoCMVlDx6LUGoZEKGDX+iN3fdcU
siAywRr/7fD00aOzegItIbUnrK5Rr3k+W+0tidFg7Fa2dOky+PArH6/lw5vdttqA
F4m3NxXlSEsF2HNe8ul4hAXs7+FCK9JidoKbF19Uwug/8rngmfj5MGJaHW8e/Xe/
ADEBKmy4eEDzDz9gAs/DLxYVJcu7m04zZIdUQgA5SaJ5ztWZVa93ZSVYPoLwBI/z
apQLdWAC4u5KEX+LahtGeGvnvkVtq/PqI/sclITAkV/p/1pP3umWK9dweAutM/+9
FHpxvMu+EJH0Zr8qSbC5Rb0Xvra22xl/sbUynaneEjiv0PZmp2ArZyvmQq2w/0Ka
yfPsUz1s7i+u4Kin2ML3PhTgoqI4ZZfEt5wdsJiCh9M2WnFuKHJNd68YHRiiRhTF
daYY36gF2MHpTQhp0ywjFGsns5ocyJCUOB55bVMOgbb1bAULAt2eSmejhPgO0THs
ScfaCgEwy54//OYnL3xYD7C7E4k8f67tyNEhWSsMMhQKHzdSAkilgudP8nxNI/EV
GPgCht3Whq8jlsCnO7LNDWa/45G7BjdDDk+CBncTlqcDs4aeeWtNRq3NDI3rCwqQ
xVPYP7RWZ8RK3u92+djxViEJTW7hxtPFVQULIcdeJa/QbwZagyIhgBf8o/v1dHw5
FFa+Di9BzshkIR4DyVjnQDoBTuzclOWqsYe5Ox8Ar2/PeOB0DHfBYM9NcZt1bBW8
llmwtIOUXP9c23rLAsma/4wXPBXI4I6+JPBsH7ktEcrM8OfnSUYJaOZTIFNQxIfY
oJRzHPM4ixYj6xUbo3HQa4Na2BKnSCNyY/t2GqHFvH9vmnQy19QT416JsQh/cDri
gn59eEJEEtFFKxN/Jv4QZwnxKdQaHWNidzL+CmqZmY0PBI87rii8T64gFHVpzseV
58kXqR7PC92ugqWmp8gHxc7+jCe0UxKegcC8TSCDq7KfIbigq7HogRHsZOGg61zE
d6M9Cg/Cy9vqhf4ek8JQOEcHbdnG+aisyrYAGXF+Behfs7q8VEFjtwejsaEqZKkg
Ogel5adtanbqh6IkEXgyhZ+RXH23O5UqalVqO5uQzUOYTO/cCosy34M8uTup665d
ncvQIvlQszMvDMPKPve9iihWUBHuytwjy9A/z9Cs96kNg7MJNxKby97LLlYhzorF
tYjItJ4bIUyqp+ntBPUfaNS6roLxfjKo5ybc+uOcnnEMiIB89G9bYGbRKTICrcVd
dxOpuDhFfFe8Y6oNsY0/QztMHSE2ECYhrw/Ei9HOdcxNqCnEIq9w08MjS0cXE6gl
P6ppESRDXDwsq9Jk4Z9JLmEVkErlEC9ALFawFOsDe8RtVoC1D9xxSnoq8QY3d/Ch
0FeHsWNfbnpRJMHjzQfmD2JMygMDxqNttElDYXuiaqQmWqQ7Y0w5QjV4tGw2wm9B
hqj+Dp3oaPFJvC3EVS5gI70TW2aQytpR1uoMsezVuwNzAMlbZThVihiOh9UN81B+
MHomU2w/mEcKrSMw7OOUAdMvVHWG9jLILSIWVxtPRcgd2e9VZaocpZUSJ57BFTzP
3e6MxOmjw2VjeeufDxLUp/s3IuC91/uDBg72kuH9RAqjcddaBrTE1yyDbkT4VmP0
ibjUWPH9MmcXAGgaeMLzq9q+TuNL9x6z/4paKV8FIjekxE0C2zg1pFXwfW1/YQjN
jBrqMP4MM/P/ft3Jalm6X75QOXUfP8hgSoFn5yiRxHNJe6KpOfBR2M5TfuS/HrbY
v6mVimY0/lgjvKAVqnYSYIIoduG/phH6oFvyytAcC/HVcD32BiyS3rpQkopg+wal
aMcVGtvn+LeIZcHIEPhIwrxB3/kb3zBphyiNWTxVzSBKBP+uSMthi0FhAUaUnYak
LcawvOSALwzntE5mWP/LwxfKd4abv5pDYDB1k5YZPNwAngV/Ro0r9lHRBU2s57zQ
Ib62GGdP6c2WFZh3cgLZJ6AwfbmwrkJytSvHAzcbAp0QBe1vkBrVhBVzmVCwyEp1
pD3ZFIEPjqlSU2TAnpnCeFsOULhQTZHzAKecsbQYi+gaY0a7pI+ZcXDUayat9Ywv
T9RKTiFwTglD3ClJJInmm5YUDITN64tYbkeJeq9HlVOrPy9+MsQDodjPdZNCWOWG
Hj7dX4GYo6bt24rj0h87wh/1Kf5Dq8/RIC2GIVuGJBHFgP+c5VRP0oEtmqSFIlVP
eg/IxWg8z6VAKCeAzMz/nzso6UJqt3hIifoov6hP0oTlsNLjI+UUofYjI/M0iQPs
6qcloYcS4jIpNficphHQ3xb/jZE8oK4ea92ClvMuBztng4HKGXbGmw3kOSpABF8s
GDzrVhFXzGpqew4+g8pGU1B4bVEeBYZRRmxux294MLPkR6IBaKd82gvtqvuuVwON
14jPWvzvNJpH96R5fxyNLnYyOyN1Y1LZ24R5jDM+75OfDa0/YV/KAlUITwT9RaBr
zWarj4I8/FoOo7uORDE2jST68Mv0qJ/lmhr87gVS82oHL6qvrmsG9zOavOTuwOsQ
lVtpx7aTfhgvApwD4Kns9F0a7ccxBB3eHtWoId8t+iGwVW7b6vXodzS65edDFKsu
dgJ4JdYmckhsu6PmQmKBZZY2m0pad3CNkMjNtIZDfPhNlCA5BBHi6XvB/t5eWoE0
gcta23x8P5MxhcJfrfEBL98iKedfr4iBcPo2VbV7928q+FyQS5L39ljNiGWhcRdK
mkjMyo0Fjpew1YEMI8HbJDhK0vAbiIKfbn/23dEtmUnVzxLVBpTpI+c9atiqQlgy
Wx6RcWAQoHPlAftLZ99ViuUBSYVS7CeWTquEokI8/Gj3nHmzh894GbTKyrFtImvR
4KTedPPoUh7kgBd1nyiYZ8yGfOj/0N48Zw1WzIxzipWkM7ZgTglh4bUlqAMZb2Km
r2EYm9ZIlZ1f8K8YDENkATOwWd1QrrqPd2EzJkuyOT9BYRVJQNCKbbh4uMa/poZV
MM7agIIgRsJoC3cEtV61+sfV/DEk5G4MzGgpage0VtNjCGC3pZChdtDiiAf6UoqF
xNl3B/GIz1ZIgHXB8Enix4fhcvKxQ636CBUixtU2v/n52PvDrzwgGOXGzTZRnpf2
A6G2lOFzeb4cPDD7GX9Dig2SOiJLdh1qpw6eTHdfSkJ5kddOZq+i0qcxi+SCIZo4
ybt3+3KxPsFqHg1VM6iCPjkrtdpA6qI55d7YK9j6P1LtwfvVCjXvXYl7JL+qrRAC
OOHpT+YEAHl+6yinXF41F+RvCL9YzuZng9WnKKxKzMRu01OS8OzdAXD3bfTVA/ZD
DmmxiOX9FtyBE5719CSYT3Lakc7vVOxYexL0xBstAY43tcIbX410MYVK7T1QkX2b
ya0dIwdaE9y0+RJaFrxOhbkL4uJsghotwrqiWXtIsNiVFisdMjjcIcaNjJJwIJxB
IU7kUzYKBFzWuiArytEcCBYZRLlMkbCJ8EMNGivZnZi9pAAcR+2D4WvCUhESwJYj
NCYZqvxs3Pg9nUAWWyf9uFLVe/7efcQKuRGYlbaCXz7/mzyZTcY5XPeIdCa3HEh2
EnTz4u3f+Qm694HifQkgx8OaTROxcVfAqWeX90iDmBphpP3WuSTGCHJVuRbpRFTX
dVi42W+ySYU+meGHltNFLoXRQGMpjm0XqaSCfW20QucBSfWEl7nWzhEeHk5UY/FH
UlY1RZo3aUKFAxF35+EFpDlbw9EzQkM5+rMPaEl0cFe+zR8ubawXcT3tP61YPvIL
Un6nWo+0YmW0tTd4/WW/gKsvgPUwcxutNH1mIoa/He3NtaFFMoNaiRaoHI+dtHWT
zNPVBunsHxRicDCu0Vd0ue4jwchD1pY6O6gzbfPcYeWfQiU7XBHP5EMyWJ7LMLYp
hIc+5y6rdpbqzM8DpnuI2BUsijQ2kUToXDI8R+9k0nYLLdVyHbdZweJU+o7ZybGs
OCqs2HRLd2d+DkHBEaZwZw85qZXwGJUMFzNrcZqlA+C2Zon+AYNrttBgCDdeztmw
zipZfEbpxgkxlq3JGfp/ClJFTM56wuzFBokfch94U0YLgfDvUcZNOfRgckZheRN1
AKSa9uOy/V1VOfTmPMk4y1OAloRqOt/j1oU0wHBHar83B/lKKvrnsxoGV0a+oUbR
f62ED5f0OjwiOlMELwSV8/NwUOdn+FBZmGxbENmQaQviyOmhry54M9GpYAafoSZR
IAeOatgNm04UWijLrmgNU8u6HYUP/KptndN72tdt+ACVXdLiN+BiWFRvEc2f9Lpk
64M5i6FGqqTyO3mowpadHhzWSfJmTzqt2UmT8mZ/cH0nUJtACJ315kCDyFXApV9L
mOSnvnyns7CtQkCQdEZF1vCzw2ZX/bkQvzOoAurmBnLYMXs3YTjbmPbFhgpU8USp
vPrpj/BHMR0RxqTIU470y160qXMrKyTNA/trMY/fIxOFidc6kS3wWan0mM1U1kOT
NrJ+hvontvaA5SaUUE+MASaOuchthtc5T5bVgMACxLxP0R+vogdQZENh4yMvIWA/
FzJ70PwQ4kqXYM119r+XpMoHI/CpAEUqh4LDvrGdVdHWvGYrjwMNBwFhuwm/Ma/P
Ex9u0t76hXhYndV1cPaVPF8oEA91jzTx0NDWsdn70KBCpZyXAnpFWlXgT86WsgO3
zHPD54G5SRYgn/idOlkzFUqXiv7B0zYJf/Ok1ifnKf5DprjGWJTeQs/dlfJb22Gu
+cYmWAHxsEai2erR0aBfzGe/W5OTZpdGx9eCKKGpGEv428BQJVRecZYWwGRuKnZ2
vUfY4XZmtcUwfxJ/vhOoHmkAS42IZu9136M8zk7HoZ9C2zNWe8iQ22kH1N3pqRTX
dHt098ggT1CsC/g0AhXI7kxGF/46PfFOCyt24NJsOg5E9GIQ+250+bveW+IiB14r
F4J3c3Bd0vwUDmakWTHeyVi7//E/DvW0Pq9soBVXQOAQT2DT6m7WSwObyALYKiAB
pV+jsa2fyP5Jje52HIo9aI13PXHtAfbNkRlALTHkKfKVuf29q0tt+EUmyfmRm10A
BEaCPFi/21gd96JEPvmq+wAk68hrUVXLW4IXduOkIs3wFfdBqK1kpVSM4AaB/2B5
rhooTmBPErecv3MCKbexsJP96WWEEPh2VpFUHpvafkYZEDGKfaX3W8zURREHeHKZ
G61Qqa/54FAo5wbdg9EH1bMfhjCJG7OwjE3VIc4GgMP1GDc6p1EoqCS9QBywY6w/
I53MAVO9i1DC/WNzgloPf8+UP7z08ev48PA+PeDBHXar4+hKUb2zxqSCu1aspset
Gbp/VLSccYbv7kyXdWynTg==
`pragma protect end_protected
