// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:39:03 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
fQNt7WTr1F4w+aQYBz2vYdWfwrYgUrHnGFwJxaXpAI/Lwoi8c+kyDENN0t+okKlx
qq4h3RLOb+RFHGGokKwkrQcp/eGGorBwdXemMGnjWVZAcFkKe1ZBx7fz3gPkpSYB
x4Rjr6xjvyjz75Sax5JywLCKK29absDcMvXR1b3Yu70=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 37488)
RQraS4XcGPuTv9IACpAcVPWhHzbzVN1UTOMZfzeR/4bLUlmhLHdEj7f7kzmZsNYf
3ErXbyPPAKHMoJJRgbAJwdRUdITtqpb3RXU77Q7vxLWcMdDVxzZXwwyibASclILl
WBe7VYl0FPQduLC5fKHRIhc4JWtVWfMBc/HOisonC1Siv5pxztQ7zBG7UJE9+zC/
ixz6DIGi62zv7YXkiiKwktwjc8GGzmPOPrJV45PWUjURgAecPR51W4XY/EgA4Obn
DULy4tOPIBxwGvrUql6KJsIdEqLbhniq8yqjShH/zWeo3SMGeA62oPnEW9WK753l
WBhRNqUWNzqzCeZ9GztydybBWSY3TEJZXcM8UIDHzy9Na5b4TGJArTBDCmQFQhu8
xPBRp62Dfd2i+3y/JZjDFMws/FyFfvG/+Dw2iUhUmO0ejgiEvYxrMXIolB6IVvrg
gpD32u9ykTW9/2LtFzIOe7zl6BtTdjfCEYfSoxnecgdjS1tj19fayyAL0xi5FxYW
3nGkSgAD2jrLFbUTfrMQUVJuFU+cLXOhcw4p6ifgI1jpfZjvq6fyFQ4W5eSq1Udl
a9XxLdAkCiHFslKwabzHnWPdF1l5l5WPtj7swZmEgM9Sykvh3ttk2oYyUDYqp+2k
YxHZoJznmBkQDzlDPSIU42GuCdCNf8CiENCLpGnEsBGnrLkZAMYNTyWq+6A1zXnL
IWQIdIXbcJYqrm/8f2CuSFELe5hsz7S/1V0TeMb3Z2W2cTndRL9ye9C2wvsPuTFB
MJnr4ggLwnR06CW9aYgjSizJSYL+xgyGe6UkQvqpNKj16W0NAdwLcWmMsiy8EkOq
QZtXdXJPGmrYVrxbKoFoNZpRazFhgn6CVzVrgTI27+H5tQmaZmNuVv2WtEzw5ouH
klaY8lrueqrYJl/dRMdYbLQyimBunwt8dCIFUPEeg7BNSz371D7GAlMK+29KGa6O
XqwXFbee6El+8h6LSsEfQ2i+qnuB7D8W/9MVtgKFZpHCEA80y3vuccsq6T5SH9MQ
bD6TRBKdXo0aBW0s2/rimgcrZIj7HXWU1wSok/cFXLx20M6mLgDEY9Fo8xTf60Ub
oXFkrilc9J/P0sNx1ph3aFc9VpZEvGokTzwZbV8AJYttNVA/xlVet4/tiBScT9/Z
aocgBrzhyR2Zsjwb0DM7Xxs/guEKisdUI68rWnawCK4hhiYje0wgxQl9jdZroeT9
oM/3Y8s/lZrAR34jjMJDyT0mj3nPjdRbkpcoIsLaFiJHzfwBaA5pX0NFNaAcOXIN
qpfneN+0OBjG/z8YddPIaGbx4TRb/TX7Ss1JgLiMO8CoUSbaR8ZLc8vgtl5Bk+sU
lyOPm+k3KNB8UwIhc32Ti0ItEULFIJuZhCEAPJp3/6DIrMu3FAgPyWi8lhF3PSGr
lG3GrnI3rzutd4enogLaZCwZ0BiRolfUYymA0KNDLWaLzx/5hRu70J1i+Q47gvuj
4XKirMbNn3QGWJEOfjkE3NRtzQoWusG1lOarqDuOo/WSA3TByhhhbuUSjDLuZ1UO
oLqMWM7Cj9sVKQUQYofeYMQYU1itBpAUMZe/xZeJJ+0FKJ78+o8fz8wJnl0MW+Di
/hMJUdEcjt5Ahn47BS9irZP3EDZo52bNDGmTjzauUlbb3ITbekpLFYNZ/nQp7E0V
QgrGnJDeAqFkt/3VlD/XtQdhvl1M73zFc4yeqUdyM9MJas0kyZquWk9A9S/fgi1x
wj+UR8+QwFCNtiWWlQQo3SQFN/1voCvwOkekk6hJy5BwEWqi0F4eGeD8OIWkd0p5
rOGnmSK7cvQck/iGutIwyovazPKvyATpo+5JLmQIk9uV5ohZ3HuTEOjW6iDX8qk/
ASMcAUJJ4kcgxQW+sbOURhFj8u2ElyLSKoFVDr0RH5oXqZtlvpYzAX6t7EEtunvU
KP7ureSKauJTsCqq2sUK1ddXNlnk8KKgCQ1tbJaQhbWL4Hs+4Mf4B6XVjs1pZ+B1
kmUaNCcVcVkRdQICDSayMB5q2EJoEZ2YcPWAsTuKHvgeOtOVZ40bEDPhgOG2Ot6S
SdJHjCEDCCKj3x8qAJoTt8YiL7cHYkaPNDbwTaYNeDZyewbt1XGZ5+/H0BZsMcbi
R9DE9v3/2uS0tXESsaZBaM31ANxMiDXTdEcUp9f174OB4k5abXNpXHWEOgvv3Tmw
XD4SPuKYx4/5BqApD6OWdltmNtEplOgeKQwuEPkKDp2IIP0Y1I7S4fOFWgOb9BI8
/NNG07kz8VK+gX9nuYtg1rjVTVfX9WDmTK3B+rc7RR7YTpBHOlP7hszvcL18dUBH
xlPZBbQcGyoKAhCBQx+vxgNYjGcQKM7glu+ktjMT3VY3FkpFtYUVYRDichMdvdCI
TDaBhhZAb9J8iQB3yyFNUkAY4yJ/exAImOvAytWTpis6dIe2MG7cdr10xh0r8XCA
iCidgs6yFQyth4fpZwB1PoPt90JwVUtGO4Scj7LiRCfUGAzYv9++JfJjIji6DOKT
ZayZ5GF5BlCtp+l3NA5sfarLICMRDJRm4grRkmKXCP1KcPc2+Ijpqe/HsXOgaeem
5JwBr8YD37KpoYnvl+ZUK+mDN2/ecPeyYhl95tQ8QX++chit3GOMUWBTytkcmA9Z
qvNF79Rnec8iapoQQklr4ptRypVie1T48uaDgpYpjAf+Au8u9NamFuyg+cxS+iKR
Gmkm2JVTaVjDIuO4vgx19XzHdAOYY7HhSFx7DCiJiw878nlNGkagaHbMBVyzybBo
J1gQDgYtFT3ng1pg+9u6AjfJi3BjdzY1W2DMmBYYlwVPU4nFN1FY427dF/+HiQI8
H7w345bS6MyAQ5O3lw9g3LYQ8q5qnopdoR4Oi2eAAyzP5UfuPkJNpXM7+XL36pQX
nrhN14YjmGev7sni5Dzuu4DpusWaPU8BunJ6AVVruVCv7/tLJa5yzvP7Zv2F6kAN
Y7MuEmU2c1JeSaS7xVaJ7NIx0UVDzyEMn0qKzh2/fqeno/eBMav6HOd0jfXCw6HD
SisZrnjpNC9TF/kBe9NX3x2VOiUqEZgLkKf5SqAtiTc7GVypmBF8BP3TTlzx4IGR
p0kUWhv5oW4lskrPXVYwmw4lQiGTAL/9mWnoh8z6QANgRAq30kKwElYYBOZYyPKY
Mz3rgo4oF32USSvwHk8SeAv4Ow5v61vDDUTqftEwgwjdlVd9UQ8Enrtadd3jeeaO
srNaIhgVormd2AbRmlexjvSaxMAgDdes1aR99KgvTe97b77gy0qyTYO7weMDIydK
cJRoEsXU7sVA3swL1w0DeLlPEbNJTFOVmpZG0WmJS+wTjAaVnW+L7CQ+jRrm4pTA
leJMU8WcEAYy1ZL7wOraoaA+st2s8+xl2I8ose2miehNUnbG/wA/50ugDdPWx0Ak
C9z837wCxW2v486MnioGyGxDEDWJk9pmKcC4/KbOwkNFoS3U+sbHpMTuzYgkvvi4
Esgh6R7GbJfFD6wSuTaBFY7Fzn1Oca0T1o6eJrJLyUqxN97lSgvW/wtP7knlmgYT
Kkc7pdrjcFvremKcqduPMqYLGSy5jTCqRefcDNuygstfJvOLqCnKy2nimpQkY6Od
C7MopCopuv3jnqZqs+CfBuDBrV2Fh0sGEpCuKRwnKoZiFLA6SAP7AcsAZDyQROTM
3sKrgXLpkdqONavRGvp84EZckJ+xRf6o6t6ynqLhZgjwQh8Lglo4M9FFvHK2UaYW
jS2v+6QaH3yX2TpAtLazhJQVSIPXqCGSe1tfWLCyyF3esmuElA8wOubhxQsrQD0y
iruJhwJ0L48/Kv/f0nv8f8RhmCgs6WnLheDQG5MyQaW2GWLarqAQpOZXIeN/FNlD
IysgKRNKotjtCqDCApvDvC0GRKqau6gtASnCZTfyqp+84RN0Vdz857CfvHFV9WgY
yBj0qGPjnjdsU/UYYrNs3cINDA/atptQyTz9YAyFENhQgMb2Hd9hrmag6yuhXUmE
iPaebNI60ZBViJi8QwVSk9cn9RFdiwgDAAwcsEMxssTJaIxuQNW9UVlEuBGOjUNC
sOZGNn1QzgLEdLn0baiK0QjkPYlZcra3kkmZZiuUc0Qq/UflK9lGUgXp0cpE9ZvT
e/HscLfpCSD+oZO4h0aCHKNTK9SzwhVh2iavqns40cteb7BOt1djCD7mQ6HNd2HU
vBvT7hrlVNxUYHJApWqgEhK2YIJTWcWTvjvQISb3j6x1EXgeFWeVMLNLJvjqyWPO
ZLCZFXzpxRfbaNmbO7luKGoJMXXPT07AboWQMNh/Os7B0o39CpCvw3eZ7wWpZFgf
i5QhSyqrmguDeGFFdx+IeqGBCPl3urWtGCGhvuGToJLmsU0EJaiiIR3lil6bd8va
4HZP4hqcEev+HibcG//ZmIE+0opW0tMEmHSaJCA711AOd0AJ2nM1Gjy649XXgs72
AaSM2/jFW+5eEjGYNxdaTXBoKXDZiH9DJKkS2ueNd0oyYn8FjtAKM6rxQI3IRe/k
q9ZoQH/Y/uQQiCRblNDiLX7k5Uqyy+sP44N9up5ucDeiKKxn//+pybBF1oCVtLM/
PTtItvwiJGXCe2OF+DqRvoaSvvLtnGNFljuBGa66EBQkX3Ucap9HbhyzQiRSxzYy
g9UBIxinFLk4Ey3UMXfNdF3SJzRQrd6Elybx+P6UNSs1PKLYhO6CcIW8YJjLlIkh
r8nvJZhVyb0Uq539EURvu8l8YJDYhNTcnGEV01yZEmuZJ0FV70VWEWN1R9XvedP4
++aUrGth7dpWuvC0r+fwfiHRnwdTgAi8LkF3A2JiVL4LBEXGes87T6p01r7uXqTk
NvK0xiWNKJ9Bj6EzSm+5rPZeQ+GIdaRc7cvwIgo549k7WdFiLp/O0pdCEL7e+6qk
JVmMnNCuT8+8b7Wt/9QIfJygaYhNuIuCc++n6bAq8lP6BKF9FbeFPwC16AIPAwSr
1hb0ncDspzVZJYBAFfY85EFgMvqbcvTAL1q8xCEK8bac54nPI5M6tPwqmJpJ6q/D
nW/xMZpHTAw8FEEB3zfDyL5ns67PvR0PpspP2c/8U7qM+I57qhAHlu+YyG/evliG
kG81tUyROQUu2K+J/ozLvYiuyKA+KsDuv4Vui/zfYYJ2Mt9p0TvhQNCYXK7WuoUv
x+hFSjHBBRwt4eVue1BBeU13gSLuxXMbmNMdT9As9Z7rcMiNF8Z7Nt2h8siwLG/a
GtMTDs0jY+sERMR/LtsAJO/xw85iU/tBMpe8qrDulzgUvgcLJr17DEfEgbII5Jw5
iKFOc7LOzr+8VSYIxEAzwoLpLghgZ3CwaiZP3PRmyA4tEa45bqMcKhqtR148FASM
cUXBfVub14G5ttbB+84fsAG+51HacJHtnIEvwqwQvyLaacH24A7n2GxsWhARz7HB
OWdTfIRfVMgP8AZ4G76jv8I00wma7rofgAFxrxHi0g+Zdw7AOaL0BZY2BsF5unYv
zct94ncyR3m14J9dsMj6V+4dAb8s1mo5FeluybDT0LEjkc2CAKq8q3PFePWEAHZ/
p2tEfu1uBDCBjBL0o+04AszC95HWvhpG2pOi2Poiyt4mpTZP8DBVVjvQ//UBPhhD
SuVEGWRvwwKKnOL4j3gubFhphyCSOylqAatHZ6H3mKa7NLSbpNE50+FmqIgiwXBG
AQx+dJloLaj+ZW6k9Dzhz4pR8lAdtK4dtjjcp6Xqn9ASwfJugdYtD6n048FNd+u1
uuzwpprTZSkNqnD45FAJQawYu7ELnn5+nmdGF48fJ/ny2ZceEaQp88siI+baZNJ3
35HYdjUlh9jxCJgCNsIxwptrcOiEU9gNKBrREb+GwnW48g1fPe98vkGIvy4srItj
o/iFuDi4eyPQNhxI8Om3ECvMVODItt+btchc9WFwM6If0HpQ+OyX7r3O4FMRecVh
k/vVJ2Bbo4eG/nvfAb/c6ipWDppdqzMHJUWNAQpetN39CN1OcpkY6OYFIZQgRBy6
KfFuLViez6We1OY5peEbBOC2Gf4tyI1kV+UFoVJ2/33oRZzzNAlrJsDziZsxaSKR
bFkir/XxY/mcOFEBtfos1u0m1njlOV6ng8Jm6C61gdaVOXX5C9G2BPvtR9+lMFGX
WbL1Q03jM97v5PLfHMzrVgIC3RTpdlHhU5cgSw8fkw63GPo2HZfZeuhBNfQbDLcj
HQ9sNU6S8bIrrYN1963JYvybEd/krmjk5hY0sxJxQijbvW2vpl7LHyVCdne9PzAJ
KBwAAPyMliR5SUKLtFSsYLmX29Wdkcyehoj2IScGJaf7RKuq9CWz3Xiut7RBHp+d
0Luyd/jDydaBy8dlL3Q16AvDd9T3hLSwCDn82/Fi/UCJRCJckrTbHNqteMFmnfwN
IOsu3ZIih/ygimB0VTBE9bFAaImh2lNIms8Y9v6uRx27cd5Ji3CA/jRfPgQ8vlXq
0ruk+QMFypSm8raZ8kwd27l98loqCve2XxkgocwQRL3WzRALq0/yyxaTgOdwQZdn
TZsyn6ICHYgaawu4JX14h5BrWGIbcwhaXM+I2R3dL9fF0Lt/LmwPkqCO5qNL6lbu
pZBDsHnZRAlDcX+ThjBh1KGSEgrvnMBDb/WFBfDhBIP1qhTIzG+M/eLzyhSF+qaf
I7Kv3GTIAzMNy1s1XT9wFrGlJZLnU+vXK7Z39wlIQ/OeIcPr+JUbrbe4F6qTRpD1
ABvIzxcdGsr3hoSgKd2D420VvEyrFMLqna7jXY8/hIkN0COAESWHfIcXuhzck7hg
FXlv7gJwygUYhvBzFehcChcTD6hO7qEw6j3NPzo9mYhVBBsC+sG4Eq8sd9BDRRzM
m6i+4F/LIX20fMmjlUHH+/BbHE+UAA7l8SBK5ph/cZVsgt2KfT7K+CoaXY2ojDei
npTksmVSDNe9U84cvlbIDwmoSS7HF5oydlC3L22zQsTmU2sVn7gnEYhyaFk01JrF
xxdB8jUAMixR99W3wU8iwNAMxn3SH8sIJ6UuGwgzMYTG5X7TD31bZ/fmES8q4pXj
LtJI6NUQvOxxFeZOEioO1DGu1+l5kVfrQfYs8r0bLwVgCi4k7Jcy1pzXP8s4R/Cb
KZ6OoxcID5TQmUYuOG2b3c1/SPMjHDdp/9EK0VBwMI/G4leZT21NRh217Rt8OqtX
JykQ9Uqm8PhfHhHYKC2ovwomkAtukLmxSHHmT2/xxfmFp6MDkTdZXG0sIwKikUTl
5VUrNOusD2o60KOKQ/kPwWz87gf/nu27SZJH/L9BIh3bMbvrmDSYvzFUSSAQ1Cy4
F2WhfQUYrJoJrmiJiDJ6OTzaFfe809gZH8M2SGr/wKkXmmI+NzGUkgJQfanpimHI
Itdr/yRLvMPJXyIrxNiPByCRVk43jcFRaqZ/DTMm0RNqHFVbF9n7d4N8IN72tDbF
759fU7hfUxXhtdXZBjs58FdDjpBEy02H88UoMZEPABE0kjgIXuHDWGg9dXffzD+X
n/jGolmobDGz1ec85NmASU5FiPOb0X1D640RPGRXdo6AIANWgr3D+byb/I3c+OlK
KzfuYNw+vL4hVlMPC/Q9HG6VZ1lp5CDV6jjwvt1Vm5y0Ok34mJJb1uI6enu+FeDS
GX7/JlqcsK6hj4B44iKN8mV8pb2JYH0vgrTMvHn/r7KIT0eniZuxJhckFRh+Xulr
o2EOucYEx8Hn9ON+Vn/9fcrmHyWbyub0PGLQm++ek8MWTcZjDojQ/UpLzW0Lox0z
36zLES2ky3xJ4siXaSx3d9hqSRRFMACy7b7oZ4IPaP7sgYThyI0m9aB0HpF1NGRw
P0gg4/GrRtlsj+rCJf+NPOMTuAoLz1GZ4HKUZE85OP2I14P09hMxe1kIoYsS9hef
PKIIfJKY4RZamdn7lIUA3cJYzUwTfoY6jC3UD0IiLk669nPYvjjzqtjIAJ0cB+v8
WZVKDA1JrxmmIbCOdesshJvd8eR1p1LnAHrNaEU7utpgMocfGLMlBcGOyG8Ux7aj
tLJzAtUicHddq0qlvBGn3f+ApLXrk86FJ2CdSvaOV9tb9PAMLXEwm3Q4C4zTYBuJ
YXBBPJ8eIlrZNcBSUBZFDxnj/tzYDu3D6FbUUiBpxiOxLXvhrrIE9KFgyw7f7KrG
Deo66J1zQ3Bjnivrqz3iDSxKJ10o61ZTjGUoTj8XF0LRMk2Q3IOpiBJwJUjsK2DK
1gvX+l+rqlg/1vmIPvGD+njKpQ4Oi32Xxno6205htGR8ZPfWxPUioUae1qa+jfFM
J+YG4HnZHQNy7fXGAn3WWgMbodXdYo7JrJUsJ13eEEiRnfjm76scIPBknxVp4gVN
nOa4/J2Y+JZpFJVE23DXgS7RYP6X2VmkMsfIkHpfHt0LtwmbTB23RbKa88IahGyw
gVKmN5wNgyG0qVJmRRMVnrMeSuuFPHrIP5BgSV1Ryn5gM8J7IuAd9oya3vCSYmpG
hz8cdIOgGYOqZOLqO7IaoS4MI2tQNHdp0Y8phvV1FWhM5qB+ygdAcCjTSBx3kFf3
xRs3MXzngqKKpT/A4PFUotd5kttgIZMCwOVfdO8VRUHNSO71WEhBDirrcTkcdROi
OeLopOwu+4nzIiNF3o9NldzpCV99Av9wcjAwxm4bAuYTeTrwSl8DmywcFreBDVJ2
9naztVdIE5MhPFaanOiJ5GIB8yL/Q0sDyX3ClC58onjqwgDbS1XPEll712AE8OwH
0bhXgBOZxfWEaOypF0DUVTmsWPwXEa8eHKMh6ik5PmHYcVixTJsngq3dtfBk9IK2
OLWf84TH9ISb/uBrA0ATvp9nnbWKTK++JdjRh2F2sR0I8PBV8KWjFa9d1ZoAzGUA
xU61Mkub2OLxQ9ucqcD5wo0pjCP8Y5LTiFSj5xA/GNiQyZo4LM0nYizvvgyeRW5O
tmI+OdzrwtCgD3bWozd74UFc6z1VJCNU+Tro4POSox5esUpF6zIzST3USSE5VHbZ
DiJAPL8UtmSt6i0d3ZLFPl+/GzF8GS/3kSvktMCyL4c0nduTR3u2D8CvCs+sg6n4
iWEvIXdALcohJEhsPoV5DiX0v6BcfJVSqHJlpARNcsJZNCX7t+Va+RmZZIqStjsu
FVMoQtWOfXBB11YtrPhOB4p0tQF6i7fIX79IX9MiC9Twt0hyYYtKhOuOu2+7zgaR
5BwrfTO6z8lfV9TJXhp+f8cgcZjAa3R/R8EJbio/BfAXE5nYgfO0OpswfCxHK0l8
TWoR/7hWovTe0H2sokDyhhgqfUihjKaSwTUkFVBlqiChI6vXjXezbT3afErN44c9
Ve1s1MZciVwZeQGOqBkUEL7tIqFac5fHUBW2C2IRIOIbzJr/3CFPc4yHlUEd4nrU
DTZlAkHAIvFncnhAENZmIwY9c0GKdaLMTzfEXPSnAP8DoWa3CVOYjcaqG3hQk9IG
UI9mqL3mMwnO4L1YBvmb89IduV0+r9qJbQDMFjgSIkNXMVJFngef9wHEzmHnLJuJ
bakYqExj5kXPyFfA20Y0P7Lci3Ev20u9vbQnqzftVLTho8RVn5FK63jkGd89+JYN
TjJhzeaSPHApxwaI/Z1kruA69t58DCyiG7DlNOdpEu1n1q2qt8IGMW7LLcV9xboy
Z+zYbtiUoIkFgO6gz6vDtSU9wNV4rB2r2ll3H6wS6qO/DR7v+awY7wyGn/EoEfvp
EMyd+pyFsilyApqCJZOZZyTB/Ngns0RdiGWtmK9rLK0kR4W826QaN9La6u4lpTJp
k2wRSF3+J5QTc49idysmF7niM3lmw24y9Vyd9lAfevn/Ci2Qp4Mek5i2zX6OtTpf
fLZphPUUGbdXUXMyPMWFN+sYf37ZuxzGef9B4xxWHxE2KjjV94bJJcG8WtDKASvf
YmuSoXFRUh7nYF9nQjUyo0DXtGi2qvjwrB7WdDTs4px0lPvq/Psc4XB95ghfYzs6
jARwpwgweVMDDXVMrtZNoGBly95HHopQGLtaLvRJbbiv/49bptbm7ORNJzTF6uuz
UcXtt7ORUvJb4ieZUR8+8QT4/EmMr8rLwD09skelejFk1YPoz0iVFQDTZibVCj6B
yMwlTy8xrt9KoDGjar99cb4dAKQQEOEOnj8Cl88qs5dtzppa6U7bUZm5l5LYtUkd
pLsNgJXOpF5NPsK8qzLjR2/cBPrEA/rBvlK0g1TcbIJBZy7djNJUx5SWaRc5iJQq
7dll3Q1A8dSjSxUkue8KeGTwhSkXb4ALzhQ2Eo6TGp2aEULqiW9fIHur3DC5wGil
6vzcb0zuvlZyvAh1zOOIhV+p/iRmFQI5R9xrDxYXr7G/TB5T64y7U/O21sqw7lgR
HPE3rPr1ACMvVaDVU4yrVa0YyT0iA5PM4A9HnrPaDB0J+S+mZnORBHIAOSofdz4W
RMaDjGWjcjePDigKxoTJbz8p6RgYl95fjX2GBvC++M0E5yf0XxpSe3v53xWIasXn
bBGbOxrfrBeHhGOmBGb1b3IjAgePyp57CEHpMeh5sPzgWw4xWw6BEjz2uvGSR3U0
SO1rnc4EatDDa9SChG84JEf6GAIzdeofvETRBYJGPl6Tf9ktJ272HDh/Y8lBrsGE
bjz2bQ3V4mONX2MsOetXMSCUirHHiEwyT4RWxALuNnNIy+3/bTN+gFxJzGeuweYe
gbqNpXqKN09IIbfhEIu2U69+mVjd8Dv6AA6nJqBKA8w0AzjwCPqCGi/lLkDLzpO3
9MmaFK5xxO1ki2Ys/wz2fvgt0IApzx7mADQJk7ldhjNWQjIz5/+IEkQnkMwh9Fyi
v3DeQ1utFHds+2mWPFmZTCjlwsCCO9hqhKUROajMTjY2pVyBPTlGKhhEtuBfMfep
HxSy534sOCIGNU7X5Bm7pQiNP5oDUEktjPk/2Jw/jgjtL7PlEbk49MPv9dH5O8Qz
ZxVcNzJ4Dc5KcpsCUBqMjLfhBIDOJLB9x9Ae9YzmkomxgilmvTDyfqE8iI6k+Tan
zF2r+WgUGGp58ws7doTGkrV05LshTbTN/5w4jgHyRrc6JEZdW2dgyBJQtPXHX711
t2mQfTu0iry5AVkhvGJgenhcarRCCZilmSzDTS/Gah5cmP201XcF9EADmeqMcbnX
UG4uWMmqwie6mSWOVhGfmmtEp8xisQoFwMIw1qcZXkR25MVgEZdbh37YcB5Oh4Yk
iqpr6hbNY/WQV7pqDA97dIa/wQFciNFcfa5cn6LoTBHkT/dd7fhJB81GqtWMcxb4
fcSx4Og0xElT003oW9Rzcu61elSTHNR0WuZO9WcoS4flMAjI1O++zC/EsgK6d/rA
GcjbiAvqyLRHdkAryxz04hSsFkjKfYnaNy7crQFwt/GjTtW1Iqw7c3K0/vGdSFkz
2XNFonRiAZDwBXVtKmkox57Yp0THIcPxzqHZ88CpUZH/f2usVF0vYj8n/0BVIZzn
w4cEwL7hy7Jh8ApBm+8KeJfaw1aieRNPcppLhf9QUI1f5YUbWyWlA6J8FVYBcv8E
n8tOmMJDEatMXu48kyqsdW3CWO/vYJyMvDx7t+/ZqIY+UKTGuuGCTAM/ilO+CEQf
LGTTSRQglnOD2CH4hmFVvHmQELK05m8W+PwqiAvrnnE3wBUSbX7wZLx+3vuDq4Lc
kOAgzkvBI6yvB4YlUVQzz/QgodV+M+jjd5AtDUPm52esw0sM9vBUHn0L5N7GmOtL
ajJWka/BEBNX2jQ2OLgBuFQJQuQywgOQWXP+6045nEgJeAXOFESzfJ2QjkfybFKA
720V/eUBTAfZ6Bfsdx37DT/yfdU1EFjKmYI0pkhYRRydGWu9IhFPV7aJLmx+RE+1
xLFkezcZaiv1/3Ad96ptZyDHrqAkWPacYkkaMRDHXQpesAML9qupZEo+nm36Z1UI
X01gZ60GVl5x5WA/Iw3aGhMFXMH8SoXsfVNqlX3aXUHZduzXBQ+OPldFJzx1P+Au
kNs2s0A0alNsp+LrGBBdevEdLtDDLFJalA44jhf/jmweQmqdatiehh2bEohTiljW
yUt/kISsl9PMLLyWUHe0aoF+zCbel/crqP7d14AVuuSOOeeYpHhTTQxZIabwsEdg
39KfOE+YZhu1K+oEv3xfmwWAvapFQCqLM1tO4idJYk52NZVcqeMR7xTw9luIFZUK
HtNhdtivGTPgjqOHWEm/r9iR24+/nmEJtsGqeq3M93zpfxUgbUwYWVIwvSQEzXDv
yl7vmB0yF+5M6v6HYfQD+NGJ4clCk42WkolUnDSNoPvmXkcAotKca2UolOVprkSP
DAy8nRU3pLw/v2HhAOtBlwV1KwTh+Twcn3xSfaz0tfNPihm10v8lwgHS/4xNGsPh
01T4zF1gKtbM7wciZMRwKFAW1ugiOCDaEAguvxtO2WdlzRRweratunzsWrrX7SJa
yQGDEmrspsyk0tia85Aj1yodYqL6+fFRa8rRXWjrDozEfOtVk+XT0sZM+8UW7tXq
9DlgIRsBVrfO7v020kl2osBRiQCDOvb5DDRkXlieKFifKW3Vs4FrF9RE8fwYYOa7
eZkiER8MPddBxQc4eKj2dflUWkuKQKs1JtzQEELaQFtidE7iYtFvt9QUpdPyi3mq
NUHhGjr3ndE+oMgwThHNUri4JBb3G77bjFPjbRYBKJTGrasfrc6MEJAG6//8Ajfl
IHsep9WabgjALNDCF0X4+m2Os1QDa8PqwQZbVsUV2RHbXD+hXc375cZwl3a87kP+
mo0/uLs0y4C/W4WaSPNYdF7jbz1hn5V36cJGa6j9mHUbIMiZ9ZZM0eossWudkxZs
StR3U2P9QDtMzzXefFW5k74Yl/aZEEFfuhuL2jYr8dy1OA66QWbjEnjZsnXJjlZf
3tyFpSe/1HMsCon/oFE6wRSiVHORfMm52cRBlmlxa0isr6fRJwpOwT1GCHaqBram
FDnDkQYF8Zba9xKV62i0m/GXdXZlZGW9EQxfbNmz8zi1Zb6jQQILg6Lep9C00Ed2
ctbSdZza8G6WAP6muDL11R8xwRm74cO4w19fG15GEzvAWHn2zvKrYoK7XC8a3EGJ
wWtDMYA3ADAcRYRaJ9OwnGhmVvDmQopn3A1mKtAsd3KsXlrIrLEBzQdmdLe6fjCp
Zqb6C2ctKwe96lS634GENfa7lMMig+NBlRPkLr5G0YOTnyR21VtjdvBgtHZ4ijMQ
t+DuLKohxYudEJwvDg0JBTyLeBNmz94XzSacFPCV1IUxEJRL8ddrkv5vxXuquGA0
kBN0Rw/eq7EPJw/+GeONpBCGqbNPwIkIR6/Oa3fUAoX4BfCAx9C9+UyBpLRz9Cuu
RtnC4WQyQ6/2wpqpIsN59BhwUaXjxZYAVKzLfJ69YVqbgi0mXn9XPX2NlxUvm9oE
zzuWrnj+9glI/FKU7X9Oi9xUgdw+EC7/VJpMBpUpGJ16kO5vT/TlBXlnWVyqX3QH
dUosmFhuUOue8Ov8l972CGRW/pNC0hDcaJx+LphRhsjbGi0TdaIxvpmjv0DelBPj
822dFI76+PYNxl3rTrAHy685GZBDvwbkzftr8PTYpEsv4JH2ksddp1FOduYgMz/U
FLp0bdeoQcddSbA+kSNuRQFCq3UNMubuzHa6QROVWWn447nbNUW/8kEEK2BgJFDk
qfJ/8VmVpDeQ1prOLJ2jtZremjXbdqdKbXYpFt75RNO74JoEOizxnEBR0dLdrIxT
FdjZuIGvDBPXs95Pk/EUoXDw0+fGV89wTJQ/19x7Ct7DT9y0So6hOPpXo8wrm6KW
BwSn0C+zCpt2TSsHpDCk2ZGw0vGxZtn8DDMjz7/ulAVSLCwR2mJro+L23BA196xv
2LIKBWe0JjQB2bC/DuSMmgWD3bxqziLixE8lUwoU1tmeL4zZhGG5CVQUFBALiwkM
UFzFDk/0NuFODp04JF35t42y0IjHLX7TZV0LF97MQqvdOJM60Pww/pTMcrrY2qvh
+y7ZHnIadsKTknDvMPl7cZyo7k5K5NGTHHw327awKwlP8eLX9xV8zFsEcYVjuO3f
9aF9a5ZZi8uy9c2Sg2VC6NkLZAwuPvIEBjAuu75/18wWqbUKNbJF0wtCVjq+W1Mk
pybZKSqMiV79o3q9JXqXs4hhXuVuFrT67Vk6XFmFo49nhMlHBHu/tOTMcKAfaGGS
cu6Lpe97f5Pf8go4RBKehj8lmvQsXxNsvq8AwOBTNHsI9EboFCsM6lfjByOVqVw3
zBXdutbSbR/WyvKgkFFKZNX7qMZ6+cASMYoqxeVuWizVNUmcGIKANE2nd6gBQsGR
PI9erUP1q5pDFqozyF8Eo/2Q7GlhZ1OTQjItdz+gL86MbVHqEe7bP2PlIFfOUINI
NwlkRNEtqvz3HQUUpw7o8jIHQcplqLGZvq0kQezpX/c7dNEZb4xhz0kwG9u8o9X/
f+e7oA4YgQ04vIHq6+NVl4tFjs/sIO6AJnoO/3zU3q8lxWbCCB2duzbXVg/UCL12
1UsbQmBU29O5ZddxAKg/0MsbofTjDSBiW5DychlsNlMny8+EoXAQlOce80m9/zKT
TIKCPDjGmykrhDb6/Md/N/uCJ/PQZpxrNmptapJmUDMTWg4QYQxUc7G0ba18Ox04
YOoTpY+W7NwBkRV/xdhKZdiW4/C75HheIvolvkCPvoDhekr9TZUX1Fm+qo0KmPoA
FnXeDXCoT0mNaV9nZxHwBA5mkaqz7UpriHKjOl8uJScfXyUCdpteOAph0+/7zeWJ
+XPR1cgOllGfcneg3B1V/zjqewW8BShAj7qJnxWMn6XOqXewxx6jNrsmEvy3wrgV
/iPzOGR7GlrNRLJnzw8/UyEBAvBxmpbZRyCZjRp291aa+vrg2ks3OVcxT1lLGu8m
D9qdNrsx/7IbkhyIYF1mT+Zl0ROsyj50yYbqxNRFv9JDIcyRJr1gcUDL5++A9Mhr
/BojMmFs4fx6HDLpniJXKh+2kkT7w8hcnZ3aY3veLc3LAg1mTRx3nA2/onzLXYuZ
giNKlVEl+O4v1nmba9A6HHdGWEZ0EMVocYjRmfeukCj9bNnwsAGYprN4R3vXCFQz
x0heLx683k+QMY7KB6Fmqo52mv+vnMfvHTOIuUPNIzyDlvhUSxohSOUy3u3AMA9R
iW0Up2oa38jWhVfVglH/QzRJDlTi5EQNlCesvuDytrUvRe/FjCYGsYB4AJOkmRLC
GSNOzpCoan/T/hPAcM2WHK9yWuv31A67C9820hr2CMGA8U6hdGzNTbJbg68DxrRl
WpS0CRh5m2GLM59AWKiuJ9fr8ZjyQkWmBXs/jea/gD/6+NzhqFei5dkHLyYXPBpI
TNSuFhuAI5n9PfZP7jg3LVJdtNZQVv+seysHleXHRAEYeIKhT4oEWY0ohZtG8rdC
qFEB/JIQrhI5G6LVuvcIQqBd26IF9fVDxfQMEvFLix1tjHgy0rbRRqfQfVtamkuJ
repeAwqvLNjT8RWZzxbc4o3/MlHg0k33D3WsXEIH3NK761Z8wRhBkQ1cpUcMMrIu
P0EngZCywGTYsEv2PLB1+oA9Y3Rn+bhBNbeUti1kfuZMTBcV6LGE+sx80uOVZdbU
foXQkAnVndres6ZxT8ecIBFCaUC71zvcnSxOmW/Up2CNC8nCkdn3jPvm0dFGSd5P
sYGb4tWHVk27HSt/YhlUcNd6qQ4fqQNk02YY0cM7pDi0asFz/AVFMYF+u5zwSDTG
UqKxajgffCvtZpIvYJk/eyUaTT1gCHoOp8RFWbGS5Fm6zWIFp+KjQGt8TcxNh39w
ksxCwxAG1Eh7AY+uiz3+eDZE0b5c61vVmFsd+bZPKSgJvCBXcYzjcTQs4WdIFQxy
izlajKPTuuot/K4Cv7/5XobPeCB2aWjMbASrXXM2tZgvBWWSLetSQIWx6Jkp+DkD
TqdnrlNbHNtcFTwLoluF4YSABnTsF0OLJj9iE3TurT4+VgOPUJ0bOcSNl2EWjgmx
EN12oOTM7wuUon3MBm952pnc16koTm7Ewi0a+O7Y8q/O74eFyUS4dOZvW1Z4KcnE
kgK+jy4bn2ziMZ63SQxvyjBRXpG3bwpj8URCTuaQvvQCSNrFy6uGUvLbhAtE/IIp
8PwQlLccBJqzU/wnP/QKYiCZKZK1PYUTbSXKhKHG/WbpVFHPiV5NIgnsk+5wRjQI
zT0pE/qZxvLtslyITsPEVtOq+IM8iAud0sxs8NhMGV/XlRCZQDJDZ1ZDXSqXzx85
SteUlLea7vbtWZgTp2IZgw5CxXwznJwoM4eFmuT2pJBT+23ErapOt8zRgdCIVpUc
VSbla4GpTQN5hRQqzAaXL+wIucU9IvfRC/Xaj80DRKpryGKFKfdvbuQoPsgGb1aO
sXTzKWoUzWq9kBuwKmhZihRMmCMUhvtVr+ndJzRXJDI15JVED3OQrNKlfmTuII1H
SMKGxxx592kuYDHjx2nvD3KU82PAf58ViPHznXEIO5Sb/t24GjsFS67w23kKtBHL
krIv9+fxbJGArLEHqrbSgyQaiVVgYHYZcxfa6rp9vXL7v3gwfHVVp/V7FJZq9f3m
aYLDBxEGmX3ao9qa97UpIAJQB123UNCXacjCCEvgMSN1oq2RXB+6bSiyKNff+ZCi
ubkz14AcPyCRZ9dPeEgid6qowcsad4ADxrUEyuZB9+BMSbsrVIm/p6+sEZt3wior
vk1rphd5f4+9rmRf7K1WmsMriI/CnS5QpgGUqa+yActIhTO5ZwNIbqzbMd02wjZP
E3yFDn848Fgyi8CSIexa1oYG51Pw2AguVALNtneGaJs8salQguJYx5zcpzCK+1Fl
Xxy9Ko3nMJQi/+qNf9GR58kjoL15ra/9Y46dz0nlif2v5mHGzc2niGcwoFU22Rww
WTLX6zSFMuhBFAeXbKTPF0VJPjVfT8J3h4frPp55tXJF9VfcgNy5HxWtqHsyV0Zy
ogiRJOZcLjdcIUSthmwHnaQ3TEU+wzodND8Ek07dq+UDLoIzCHmdPEC07zqy8u2k
fmpqdTHgjOoyUfL3L2SyGh3g23AvhyK64lpdfLqNgHK/19yM849cEHo08kR2l8Rz
6k25MjfpoAB+cF84hDJiYY5cBzb4XZ/Wz6zR1yNPnuP/ibaU3qbUvd86KNmbcqy2
L93QCn9UiCQy0HRVEnQRZXX5OieY1L0hv0PIKsVhlodabSbpl6MY3HNXzNTP/S9g
UdFtYrxeUJyqtLYghAP8ungPmTw16BOVhnbOj2AEG1VaRBeMSUSJFxjgNOXYh5de
Dis5/Ovb5GlwAe3LYfQuJ0TdgB+acOWNTUTbDosDyYWLUINF+V11hai9UHswA+kB
sYahn3ZeKhQg9VxkGES6Hh/4xRa0+hPP6XFySt8drr5mDSi0NDeEthRpRbiY4h27
FSSaFn1ReiO2SFSniOKgdr2EvREajMDisRJJbpFgM6odfyTJc40+ilSeMaI3jKlc
Yl4e34KmJjJ3dA2+CuUqtYomERKokIX6gFW7KJ5lK7tgsy6/Bmu+W1RK9nxfSIfv
O4B6bpkj6+L7E4Lsn8Hzl4MbW66lKREBvCiL/TZXaug03nLD/ozEso35HQpyYuya
v/FTFlBe5cQprQPvQ5PjMvT+WyuDMP6Sm09RdJ4kGGJVA/GM/K2CnS1ZaIJA75DM
sPF3ZF8LhZdOG68dVyhBKmfnIUY7WNzmPM9UubWDYouNQRJZj9m4WhEi9aTWwnNY
KnnugTRHbYnxDAQ66xYoWWIalLvqYKNTyBKZulYizKBUD6pU6QLuxoU0PFu3JmG1
CSubbfmTlggSPgt7i8YESHhxiQy0DTgZ0bkMaHfs8rFaMsCRuMhgVHd6yhIl8azz
JW4NeeM+yIH/Z8IZ6XhhpoiHLmJymj8ow8iftatrDx/6wkzrJgIVbrcALpxWW8YT
uXA4G9LsKcg+7gd2FbX0qIauRtHaPNHeKWHY5XFmritl9s1+1o5TVt4rOfSYIH6m
vTY0T/6EHZZksPkGtITNYESTTFLaPq7jE4sDN3Wt5469M8vFNM8aPJbgSAYqNkCY
zhforqYKYhpmqvYIqwP8w+GOhZbmqn3qvCFUNm1oV1CTBpnedRauSHxm5ibF9N7l
ZaVWF9QwALTKaq2YLy4+j+bNp4zctoYSw9nQP+Ks5iSPUJpodmYQ8QWysneapckH
+97E8LikD9+DAz2MU9NJktgLi6sE4Mpv1XnfbLwBIsk+CSLST6m+of+9yy9ag5GP
DrHGFKZ9kb3dBePvRSKMhU4pAhlRKS0Yccu+IVeP7xd0iYYuHofT1Fc9tJu4m0V/
Qxw6TJt8aVrX21QF+WP5y5aDbodVLxMMWAel+DMfYedWoiWhIgbrSSp+exqYydXb
gdNQPakS2XqeiWlSimmtGczkkHhbtEYyW4lBJV8hQ3mlFCe7LGcncxbQH3M7FsnO
I9EzSH84FhlA01HFvlhZOTdrr1sYarWKtxH5VqGE2UcmDQNnpjPu0s1CvqaBcvTC
ekLhWFFRD4hfITOJjg0tWaofhNZsw+wopC+tymNK0pPCu08vshRWQ/9ODXBARdb3
31NNNzGm3DyIhJ+A573rTeq1v7hYzDWp9nRTvFztzG0p4f8I8/RSdFgS/Yh9TDKj
pnuNmHvpaRqbsgt3NfIA63VMXbUJlKwQf3hUGv57Cp/ZZapeyzW7R7e6HTYUDoPd
1WT76sInPHBsZVP1QKG5NbRqXcjSNcZUtadd0sL8NDHmYPZbndd0ZEYV6LqX9ySO
kRcsifazH4AY9JpTvvutOieBRAniXGJcgBfYDCvR0oxYHEI4vIKBSq4uW+cRWTDK
5DtuFSj7RjpdGILy6uAxXZ+6DLBwglu/EWkcEBVuymZMEQid03Ezt0I1Xf1UxZgX
f3/iwKlU3y5+qlxv6le5nEKYp8M2uxBbF8N8hBBvlFWaUsQB4sS6nDE5z204JPnV
VTybdWz4bALTWAIh2+W78lz1zs/ce6YBkV5L81impyRtPPpocIvHcY2hz9pQ7ShM
gUtyCPjoEW4uiXA6I9SEse2KwEimdmmsyMTia8beyHxrKz/XH4LJ+z+Csw0xUUie
ATx0JO8njtlV0zmsQOqnY7j+Ugbeq/ojAwNsecSTsFyWm1WnNYw9QI6df1pn6rUJ
A0tVr3g+4Zw/645ebHdYMBT/mlRy4B5lTASLAiwGzp19rostEKZDdE7cJI4IFB5A
jZ9pK2XktAWTkQukG4zl/6MtK3Xt80L/Vbvi2RgkhPtlmvs9614+l5HBB7Zy+7XA
ArivgRaHNuo6BxOteIps1tWj+ZxcHQKf01HmpWg3RcftJ/c766MhnhLPOEfH0ke6
86EKieOz4DS7LNOEj/H4y8wO5mTRCXlrqVR2fodJeh9FwMm1uFNkNs0eF0gtOTRC
YYO7T8z4qDxgzXb4sz9W20mUNrH2fjNovwnEXmZBcvofDPBZRLG40O2P6FGeaocb
oPNq7YQGXnBst+Z1ulF3VtkvjGaduQyxJx+9ObtWJss0d0oqW7H8YJ+Gtn5pgTGC
6lMMKcA9ImHdRtmEg1NStWMNsruq96Xz7WXFX/pazJGNNyFLb0RAz9fnnVBhqMME
GT7gvxHt3uXSSHy9P2NjSgdtsVMoUP4Gl8F115xDwO5yMcFNwkaEysRRTkqFff0R
lC8eYyN61GpmKLAZc5bUrSZyitrW5FrG9tecbMp4M/raogb4kH/0rFuUzAZp3Dt6
q1UV5u5wSVxXT567OU+sGKBFxsetKPAMtyEItmURFudSUnZZwMwwK4B0wrbDgsvq
IIB/WoHy0ZPnOdhpTMMIeXJEynRH12lug7d6olkvvIb37Bp+JeVW6kPxYdEWNtXs
mCBbksQYQ721Hnmbw6as3DYOfY5aUlAtpUeuI17vChSynAtEYwBwqKtJtApfipko
4aANkPIMr2cO2juD9KU5wYcVYKmsgKemnkRtTY5JmSaTgFNgh9RNzqsDT3tHNGUv
4uz9Rbg9QBaeTp3C5b5kM62iJkk4MS762Q8L72PN/lt9YlNANdxLVHS+0WkMlICW
4MEhlW2r+5DhyIalH5tnRSmqYnrvm3uaVy6muMC/IyAIrwII82wCAmrJcbcRgTP/
lj2FaAoJnSurVkbi4y4G72oHTR8M8NOnv2vVNxbCQAkqE4EqnSNyOQnYm5hPrhhK
ISD/20KC2OICA8rqP5l5d2yHsiFT4ynAxrtK1BAMbYRoc/SfU2p9DE+Q2rcFjhQ+
9vJvXk07TK+uKRcsu1uaGTX/drhBMsRzasITPOptNBYPAW4XBCBLD8D9zDLKAmLQ
IqUS1J7lE80KbSoF1FVLiDbaNqtzCOF9YmCaQgO/Fdczleq84Juvy25R9/fDB2t2
gUPgdzCmr50NVpFeg/wHrqtDEzU4m/6GSTcSL+EekgX2Y8d+Qq72Rz92Bt60Mncd
9IxuMwSDhbNa9AzPvEor5fV0wQb100Dz7fNEqmvQhxT5WOUavVmJ4leqzud6oKwW
Vx8si/wm21h7WI/Adiepcnq2zDN+TGW5oRNBNHHjQ+jveHnxRh7PehWvj4D2mlBT
rxAmOBuiM0K6T61QJeEn0snASiWeQ9P3PG09lMvpFT3HCrJ7ldxvRPSRrMwFKJ4h
HFwObnaAVqP806zn4E72i7e02kQmZspY6QmBNEFbaChvVjxg5uo/1Hta/cR6GbrX
4rMBZn7YmrFnF8kAj3DP6fnqE73H4ZZgv8LpfiOLoVIprhn/2MFCkvkWbBdyq3bE
2Bqi+OpR+4fXKrrpF5IaooZ1Gu+NTaeufk+Tl2zVMXnF7Hq4STxSUc7hGq8Lybil
r1q7OL36J97e6mwNEX48Mc4rU5qQ3e+JxDz43QbhZSSTuLNLbrcmK5Q/8lJMlAa0
USX7SGIR+uy/jqm9eTOFw2dSWuwxzeUzADTbJoePi22zzwjfZwWjQYtVq9sTGm9O
yCQOUnjF6v+tWMrx1er5JwUysyn+PCRUTzrOcctifKMe3XRqvw7Cd2KYP7URHL+F
P1Urz3750rrA+Q5G0NoJXRLDi30P5VX55SZpTBH0qFHfyRU8Iu5MlFmLbBnRSfvU
yQZ7xJhnxQr8Wg6uh4Y+NgmSbXSiq3hlhsv9eutUsQM446smgBMEG0RUCuvAMjv7
cA6LWrgDIQ9uLZ8MHRyfHWX6iU7wuUo3DubOYA5YYOR3bczhLGMyfuGUmpoVfhoo
iAushpCb+up8sTf604OEjJpFKCRwoLN7JLh579RB7YF7yjpOQj8lbeTBvg0pT43L
riL7ydExn1WXIETaDzaikl1X6F9rHv5ejFXYHrlIpC65Zeq4XFecY4adoVYTagqh
5YV0RfRwl2Ctjt4xfZUO3wBpqpDh6Z6Dt50rN24h8vusD4WzlME1aNyMoUZmA0U2
WBbXTRHhIlgENRGowTKdGuQ03o+2tkG3owtCqLU86eNNyZ/trCDrZOW9m7TNel+F
yghoYCZs14i3q2rzhBGr0Bdy4WIVG2xKDtTb13UsVtNBvzKBPLsk0bOX7hkeXcbP
iKrtIVts5YYywEFAtYY9ou4cvX3bky8E9YVBCKI0qUFPok4yXaC7NHvvE38c6mEL
iN+zaCo544i36Ci7P/vxk1wtPMpcrOouQogOK0VftiC/db4F8BPqqRpPoRG4lWQb
zv5SG2RmUL7Y/u7cfuPqv8Ow7g8WgJ/eHv/S5YktroL/1yzAu+E2aNP5OhfXEZ3f
kopj/8tpRtM48oeLCwH28K/y8E5/fAADhJV8s5qPrKqS4KiF2Nufd5FJtVXo6Xlh
llvWzHMpfJM58huOPWkzgz31la7YW+tInsqs2lA/AxpozvoX8hFod4dzkDdwaj2f
06lGLx5+bXfiLeln9PIUpJsLGB/FsWD1+G22KT9L+EqtY6iZVC4xCKqwRciEcrDK
eU588k8XvSMkfSmtc2l5j6Vyqkng9Fj0PEMXCkyUwwlqRevWrU8IIU6R4U1SmMKf
7tjeUgCzK6RkB6rD0OrLiYz3Ei0uNKbd3vWGohfwixr2y+5epzb6K0u65MT8v1wf
pnIz0xYoG+oEbPiMmTW2vi5M0dIptX+gZFgAVf8f+97NNYI9iZHRIA/FQv6/ef7F
ri+vBaiqrXqJvzjGvdSsTi+XACIBYd2aanuH1s2IwxTNAac7tu9Umcpt89MwknMf
1rMR4HaKxwtVshveYdBaJcgqLXlxe1mZLx6SVNxiwEqzKEcABbbE5AN0baxGlp3y
OUso3rhmcJHvBkCePA4Y6wJMD9LhyGA3QFVkKEt2ubEDIj6+SAtzjLliw93KXkR0
gQAVa9tc01fojHwRanJod+coprynHPknXWef22fda3291/0XNcsS8wBOlAzw2/b5
lA3FG+CypWgg1cdxuv0W87m8Dqb95xhTy5Dp9tdgkWnrKad5XsisAh50UERk9yq/
rOVyt9WLzAB+jqOw/rVydkctJTsHaPTs80SuAc3iQRC8/HSrnqT2dYFk3mrzQRLU
nX5E1JHdFR73ZMqVo24v0DMOMzZJEA9KZOzztRV3VVP9EK8+INR8Tt+RsHxAR1En
qYk/Sm2rQ2tHKTYUMlU6IiZQ9ZpdBjwrnmUsM94xfiA7/ke/TVCjAJ8xtskEmfhN
rg0IUlxNwiEQKYbPFbvP8Fb1u72N2zvM4faO+llfoH4bIw18OVTfC9H5xrFpG9NL
pVfxcozi0Hq18te8fAup+yJaEcic45wpbWcoYK3S5/X+VF7sl+Xte/AFkzDzemUl
vs4UfkulEtCA480jBLrnTGE1XDsKsp2zA1p6DXgENEXpp5fT3I8+H4i4OYca8Al7
C5Q5Q/gjnTxHeYxXViNsnjYbJh0laMkcl5tNJ8mdtbyZs9kKV1dAHRu2kbXf13kP
mJbemXrf0ktfHCCNba8eGJEJ3TQwzUbU1RQ7MZOY66m7J4+gqwXZGUvd0divIVfB
dG5W/JqXhLDhC8cVqNgS7+OBzPZo6IMMgLKX1xGtDMSHB8YR7Dn6zWq7fy4eqivc
vN/GxQn76I6DZKI46gqsUqlmYVcYO3kAf7ljMIL3D05I46hGSjRie1eaxFwdL7p5
yz/TgClTcUdl0Cle9ClX97fwEpBMNiHwy47JLGQXYJUeR9eWLooZ1CUCYELPBqvt
E5ZjwbARgdPBQCXfAaNlP39ZfeVbl+YbvvIh9wPlZ4Kvrb14d3vIOhYjjdJ+nH6s
GUxZxRuuq4slnExTPUStwX2rBQKI+ieJGEXuTYLzr9ylqYt3FHmKL03OVvk27BxX
/7stOfAjDFzpdn72HXnEeUjUIgo821hhZkn2cCWPxPEyph8zqBnI2VCZmIr1jr1i
dEyp18CZHMJVhZYY2jaKHwuzgE5SNpOfzaaigdKHvT7zveEfKTgnVZVO0oy/ueV1
YBvGWEryGjAvKt9O13BIWk2sT4VHe5DZm4lFyyNFD8GKUM+da5L9C0LA12Cnlee7
jfrb4dl1uKtAAxxBLwFIUn7ZdJW4ndOgBS+MV06/KOyEJyPuZ4uCCwBxJg20KvpT
IICnP8p6Svqh3n0e5N3fGYyD/5az8oV6nLfiqe0q0kAoKtHFY+jpNf98c31vcQ3S
YV2/f/HIvBmsKlZHxYFJLS+VgzS1U7zVpzVOpMNCHj4CUiRToMIlci96VrNRNlY3
G4a4DAYR2LIUd1qQ+f2y24B4k1Wzr+WccASmhh0i4gW/wayEAH20GfJpQWwc7eVH
lFtjnw1Ze9Qav+KihWQxidZYfE87+4F7tLJbggyYUbHig7eI4119dKAbZSJGmaGl
dqbPrTiZmhVpLmDtyRgriqiOswoSHlLkWjtpOvgsQ4F2IOjeVqjBvj/uVdVfPQw5
eBBRPq5DjpBxHwALFAnLksGH8WzI0g7PhZV6fza7HVoj3QN2qF2lrHrzHjRT9YoU
X1LTFwa5SC3IfZT8CnVFpKisONAiHEoKgpJR0RsPoDo+F48tqWgmDkYNXp9UKKt7
wt7UHiqZyBulHzchg9MKjYLNT7BEtrqdTUyR6JIKb/n7mkDjD2nzfg5KQwXY4qs3
pYhFmvLEaXGT8vX9kar2Yc07LJbakHSw4XSRuFtR/K1JErj/C8neu4QNGwCZdorY
v77OFXnhWYxD3nigpfNmFkJmdQAKZC99CNlnxnPzr1MEyiT/joPbg9VK8kqwPGJr
IPxIA+EPR7MbDCaczZ5kL4XlmkvQPu0vMBXYgceMyjYfA6PbIr1P3ws8MJq/Nkln
29h40FUxt/m7ABXvfj9cAKrNaTGc9LhFPjmzDyWN97dNj4FLFZc9qqNgZfSrd1IJ
RD7iro4JFaVKnM6WuotfBD9jdWIc3dNmcVhOPKUnYitGSztXq0NDAyLR6vl02Tkw
Ba/dSXDg+uVeAMw9cheCwZY+LEjcY6aQqQU0+ubq9VnwssgaqIXrA4u6R1B0QZrf
shGdbHHFH2ckvVVvLD0DP5Yvd6nA+mnr4d9B3vEbX7lb4AMqO3T0gWPIdrlOjtfh
DQ5kqW5u7PAGwjnaXqfWHSJKXmr8PWLuXRHtrX0kXRLQZpfdayxKahYjSyoWmXMq
UKJJcAVc4rbAVEwL2NHiLY9j7ZjsVsHqqWm//3b8pX9ynW5utJd/5MNizi+XxEHG
E+sY/XfeV+e9GLv0tXK2r/5+JjRxFTFJViLYRxKy5v8m9T5Z7uf+Heoc3qq3bv/K
+3zBAl+0x9PHATrfizLlZs9iBfjnHnHDdTGLkgC7iuOFFfntQNpwaE6xORXF52uj
BZTOtT5+UJ8k0M2wM69F5JWHTuZxl8e3bgLuevEh7D6ykJ/scbjSQjZjkGQlaCIN
6VTkfJUWaI2tcXYIWzdwNFO0ZBbdS6IOrOSXV7X7MoDMDoorT9w+K4jjB3FcfXzJ
GWW4eNwXjYWT2IFgO8JT+9Ix491ZLCKFmk0N4RguDO8aMOB7qhgk5O75R9kio0X9
vGnetAFlg3L2TNG0Tb4AbiqbHN4nmaaduMQg/7em8uKfoJMCPiusNSqMtckhFiu4
ffB9+8DA9cSdrijIygLBx0T3lxJoBzlg/VKlnjwOCcRWHaewAwERmy1QbpTGYcnL
pIFpBmk3nqkUa90e6884PXtKVsEIi1QbG9rHhRy0k7bXSdos8sSwQlntMGuJuMM7
U3CxV4cN2aC3YWWHy9a8gYntNW1ikvn7tR97P1iMcvHSK3ZyuzrAH3pi6dxCcCP8
HEDWYJ+UOYr3aFwXE8gA+o8jxOehJSNbHpdYsK/VDOvSCoCkhg0rDFKZOKdW3OIW
4cr991EiYhP44XnSQDvXnim57ujat222c/0t7jrV9eSJbT7B6IeW08UWZOxMEQK5
7Uf2UGeoTniU0aEjkEud4LJ22Iv/PAL4y6Dix+ThcxjI+yrgFd58R/mpcsMnpqKE
Y2gilpoZKMBpzvI0pk8NYkV1wdK5Fz+tYb4y3EXSHMSyM1GwQmaTltYvHjkVqGv+
/C0JTyi0Gk0FdreRg4IOIrYgVcI8qqHxc++z3AtjtRrF26wdh9kLExqqY4vrIAuw
ctX4dLBaTN9WI339SGnNxzjMaS20BjBAnr9bkMhKvw2vgM5WYVR0QsHlMlIW5+kt
0JrMyT1YVxAmjLsApMkh/sig/h8ZIhTrYiggg/+ObagmhORPETGwgXGKXtwH0BNu
zMUmOeBt+WBDHbG8FoGWev/v6JOf7popKjaNjBASv3Fo/AkCr31GVxYNTVKCQDnQ
3/PJ0Y79NuHQpAmSEgaSaP6sNa3OcXO6NAZkq1V4YJ9Ilv4MYGA8JYESGod97Lou
wbBgEdB2CXP2napnnml5zi2OeXsE3V3rEd7GmVv5zDA3XD7zf0mA6PAHVQJuUMck
+uDU58ckfPxdGTpOjIcm/bKPmGC7RfDaEEwBl9t5l1Kw9TEvLdJqDEOmWOaX77jM
8UtRg3/3owYDNT+DOv1wpHfIH9zbNKa8ct34ZNd49NTYAJI8JkBPb1JfRM2qsdY6
ZTowDrKkUWDRY4zDDofQiqW3it3lIsah0OlHhWsGaBeywxPIeKETNOOhpd1HVfMV
2KwA9gGfe2tR916NKhiCF7cZ2FEhApG5joMa/20trIcZmeacryy2h4BrqY+5UWoW
VQwt/oDi67osHXCze7lZlCqeMOg4shHsej6eIVW60GQU9L83A1Zv5hDiTgfzJ92V
vuIHvXx7xvS074s0leMk8iwwBFkAz1ulHLTXgSNQYCru5/vPzut8ZsAILKdaBGbO
G+07foOoRv6ZgzBXEP2El2iM5oR/5WdMCAPv8U5BrSWGqXnaVFIbvD5h+h5WbjKt
1qOiVkEZvgDmgnfLTklQtzKACr8GQIijiHEVAWDeEpEBZvG9NE7CE057VwN3Hic8
zNmCu68inOXZ9PlnZC3ikPLWHxpl4EZfeew3GHNznfGr9ZhUFbtEZiUOjv5F8R2i
AQthlBsmNvDvLio6snX+oN46D7zvOYb0ZNopgwOPiezllM3TfFlJ4+UFlRG79BGB
QMO/Dx0g1WXf9urb0J2yGDmVIhAcqgk48Zsmu2WZUyVzP9g9k0O+2HYCZfLzCTJM
mZ4ZmiGaF47SE6V92fA4sOoLJJ1p96T+kEsJ+Wb/RZvgC9LEOLQiUtp64NOkX96b
9PIDwYccW6hNiKx8addQU6d6CEdYjGyjGwFaCJn6WQpD6owIOoDWF3DNLGX/VHxp
sxb6AOsGMrGAU7tbDUpYCCieiSChsBFaw89Mp2Yi0zU3ybrqY0lntFFodWu1TGpA
0Wa4sAmuaZh1Lx4YUtCZ/UHUtn3VYTww8m1LgExlx8PjYQ6bt3moR4gUpuOUQlY+
FqWKxWcmpjsBuOHBOb3lBffxfyy7QCYOjdd+2K076FOcf4fp3/W48QvycRtvGcDg
3lrUWWsdVZ1omlIDuXc2v3JD7gm3ub7xEZ+MScQjrGb2RqEMco8txdSeMQheNpaB
XJl4/XR5KVcwaSRJGfRtjvXTX0P98/oGvHylUq0fB2lwHucpI4SNXWK+OIE9lS8Q
LDuUNSkfLWAvYfMUmoskXjisRckEk4rbnFOsDazRJfvfXNzL4Q80E4CEhyNspaJw
EujSVEKlZSqvCtUjp3PS4CYpNKOzw1xqFN6ohGk9H4LG2VMpIs00f7mDDpNUnmfH
HVH7IOSq2Akkju1ch6Nd6Qmt2JIu6C76C8tWpJdyZsGoepLzYFSToKtPnpAlSlCC
epXU6OYXgMLsTi1Qim4Nfiv3EgQVjsGR6xDu3iNJuJXpM7+7jfkxSyJGIvtB7IPG
chOi6iXkX4eE0uPoptd6bAYBPdRmc4v3M0lGiNHp0JhkOV/BAz3f0LckKzLd1MWi
lEVQbcoGz3MPIDYFefWjk2XmiACBsP2rvGPF3dynnzCDVspHMIh1ICfWVicXAeau
1Rzyrrrbqpabuy/nEdoyFnCcr5v4nHQoeFs60rvRKqoQDDGFOCSheaHgiB698dcV
0ElXCPQQvJ6FbC81dR+tNNsNq3DXB93rsEuhWuzeSOw+VMGTU0eAwLNe+TeZgZ0x
aTxc1GEyAOgAoWTzlqln1BBv/a+W9delMG8/cFLW29Y5I7a9T0ImcMiB7h/JOW7R
wl28ABZWCNKm98r7gYJUngpjNeXj9G6o4/mNd2Q42iM5BMDvc5ZTYqale3s7eCzO
3j0EkjSQJnkMg3K7TrVhw4bgV/ojeByTDsOa6J/zDd1Ntnf8lINrzWBVv9j4h7Nb
AgKctMvj4H8j5t3T7Z9vabxjBVaY2YcO0v3MKcKPpubkdgFey93l0JkG+2aJwHk5
pT8EK1FuW+EVg3nC9gqizq+RqSahIWH0MrbYScwoIUJ86bfJhc9aY1mO3oYOJvrs
Zacf1IXMMBWkzr4hro0eQHteXruynbdHCFAhQnaJLMMf7b8Ynh4BEC25Blcsyui2
ZujELNfZqVC1LeFH0XfH9AM0BmGM04fjGeAaGunRjhLufLxoI2WFfSRvrWz/cVt6
IkPW7cF9JYtiWUlKvmGNGE6n769W5rswMu/9cz10q0SiZY9CiNVJ+tm3KkZsfeQo
trWzUEQpmEo3UVY2HP4V157dNJKivaFUv2++c/RRYrsyfv5aVxFFq7Sv12vAx9hE
BSEqSIS2OIwMfz+VDr2c3MRrPVWmuwJOL/g2kGW8IlarDoZHb4EpLO/x0VjyiGkA
Ocp3QSLvILz+tNsSXzDf5jPPG1k6b0QCYld7hEG54rrU3ILFNBMYzBWlj24qESDg
24PoI6wjsWQhB08PBy8iYqSik953AzMZm5ER3V/5L8TVuy9M2af14f0dCGxYxrG4
7qMGp3N6VQJqQSizrk96y47XtbXpNoo7QAe/Sc5ralPMyZa/I28VT/VzTs7gXc3e
mZQcYJwVTWn1NGx2a0GfX63aIDKS01QxFeIfLCWBDGCNlrEMA2U6PL8lB4OXdafN
MpAHq5UJJaCKarKsT8qFANrhYiZccd/77lGvYZ/Ha7zuqR9h067wIvBwWAmUCBla
+pYtz1k5p7aufQRNd2oJlxLDCB9Y+ZdVpr2+UHRaagEOPe04Znh8LMjJ7bwBPave
0IPCrhpBB3P3mCePfmL3B9TAzDcvDhTtyq806AbNUOWtGeIgAomOnP2m/oG2FV5g
5KnxWEOtQ3zAb4GMN09Hn6ejX6mbpiZma3q/u1Rk/Wfhbiwo8ZSabtkd/rKeDRxd
l2cVqc/GWG4vZCjUA8KdIsc2OgsAYnShfPbvidCUXGmuCDYf7lEPmQdNBNeGBtCI
Fg3U9QdgE0KcW64XuHqe8/kftm8BOFjaxaoi0BwOPbAJiu3vHu94f7RhfE7lWf4Y
rTVGTQ/mR5f0+eWi5n7SKidXa/uCaqcXdd1s/uQFhw2wdOvUecgbud5t76ndmYNH
BFkHql6RFhxQqKxsYh9RlGgNdriI46hLXBHfIpHuI9duB5UYaqexxhIxAQP8HS1G
mJGct6stN3a2zmsQW/n5OrzKSh7zvImpCmQe7zLC4o+gFuEtjN2AkZKrqE4aHcMY
7beRwQSjTYykLh9O6CRotft7TOZkEAoM7AzBikLlPFPvlIR0ECS4TxxfSOhxnXqz
ZTJ2r94zqpKFA4bWp4SPCD7g6MvJqNUOx0zuzSH6mtybhyJIyf7OMon5xSi/7fRC
KQ0bCTwSGl0a1Ar1dJdns+o6qUvy/N4GlgqmYfL9kYqVbn3fknFETkQBtQMmCzZC
EtbkXkfRRH89GVE9ADLf+8V9y09XKT/H9/MW0H9unlDYvPTr+q0irVZtT7D5w1FW
RnwikLGFABLG2j6VR/UDEVICsJ5IrPI5Xj7TPYSog6SUUacDappizpQsO0HfYb5t
JFnAD4E4FIIjCfvlGQt0ArLYBPQVm7aZVwF8A9tFTlFSp2k2XNDQKZGra454zorg
1dHqqfoVbv+fxphhHCGmsNySO0kzFU7oAe326Ib8jK8sCzUFW2oIy/uR15uaCweX
Zj6LI3oBfoeSUHIJj9Wc0Sz5Is8IJErqkgNFrhcGy6NyMs28oPbZMD/L7UG4Tq+u
2/jUJKagaz8gv7339DjYOpbZfUAyZqfcI4q6tg+cuiJmRrT4daD9H9umWMQdQVMw
pyD9gWQpJFokz9FZvq4dfCjTItCM6nbkrWQM88QPhvxVnNzC4auzeVsVb9dxWVHG
ZOhmCYwdwHvfooNHpk9fsH123brBNuGNAeMecpVP6uVxSlaSylC/spyv7iJYAWFe
AX2CI1zvSX7fUck/I19UOw9HfxyjUot1sflQIIj8OMkIpHUNRh17xMC0fIkRz0jC
2aewrAcsHgggL3ZrEDQLTQ6GkaZKHDJ8EtyvMIA6oY6iE5U2ZUSIaffw1TZ3aU7B
R3ozLnTRXRKTtc6827pf3mh32776vBJwJK6+Hn8aWk1A/IORUhzEHAAITqYa/hdU
5HwzLmd9Rm4xj5sIgsN8LK3HPzK6Ir7wLQiUDsjjaasaDk/HpjO1gWoFrBUWjmdG
GNljF1u99N1D3PRQDgK35ohlFp/ui53lFu9lOFk5y1ZOltEusXaWGbLivLVpti8G
SEiN/lbDCpEHorOKKaG2CgvsIdQzCiXvW2LHcyNi65TU6swltxxe17xa/vQjiUpM
OYya/3vKpiAmRewmS/8MnBHTKtCdtx3pYtjMl4UYQTWEDSRi1JE4prFctOFLy6/L
Qz6+NEDvC0v8iRk956sZvC7/pOZJmKZyiflRwVbjCTRYxlkqgHABiiSTcwKVeUQh
9O2i41igbXsFSk6vPcHnot/UpdJuJ0Gts4S7wyLAt07Oqm5tJUj/XzHBtifW7KEu
7z7i2UjUNHKmhh+3RUIsBBtO2WWNleOyW0Vs4QbIRT4ryTjthC9CvEglJqUsDaLM
SdBO7JM4XaYC+sHoaOzrvluYpShQ7jgXOOSwXBsghvo9i2cSKX7GKyx234M4zxDp
lK81LEszWFmFmtXaXnWqaY0abjFXPAet/kvO+AZU0h6x1CCNyZAnM3nHqPvM+CZU
BSv0RsCxbgb93WGxkTggXtji1Qo4Ic195yLqVApGvZAWe9cmppgiH1FYxyTFgLmq
3fLamaBLKBWwr7MmCva/pzo/fSj9sCy4Rf9829hxDJsQQ/WyDOTWm9ogp00Kb6mT
iTiotmBUkZjsh+brAw/CBIH0vSCoJ551YE71EfU2mF1nuk/0JM54n3uS2/V0NKjJ
u8qi8T2BQdNMI45/dfHLT6QK1NJhskaa7DPc/xIk3dPa3qLJjtxfRis5LQCn21bi
34lnDivSYBSEK6oaKBUcl2ctq4Ux5JQXqUAfZYAePRzNpXHQOk37NBxXVf77hZu3
ZyYNCCZwvGENIuQ44p91lPRT1qAqUxkhg+ivScA8yuMI4sFjuDIXS8spjYKjl1c3
O4LUOfrS06riUwJjKSQPhotnpZ6KEs1+kq1FZr0t7BQfpU3m+0hVgyrCGXdX0s5L
6wX3PWF69gilT0FEinRKHqN7t2ATbz1+Z5oCSh7dhltaq+bR4lR6ixHIuy4zmPY4
o7fllRTmPI1J7OXzXt+uQXF+oSO4PpSkNimZ6lkmoR1S0Vxuhatgxk9Lw+hFi9rR
GGpLegKrfw0arwuWSS7zGOpVjKLPjVhLBMtTsaJPes22+FkLsEBBlASNXwibCYF5
3lEnkqvE844lhCRuVcUcmYpBC2vrnV0c5NBrHr/n2cxPcsPr17k63IdFEjp3NW1C
SB/OodRRZGxuWvxmfseaEJasD0E3KXyLXfLi+qxrsXDytAsxfrJfyW1T4ucUdJKf
H8dRxSXJ0MCRqWvaxRm+BqvS6IQhl/DejmmhhMFJdnkqw8CSEXliJEUP4ozmYeG0
TQxJj4ug4+Q6ZtAkgxRnqYwfUrqNYJNAg0mgr7YlD3dAnp9zVXl2MGSUJfn6bUPh
dgGS7JBPH1BOO1SVB/Qpyn0XP5Mjvhco8PBLcvsyZC11lSC1DjwE00GdfL2viKvv
LxW665zQ/ecdaSS+u+8yPVNxRlgZOlBO8Sk54ZgqfsbV3bkKDIaxJL0fR8URDkXB
O3cRAr0nOnQSurskYOisxUiOY+hp7O+NfyB7XaJy18PMelJGC3A7SA7Au+Hr0AAO
Og96kUR5pdW7FquCeBznGDwP/xlQ8fzUhdWXSvLDK1AoO2i56TAQziZhLEOhSpxI
NMjDAHIyppCbcfI3rMrIODuIGFMyNWnZOdiaswzNKjS12Cw5PuS1gLF8JXwNoZTR
0oflE85/3G7ah1xcQY8/lWMSX4Xz0BfRvfxkg2j8q4C0GAw1sz8gaD+36/Lx3KzO
9APLagh0bUr1mwbFNpJLKpt2+N+EcLvqVvfm3oVWbBqIpz/ZVub80ImOcNiuIaHq
yxhhXFS1WqCpw1/tk6D1So8XyUX50SYMyAjB04u5O2+SOQNXrh3KSGs7/fq0BVV2
iIe4XxyHyawM0Lhro7EMcYJcx//69qNRaDXQ8TrSp6epuRCAfg65plUKnNMnasQR
r9a71NcvN8C7pjMItRr20GvnFl84jYhjxzasIEHY0bR4WTiDfpzL2kkQLGmISF6f
dRNRYDMQSqCChVHnLZ/Jsr4NSXwNcwszqSV+nRVa6j20HmVGNS9xar+u//d0IpRc
CeXRlpHi3mlM+1ZODNglJ+dL+oSO6h6Ks2yxMn5Djd3/hFgrn3aa83BMpjW0VJLo
bIVeX4XANreMmDrX8+ELLnC9s8maoNDuyxzUKUJxS5xEZaFccNgRA0Rc/v26X8hw
FKUslMUKwyV3MgM3lCrlevb3P0kI32NtdJ4S50WIzS/l1VhhNjMzzpHds/GT6Ri2
4t5lRxybTD47o96CaGvGHag67EHgh/5o8M7X+8+RW9Cx4flusokpDw8l3dQEl+2X
IFHCDmUkh2w6yOhMbczNTaDUhSNh7ZfKh6qOpnhiOzgCJyrZw37jHnZtC+E8WfOt
H9boQbJSrPINAnYegF3pNHVn34OXe+/pcNaSi12z+jL5V/npZZqouIcMi3/UFdoY
V75QHKsThJXuCMbVItRcqOfq/uDXPAjLPuo5HGFGekhnIck3GSxN28Ad/1dRXOH9
XcbtObwRG0ARuGl9i9ssqP+iK5FcMiIz+PNd6MW8WAfhfL3s8fDL/U/tVZHkWTrU
sZebDKbxvt97L9rupoFLVnrl670yDKXmH7Z+/WjpSBVtFXS8jXfpy+bbgFmwmsnX
H0ERPiudWcqe4jlP86GVVw4SZODP8CG4F4svof5sjh80RuaLW+SLj3D8yQSFBPvt
s+Or93WwteHKcoN/7pBpJFv9usLL7OEa8ip2xlzzF41+eKJ8NoRkX1GWHPzdDIAC
HxvDwtj3Frtdr1WkotEn/A5rlpdsLclbqPQ3XqPJPL+UkNkYflBS9nZ1BZvOrDW8
V3YhES3imagWsvNT6tOgGAZmWdjK2yBBVjAfCEHplCXf0brEL/2QzYrO+W75N6VF
0ooseq9wz1tSlG3nVI5yzsolFWXcgLVDJy462Ig9pRinZ+i9OXnYxVWprz5gohPB
h2SXdeKP/C3ZNvf6Gr0CxnzWJOLehsxUYWdp/3SoWzUhaWUYthBqxeehMcLfz2FU
SYt3k56jSlZw3RmPgIsCFU9gaLY+ONl2HnpFZ4lB6Hnf+JfvGXC1pSvkSHe9EN/B
1pQvnwQQ73d0/jJCSWc9EhmdEFtldFMEK+IJ4cT+4FX3sku0lUWoPz7z75le1jJ9
pqtVigoBADiYWhMNl2wzzztSo8+s3hm5Lx3hRMR6IFWAleMONKP5exOgPyIFU5dx
lO3pjwovtl6LH9dQtTBKpaB3xt6kfwWiAjM3tzijUskrXS/3Z2YTObmmW38qqvLz
RkzQke5pml3ofAKNh8Tb87zxB6kIfpG6fXYFZbCc+rIInV9jhJbnBsyCvMfxcva6
87//O1dBfxCC3sg68Ccov/l4GWXVd9F0hQ6WW+yXB2hxvu29zdxlJoEHUhmo5cOU
pAyhVifc3jwpP0S4ZR/NRfdAKg/rpvyq6jNUWDRmE8Rxca2VzrdFVyhRc/dQFtkH
sw2i4WCi59JH2ryD5V94JuT9RVt1Xej2L8ZUCSs1zHOcfMEW28sLi4+jme/HKcYU
5z8Ok9yww/SE5w5eiZ8tt/xpM+YOF6G0wpRSG53u4ktMc6qNONmiIJk3gPzlB6lZ
KY/o9iRDfbEg4+DeAZtwCUJBMLw7S8d2qFMiyyLQGpg6g47yJnMKnrBJw/6LTLC5
Iqg/gOwgiRqBt/IQyar2JZ4VuMgGfD8axyhqLr12vhVNj8WMYE5SyPDwpthL/mxY
zK38yv3zbSwEzKN5ifg+fCiHvFs1m3gVvaVDsYeE7WaJl4vXh0qcGN9RYry1oI94
OVNwvuFUpNCCPE+PbaubSDK6k+3gB11wGAsWf94nJUBBQHJdIhNbU/YiTn69v0R3
dMHeM4+9wEqqcH2eNiJ5J48icNIVXDCINCCFeQqefHMrIyaFXfkjrQuGlamH3uZE
ex3iIb/WBNLI8nvW1+UzhUrJZzcsPOUro0iosebtmaAbVKNnxP5xd3/ZMEN5u7Bh
URuESXL30O1Ylead/4No5PMkoosdtH27l5O2xH46e3D8Trz8+oRGzz9PheSWVlYu
4yPl1XinoaaYEIf6cZ7rS2aWL9LmOWnl4WUYJFlpI3sCu2+ckFiW8xlXecc6XNQA
o9ZTWx4L08kkRXc7HvuNTjdM8+WiGy5Z9XGFkbDLc2i97GNGo/RNiNxkww5Rvt56
KLtNWwHt2za0hATuqw3LFiIXCqsVApcJ+6/tXJOLNAgWZ+tvWOaHK70UacYUPobv
SrhAidkYR1utQauuRjXzvfKP2bvTu1zGTYyvHsoggcV4WfYvqcFrdkj2p4eXoPgv
e5QKTgi0NjaKJthKq0DRCFc5zRSaL1eRo42AubtPzTUUQqKqKYepfHapuxT2CL/Z
p9LQIrQA6ulyvmcfkPjOC43AIuJ3hC9vxzqKihMOCkiKyI3Nfc5GBRd16ASbmFEo
rmSYqsBxcI1nAOEXDgiFU/18sGDIRkP2ajjY7Nm3fqvZeLr1vbmA2z+vAp5ZsfCL
/J1Ix0Qis0BQ1y8GK6f0YUFQhFLcA4WlEyTeSHo25ueq7rX5Ny23TV+Ua6yfXvH9
x0QQPAhHgDrCJd2h60Tc57dfnW8pXkCsijg6weWepsyrA3nRncbeQlvtDLdLI8W/
0imO4JlLhzkgjHDv9Dvcu2pAN/ilPVARj+4ADGZf9bh2NHT78H2gTofxryCXnj5P
hGrCeVGxgTgcLDaHu2TV/V/FqJnYV9pF4ch7H+GS/XOSHDu3yJYD5LCQzlL6Uz5y
jyAttGN8RNDzoOC7luYIFFZeOF4/JYAsIFdDVRo+UldR9N8I6d2jgiV799N4aa2W
1kc5u2/+J9SWLoIyT12n8Cyn+05/73mqrxWPGyJYph3kpvpz487PLzG63BZvsJLB
dDHnFRgQTvIhZy7vHcG4mZwXDNY5y2PhwtFCihXnXr/rKGVO1zmsSIeHyya98Z3Q
peiL/wVrwDlh1jmFn7SvhXOpinBT2RGvt6sMSKgWzvjcCXVVsEKetAdUVHSmK3e1
Ea0wVk0wPxmFYz40BsVtyeLcAGKb40p2eiYP3WYj4FTpeiXwEnjb2q1xAlCDBmDR
oXogz5bN07/rLgMSBhZaEQZ+FzQQOatv6Wy5hS/zdDeESdZojv64hbM94EJmBhPf
utdHXwu6JHcVE+1bO9udk2+KjsdAsC5gNEWkrqNB4GfHWrnfyGXigAvT4v4o5L5/
S+zt6bNFMXNiYL/8Oz7EGYnGRk7nuaSpkT0D0pM2zruDY00NwatAAz8YN/z+WC6h
Lj4MWwgnKcKmZOGGw5uEtRSG02LAFFyiMMaHwAUrJhrqC2DQj8fp2yV/E25BLg8I
SKyreRNofmMAngq4N/0Jmm7fNhQhqBpufxGNjTUa6CzDnsrg5ApGae8/Slv0FSlt
LXr1ozTH/RUMkCVE3E3zfvV6JpBnXA6RicyugaLIUQym0beZRhITZsnRgK0/uYiS
B2AR78ds5eWPW9YgVst4HKI0xiM2gP4L5B6T9DCRyicBT/Z5FX68LXvkj2COMXAN
Zk8pEqOcwnDh8v1av9OM4Df5MCDnEUyg46PQ3YJVJ5QOyVnIakKworAsTbR77mIx
tqcO7PtFQqUSRh1a5HxoE7G+Qhq5lS0OedGJp3vihTIkQgMVuFbZH2DnJYUXuozT
1rZIKlvG6he0QhjvuvMxZwenQLwVwxHcqsEwv3GY/Gp6UvK0YIEZ7OCHNDX5hDcb
eXL/uyZ4CmjcDpwve1gKptlzalHyEwaJE6Tv+I3G+HRzs/qhhrB/7q+WpkySZcPr
H/8+yJIZy1ica/mVAb8MvwVMo1W+KmW9pyz2CMtFnvAueXqQmDaFO+V912rlTuLV
i8996Fgb2QL3KkcJsYToK5y9K9y9SChont2mmswR1G5Kt4j58O8DJv90ETgc96IN
1VqDGQ1zx6BGNftW1vnlu2STA+hNuSNEeZQWMT1iw71ZQYZH1OcIGooQeRy3jQAd
GQbbZMyJOHfgU0mapcbWxRPGYEfqPCZGFDjWwwLysrfQBgPOq5xCiCwvuAZuzY9D
0/MP8JqWabgQVW89bzRSdT6TYu5O4lK+h+HJ/B8DCj3htF+e+CqxAfhHNn5/ky1l
7qEWymkJ5wcKX/7H7B6Gx0iwAPbERC7XJEIaFuIhK3tTtGXKH8QZBXGhD3L9oPJV
861CfLjdSTmApspXw4nL1ADsHsG8KFHKSFdJ4vxj/OX3ifbz+X/00lpJ8bS9FEn8
zKABb4r+8/QCYxE4qmtL9/IMK68bE59ZiHGqVZG0TXhrHRAbgt6K7sEfSPARBB4R
28/9IYMUZpiC8juAJ4w6edFDrTcnco8ZEwBEWtvqBsWKw+T1y1yIJJVXZw7vdO2x
zOpODAzKKEHSzQSF5LJ7FdmcWR9nDXzVf56RhGGMkRvQwGihHJnwvghNZRFehm2z
v/mQHdm5fTtzCDfRHm+lA5hknG0NeqvPzX23qAAebYBqn8baKfslOYE/TDE5w8Jm
IZdsQMcNsioC1Y4Aug0lDkT7YcXDie5ihbiiMQnArsyQsI2wSi+HyWdZp7TwSk0V
7FH835wVtlidUisXuw4KX8NcvXNKOmz/sICSR2Ml0o3cXla3Aw17eJ48PJuFi9kU
0A91sNKRNkR2wjHdGDLjJup5m4fZ3n4C8a3sb6jqTEde1E6Bls85/IAzIvpFiFcC
YDlDPhDZhvIOCRd4a2thZ2C3p1tydpTTf6beDjOs5MJ3EmPAlVrDg95p/yXkrPpF
andBah+nhI8ixE5KKT6g5f7NKWd8bPLQpcyDStWGz4zMoOTU1sKXUvoy+uGYuc1z
Oy66E1K0+fKNvKuoo3O81Gy2wZZAwiKnLYeRPiP1LG8Y3jbp9gkRbaByFo0zr+pu
TZOSUoV2aX3NIccYjK0wNKs6O+UBuhNaCBLCSaG5sTZZIVuC/l0TTyw5FLiGfjGJ
kH94IUZDb9kuBJG3EibtHqLGMHh41FxbFYyCoB7mR3zf9eho7+uwfLIXyKSWMYiH
pL/S5BhVBt0S68ZtN/rkP8pVAgMiS7YeakSFiVJj38AGekrWxf6oKeV+D5HxK7Y2
2FsEDWdoVAfOhhBlcput9oKyb6P5qLBBMwoJylTqDjLvK/PVRGEUoBeQfPPW7/WI
BVODZ55iUbmPkMYc6dREpG9csZqSkvSJ5V+4Vnk978ZmpqyaYYJ5EGaVUHq5B7N0
71l6bVoWtTE3BeKkhu2/68V8m/0LNyi3VPYXkOcMPJr3UkAKk2s+zVW/pbUsPoeP
2dgJAB4vgOWkLX+uww28+kBphJp58pEaHnUnAz0rgK45JercIuYGmZZpAFuLjC6L
vRMdoy0yaogvkoDB1Auz/CQNlxaZLoR2AdU4yQy4AaDv32jRr4hlL3JRgzXQLOVE
8wKa8W+63xLytbVeuT7wZqR6K7ykPQ1sg5L1xqKljNkg2misZEudTUyw5UyOyJ+N
/qlmcgDeDM7ca1LrxhpwRBP5PU9woAuTaoDYTEezUYVz4OErWITYiPROFBuv8nIQ
vwYWONimjrLtvzoouLSdFxASFtFZOMO4ZYSHG/3et/CR+/QIfDO6zWVdOV8t8t1U
zj3CDZY+kOsTJdh4XwE0bsk7+B/lNH5mS3e9GSlEA4/D2zgu6X6gTPqnOVushD43
rn3i6cMopGsCiAKgwGLXVrjmrLqCPYSP/vWzD2UCEbRHGredacaelTE2k/gk6dKS
MiqJH9S8J/nDJ1sRosJZZPXFAJwq53CY4I9pifPZCt4BwhQxPhyZ/jvG1w3rlR9E
FtXa2a4YRcu6NmX2U0jcppeqjtQAQhPp8nHkQaWPZ2mPDqCznCSbvx9oxB/gc9vP
6gVnCLkpOt/puv2kBYrvhCZGv7BZJG5oMy8ct9PsBZKQei9J9bPs8P1hfyOtTxn8
wwePbwMiTU/ayypnXYCM648qasbVkvSxeW8cfInM2QmjLN9lUXiNsqcNRibPiE6P
jnAfsRUv38i6Klx1pXGlTZdJH2QwzDdmnRFb2T1JQvt9IQg9x25btPuO4zzplBhN
G1BPaARNklUiXT3wmrZWxkiKdjbOcK9zHjBS58/fmFiSPQvTcINhUaSKtCCJncw9
NeSd9dOfDBjVH6KjETAV012wBX522Fw49o7ZpOlOsl9yaMlgFlmvbdPbMpsAna3S
58+6sxQY+U2kWfswA1JOhgD/h0XCAWT7npYHKb7jy3DMWM18F89hnVMnYm4L2FbK
MFCx6W1AMCZnXGBy8zC4datp0fVzVcTSVam8IzuXZHTlKOBjSPQyn96aCcGqEYS9
hof4oXaKeg6RPCHci1YLdzstNICEXbXMw/AcQrKzaJj0bAaON7MsbYmAaJ6O8EyJ
TmASfKscsLr3bvVCnacqBb+oKBevUsAXLU7AZRV7bCwu83WWEsL3N31XUZ452CnC
5Pk2bbOuGNHLAelDD9V+mYmoNfm9Ctu8/hl7P+mQ9ZYf0ZW2VEKhb9WD47nwTTYT
SS86CMXoR7CtpFCVg+AGpZ3g8Pv6UOHZ+tjBzfSrOzD5LR8h461zw1Ste1ZYfvQ3
8zQMbf/frToD1BsstWz0WcZfzTxmXvvR2z6+0/q5gxdKSe/jMn4c9ATMKQXFt18E
4eDhNUWY0ssth8JdUL0iRm5rPRfKFppzYgZ52iNJZN7q9wY7b0XIgrr7rIGCJf3y
s1zA/Y5hgRw/51s3pDr32lklkndZenL01iF9E/pfgI7DPBkbK03zyJ/BkRZUXZRS
tzGzD6UHQ7mrsyjIe+coBMa6o0hhDgzowYyeklnynF9orsWlUj84yx6DCxMgxIVB
LbrnTtnPYtQ5pUbZd0mZMQGEKfEfRqxm9Asxd0yGR/ncFYDIIA6fmRHM6LDoVyBX
NTItNQKdtZrlDmFhWkIXUElHh/nVKPiLZz1Yo4lKS1z4xYj0/mtwXxPZSmaKHkrz
gwBvf+vPuo7ptjKR+IPfaq9ZXaBPbU+A6WWIZ9Zq+Egg939G7uM+pg2iC1Qn5LeE
kWtoOEnA2+RO3mTlmi2sRH65APnsmvUEhCsJGZhFR5+oJM2Bm5DO8PGeVxioBxIK
WaEcDUytbsTsAZwNgkjXt9Mvye+VcaIehcwTNWyN8yw3kCH/3nKAU/m++Qt/kt+I
zjGl/Zc59LZh257uvFbEOuSg5G7sAWQek6VWrwIhNectZq0nQCgqNa8cRrbBDRm2
uhCp+FdG7fB2TViAn18xF9J0dGi5PcKXLePzVvhQUUu7EtsWr0r8lD0AM1BXvnZS
xSzkoUH//YJ7VRkr8X8+X1kU+h15lpGUzELYVHmzpderrHI3Vnytb+M+4sur7chG
GdkPH8w52y5C/njn7wo1CM9hBqKN885+Sxzd5ohH1yxPeOgB6JN92MlerIoJwPVk
X9pO8XEKzYVueL6uqj4Kus5jva96UoEVBqUVyDnlbqEvsCaA5aVpdBHdQyY9D4Ay
VoG03fyyob3gysN7JEjQpRSExaODZlSq9N7dwUGvnNEfZG56KhTfSfhQ3EGVeHf+
95FV82mK0hUliJalcS/laU4dEOAonNJ/O9/QEEbWYSg1kfFh+vBEhS5nsB0boGbl
0PwEtg/jXWyWSFpey42NSJK7tzLq7s11DHMpOibvuzsKdSsZQ2nLE0vbYU2QNG8T
N/hlzB8NhtZm+yipYH81aqHPPpIItocIXvHukdIkvYdv2jxq0M2vocm7jwpMQNl3
49OvSMOmRmUZCfE9hhXOQQbrOnvLLqYs8UW8Y5x+6IbNhYB8FCH5ICZ3h8rHbIH1
nzjngf1i+K5Ctgx5NahFd1dTjhkn6OGE6tZHqvBnCGPCctIHV553RLi9jxaek9sl
kcNdLaAl/lsxN5j6CsPD6mymIej6sGdTxGPlLIOcNtGJ1DyEFEViqlnJq+WlT418
2tIqIKvMAIu6ZRhfScXzuX5U8+qz2sW9C0cHhhfaWeUAcYCYR/P+wwtHi52QK4qe
K43Xn1IL4bCYKe+cgMxUBDQeGxeZADkHIBchKWowmGPUVRH/rqcWKXwoNNonPbFw
MYSuuoxg/ZHm0NwVEJuRXw8FpjWXzmBqkjpv5qPvHVBIA7RFbkZfdMXorqiigI9q
itHi5R3879cfouXgfzzBQ6VgzDt+k9qIhxCmDoDmACPK7AubAgX1VP8jkfhs6Zw+
1uWgnB8GrJgCcXykfA+wHdPqKyMN3nYTaF9TLyCTv2h/aijJA98rsD5FKpXjBINC
3xtzV7fpBhSVMXJgYHPblyLixwaAf4XOgHPnDpUwR9DB32d0TbJNQMap2qwp3tmG
cpCIF6rc3XZ4Tvwin3MbkJKs/Y+4nwavp8VN7hknybSfJSuuLrm3HJ3wiew2wEja
wMWgjF7gWC9t35rb0Uh/0sBTHXi5Y+nOnBM9YdGOSgV1H0hEACCpziF43xm0uyKs
ggw2AdDjccoE0qLRHRpP3c5O9+dhn5wm0+lLnQ0S59YpaNgZHXvRYtwwK7XLn89P
MTm/EwBCn13zPTv3BTN4m2hsmYENURi4ZPMhNZri+L61oS3lur7p1eymq4hjJS7l
sL8++x63GGoPRt+yiDR+FRunRhFlLsPWVfSlD4yKSl7kZH5oYMqaTQssaft5/dy8
g6zgz06H/B9daqHrYii9KCP2blI2spCEvSbYw473zWbgco9GXNLKVxNNujVSpKXo
xUhe+Fa0Ha3Vy3Tos7JCEaAvHyvA1Vgu+BcT1WzQG5Sqq/sdNqcr8fc6RF40YWqH
a880SJ8CZM4yAxYsl6rAvCLizamRZB7ce70q2hVUkfOtRV+vwnMLPWMeYgWkiSxv
kvBVS+RVnv5rffNa/b3bRGljQDfS3JbnNJNSzuP9DoKOpcxhMfXbjXNsYCRFBP1y
CR6sJEIMIh6w8kHYXf3coTZTkBy/yfQfWyUfeDEQhgKK8rfdbPYduGHHRrugnbrD
PylUjguivjjUO8ikwXjHnlwFc6eP2rs/Ah9msKKYoIxXFhhUjrvRcQFFHrySd58d
srvCNhM8J6XL0ZIZsegK02j+Ou2XsE/eua2GKLPRVnejUKgv2aq1q6ACWgvQ9fol
KeQ9w7iFZvGxfQGuKsbfBrVNHjhXL+DNYNegvTCCLZsNLy7rf44kpkcz9KuDf17N
bRyT9fHBnf2pqejODNfti+RoV2aCnxB3Kr/Hu24adGIa/LdJezbL3RRPLLgqJsYr
2ZWHs1JEwamDOmLSVB+9TL7Kva6ZAH+ttAioGYOdkDWdnmTPExy5l1dnaWh6uLR5
7eMQ/JE0fd8pXB7RLdTZ4nxQ4cm8+MgbMsIRL8BXQikXb9aTjGLoa/0pbk3vDqZD
MisTXUSfe3NYkREF8XcDgMiK+x/rWgFRi0ErpcUaJLvtof2iLtD3A0S3A48/j505
8PT4ATxL64NfhpOJDRTxxN72yqXQcf3mmXh4SGuer7vB7OroEmpBGq1wUYVsNIA1
uTK5uNN3vRVw8oP7/HZvMixyEIRLIjcURexNdyw72GCzB/uYzZo3s8Q4DnB97UNb
gVeAQ4M2qy4/OPHihkY1/MzTqNuvZGgjTUNQU1bPORHzAfd510FRq9i0WLEl2McV
W8LgXWTw3kTgi4VFufwgpdIQ/YT/ssl0gkYPdAVIpmFMfGRpE6cFW+QxZDkYyAa+
OPpeh9M9D95/Zml73xfsYNxwxrUI4EoUJfSi2oUZwUOHEtQqDwF8xZGd42/9l/DA
8vuUhq4zXY27zpQePNQF/X1494VEfeHROb8B9zeawJ4qbKiwibUkTC9weumD3Aoj
8HalF6MntbdQr4zMNp7+IPqpaG/tqpLPftc7uMQ5OyF3fO3AqdEQXquuaqQairKn
d4QY+2y14u5ybU5Q5GaaIxHdJgwOej2wprfpyDoDhloGQgCsHlM9WU3cyaeBarxt
TYsOKxEK58o0mysk10Mp/w6EOUL7ZvVzb413lB/123Ma4+jhDbh01YwcZjQXOpyk
zJmNgsjqLto1igOqBzV/VnWFBEN3MbBI7Tp+tSOV7KnxtKug2o/3MXcJNICPjIA4
WEak/bIGvDM1e7LKa7Fn12xNqHXX4O+g0mC6jCrBECckJH7dIEL1HJKvi2dPXX9n
H3oKJr7wiL7hMPQJkYKC+/R+uFYHwFC6LzKatyAgjHVX2vU4WXQBiJAIRYad99ZW
VqJJsRBxWFUthGURLBXdpj6hwhJ7KCdl/1ns/JsbulYZDmUEY9+rECD3SDrVt20c
X4Inx4cDGFm5zsbxXYusFL5WuuMbhrJ94BqV3ToliUCaefcTEYeaOwoGc+zR/Bhq
RdVxFtOgWt4j+qkR4NLkAvPZgnowHNbLhxmVl+yJS3mVvW2C9FOqJgDSIMvPEjwM
ROnCpJlfKilZKa39xr3a+VuxTJBz4POUUdPGMCZX97sJVzLZt3CEhW7h6SCnipBr
+OTQiImsspNrLfKUfY/k3Os2eMxdlgFuOv+DXvMhFPLjNV5upStZ1ABMfOY3tdI+
tEHL+QVxkg0+zJuuDE+laC7o6QnEjUUh2dLOMH7b0TnDbBrAPeJGcRa6zBJKDA77
aGUVoaD76U8Aw1sFUcSh+IARXcuizXGlhzImC6Tp6A2MZWU/0g1T9BoWcxywRos4
hHq5BoHDlL36o85uSsy9fwfzZEZj/M/7jpmVU3/U2+1I5/HfGUXcRROj2xalUjUK
efvigl2tjpmzlDCsRpY0j4xx2Xgv1Bluo3cvDrHA1B2jLvMldOMDvxepXcm0yG81
zMttGTWLA2jp7f4aJnMTgyjZBqqanV4TyFmnZ2XhX/IZ1fWYKPihCUMJGe0xn9pA
3JMuud62+YExbxrHwGaOYHgcYTSW/j43WsJICXPIMSgIQKap59zvRftxQNCOVso3
aWeBAn1FiiLax5z9hBAirZtlZmEqwONJw56nFuedKIWkTas3rvD9mNEKF7paJbff
fpoyqgFMK/4e9lgqTJNbBltblN2eORW5j08TwmEZAVGGV5JjTwZqi/wS+NHPKi+e
YSTf9/iXvmlA3BhCy8eZDjvs0quga9EmTs2LEnqtYEoKhIEJezJD0oym1HJL2d5K
HY60my8hFyqTcI4RhWU/MsKQxximmIzyDcyXIma3iWsNr264vIR5JB21dmzzI+AG
0C4N/xuk0g6i8on+crWr0KAwjaZ++Ut1cKYyImSlvUQ3e4RLtd2fz1sBoi47PqJe
t6IAES+WYmoh0876yrarSYoeNCLjcLRtbzoCRPoC6D0/8TdN7u1WB/nC94EnxZWL
jkQ6T2+AXtewzFmyqxTMDCEvgb/u0qxtJ7OdtTeu/0UVB/t8U0puQ5nyITc+eI+Z
xeNTvVU8XBxknqNfN8oH6k5w3s3oRwWOkyUIdMR+6XXtyy1rDCIQ9n2XNBq45fJK
C8csKsm9Vb9rhrLdZC4XOwlFtBy+X1kjZqOTwd+9wqwkmMA5xp2oBCOwXFNjyO3e
UGjPRdGw6imfo6x1YUqhUxJ2BMSGpUITj9EU0QAjdbUG13I0ar8ED6pyFgdU0Aor
lOnadzB8jTAEwWvSrBUVVsPD/9oDGGWOUsAz/T06R3EuTY6r9frk067FBCYTBLkk
xuuhFxbv82iC6P6Soul8kuReQWwbRiPeQQeADGl1tL9a8bC944ZlxgfAMs0RhqBr
VqgXXqBbheyDOwNNbV3/gmnB44XtJC4KVONwc4McoQTSIlYrBttP3zLWVz7uataP
5UQmp7EHTuCY5dK01skADHzNV4mOMwvDDFOX3zxy0Dir8oVVsz+b7ahPDw6ohB0+
CD9NiSBJxNhZa9fU4gosD1yAsUWzTKqrFtvAV/KO0Z2fCL9Vl77Cgv/zXtdkMw49
mA9ece9V47eccyQbypB043/AGofNJZ0ujWoMRT2aSre5FSeJ2UQSszyLqiEpV6c7
Ou6krJHkqPn/4LoBjGLPAqqm4loDBpwecqhsHuhuF6yQ7pfagyFP+qJMW+Cjkhp4
QQ0QcSa2iuvsBsNQMcncx7AKrEvP7jVOR3K98JcbcQ+PZm1oJ3idD4HqlMRV+7Df
spX0yhlEZG4GKl3Bhmi7XDGIDCdwbb96CVHQQtggZlDy0BbDzhQQeUZUDU0lPLK4
izddallbVuvts1F+NpdrbiPf81AFcbzSdVum2jogYx/ZDk0Ze0S6FbpssKeqFZ1l
os3TJpvkAF4XovkwwYR0T2+jhrY7+oMT2TPTHF8qDaRrSbpSVSo+JNAKdWCRux/7
+kZhlEO/CSH3EA+ABzMHxbx0AM7N+F0lHy1gq5bcKxYtlXo4weGZ0jtDr/btENNR
zWVPxfiTaPu47rX3yuIezlZMfFPA0/o6Rjzx+ebInmkOqwwwgvxOf8zgv9u3Diq/
cmm/bgpuEruw3/NYLgd3xCTXw4AiNAbH7FlNlOrQVogz4TeSaDQYXS2dkctdbBz7
UUIdfXolFbG+1FXszCQnpj6Kpypx5xR3H0bab9pHcR+SG1moysyArXNxbEtOmhIi
5tUfAxZWnVU6S2mDwN0pT474067PdDT+zKp98uwOvttcAcGA9I5Orm5g2l1Inl7d
gOuMdFcczfkPdzPAQC8spSmgDqRwM0dQTaHhMuHpR0U9a9wvUBf14tOI1trXvLxp
f6O4+4Q8z0dENnqh1+s8qBzetB9+hAxOF6mSk4evDVTYi2AhZVxzrCssAeqA69j2
ZxVIjFZPJ4aaqMi15tQCMZAnuEx8+J3+yoOeYfXYjeMn8RrtlRh6mZNR+9QPkxGu
Os7kslDTmgYxoTen9YOekn69JNDpYwR/kL7z2bz3GIkL5DaZfP9ZZ8jHZ9ms7BEx
b5WR+H8hXT25EuWOs/M34T3vzZnx+cQc0PGWEkeL3BOI8qJpR3qUjKDgtFxJKNyu
wiYPf0O3FKDarxVjtBteIi8TLDmVjR/4xJoYGCkb0WX30E8itW695z9nqcDLHYPz
tC+6gvzFnZk7JmVMmVb2Eh4GiPcrXx73ktYgONvcfwqKqIKZeh+Pe0Q4Fv1VILXp
BMeDUGxqp995CZg9erSvLGRkq0WTVAULvBMl5gSsHplVGgNMEbMVeTw2OSNO79cB
87MPpnoiICmz7Q8VN4wjvqJd8GG7ZO1uWdf/4TfPUDyJGTxVI8jeO27Ko4Rb3MVA
KMaxZrNH0RFbB/mrWyepxfGoGHU5Hrcjc77aJVkY56Qr1xN/NPUJzVCEMSt/PP4H
UzeXMuJaJnbnPNBXlEsoF8k6beiJceNrI+0pPOvIri9DUvgfKga9TX32Q/uzHZ0+
yAXNNsqexcx6tf6TfcDgonpi3TJ7clhcd0CsrCgEqxqobD8IDBhkdrEw5ParOVyp
5seCMv8Fm8dBUPv1u2Dy4GmmDMmelcR/OP+aHgHzW9sr4Aw8l8ClSn5l1ukrLk+b
CRq7zq5tWA9sQynNdXr6R9mkg4LACx3MijJzO9Z9vwIYCYU2vLkqf/km5gvLaifg
Fr6W0qXxRYxYdgykC13cP1g7eJ3FW/6uQSL5PRACRtlPlNyff1pkBZqblK1SPlXh
Es/C5a0qajCLlq757i7hO/w04N9UQY9qgD+fYx3kd0+ZdvGViSemtcYxdQ3X1zWH
lxM0llTJZLhGOY5viV3DQmfD9KEVZqVkhZTdYjXaSQG7RuPgV+4Xsy74oRuccIMy
CqnHg3NSvh8t5Q9gRfcaNqYfhtxoqURtnHsATFyDOlpC1jRwOP3RKIPTtzK1pgVt
k4htfGv+tvVFV4X24wqiK04RVcImErylucV+lkl2wwRaPNwgxdsy7EeoezywU+86
EAMV24lS3mf7B4vBhzSRv7O6casYbK/qP/WZGy1ZOMBPTC+jnq7OreC/ujA3tEK6
a6KaU4buoLNNKsPojDn8wA24mRppOasAcNydT4JmggxjDulcxRZ4dutWTqidZ5ko
EDVgWBSZcGTdoj+3Soiw+hDBJii0Lj9Dh/1dnJtNTIv23tuF7nlZpULrT3OJbjkD
ModiG6Nsy3/xdbI/p8MwIDiuY7e7gOLWzBwc3yktZlDqB8TaBPrtccl9x7S08UtX
VeXx1F3ii4Cc/GVh8G4n8dq32LlLRft6uMFnVenkKGOh/C7Xt3YP/HG020Pf2VhD
iBBP+CenbUFdiiI0blYpLKLO92cV7t6PqkzCvhZcpcdBnH2HcatyXDLrNu128yRb
Co9Qy9FldHS2+gGlcX5mhOKzLRtRdh+064yQgSZPjTAlPFBhCeLejKsU+1054rFR
z8q/jV5XoRJtbxbE1wIO/QX9o58VIjJlfsXIF3ieiJz/lAL3GGdytgi1ZjEadlov
IYQvoYUqWF4quRSPLrjC3yhav5fMcotK1opkFTCfGGqFyyOAqaRoAh5TZVywIeN/
ylrQiqs3J4T4HcAyHQkawDgp61c2Uk22hdSv2h8OMuHyLcKCaAmHdBTS8GfMe7RR
GRRz5C+A6lTx8Sd7ganFYxAsTL6YuKOv0J0ovTYcKoD8/TaQkaxuE+mQNkBzmJxv
TBsSLJDUdSZSTVjHTQZMcfPTK1Dx3fkqHZecbaMmRqL+8nW8KPaQOjRZQ3ApHbCp
F8jqtvlsAmP2NbWtybjW5CdANjbpZ64aRrTN1IOnqf2w7tRDEOMkVLWSvjQnA7zi
L9fzQqa44RCN63szTdb8zddb0hPCn1o/DyAtRsbR+R6fw+uAxcWwWvPGcFvvHfgY
qPsTjeHeT/hTTyuZqIXg7VAj6q692ZWHOmTh77RYjl2CL3B1xFuribP2PpRbjuVm
A5t/nlZVazh1JKJrXY3+0lh78XUTec9xWxG1LMxhDEMBqpZS/QuEiJ0sTP8Ap6MQ
b4c3TfWLLc7kOogIset++MBukeC7+AS8qm9P2bbKKpT3Pqlx2rPqKacnu9h5klLR
bJ9fyGUNk4OX0QnhLaanUKQO4NHIVDSpNB199NsFDg1sHsBnXWYWHycPwigpsAA0
tcdQxwthFP9oDkDHPfLuwMGBMJrshAKCg6BFSi+APwswrgc4j26Jkiyj0dfLhyM9
7anaTyxdV6yYbqvM0nO/fJOMAAndS/uzI1/VOWxRGtSPTHOW0zeR8x2N5USE8Uem
1bKsNfBgGjpgv3r9OgT72qKU5H6gqY01rWr8ilnlU9oFotjYuy5Y1lgemPAyMhja
WmHMpY2dqVpw6Lx15nKpZMHKTE6hH2oDQqEF8gFvYdJ30jZN4Z0DBasM5DIlJrBD
XdxLeW22Nj0Ol9sFHOPqjpvlZq8UKakVPZWJ/KPMbdDy5xAjk+L9NmyBWOxouIHK
w6ZFwBUNiL/Q1RXZhA0/CMabg3b21xr6Oug7GigpU9tRs1EeCQBYf+OB3ijqAJSr
UikjQ+Pgh5LJWbO8qFKOsmg3zwn2DcA+ZVg3yXOst1C5S/5qvne9Gfu7FhvAdUgo
jLVVzQD1cQ+UeJdaDruHiurtU2jzjLKjCsveQU4X23uYJfbSxSr1tIIoxwZ2UD9j
kNSvtEVZGvrwKKWewsn3IDnQdul9bQSNB9rpl3ojmr1QuOiEXmXKgTl+PYfcQkoC
CF15PFqLo/5wzfwbtYEx1qbAzbmgShxamWBBQuTnGKbR/4546I7/NLJJJeLP0Adk
+E8WajYgHeatx+ot+N+nsZXyiaPen1bY2UMGNLL85zydIfZOF3pt/C8rTVOfQnVu
eelnD6OjX4ug3SscGi0uvvs7CelMPj3OtnTZU4z/sNpogD4r6ua8EVgN7t4/5Iap
OVpjC4GzQy+DryJiaUvcPclNEVlUptsVrNI1PmjOktXWVMEC2h3YHg1FD8ZA7xRo
RVxtxhs73fpriPxJPz1iinpc8tnjOB3b5FxkDKtQ2YiUk8IfcpHggu1/eMAUD7Xw
AOjBOE/6q5gNReqs06yBGbD7ExSlTgMjfuUv4zcC/CWbfTg/7ifJjkf7IJoaZAP5
l5bgYETsmqS3+QQ3OavwCsSGOmJD9ID3Kk/A8JtqFpqi9ty+FDOONEWV0Ua6c/yU
A52yhLewjdmELgmc3ZaBLoFpcL3odfYbWEvVNXUcIYAb2nXzBxhSO9xKV5bIk+MJ
DvFMTESfRQlRZwcqSyMml5rCzLjRisIHdJCuwbPAjP5qlPFywnR/6tNNAKZJNwjE
f6CEnea6t9KOjH95s2YWZ6i51jbs4fVMfY2ML7iwdl4ya+yOufssgP6N0/0JIVG+
ataZkpzYWTXXybc3BwNtzJc8ElbHKtGOkbmhp7vGH6jZMMVCnvpQWA0OvmOZ37oc
qaLm19CL67HDZJrPsjvbRPbv3k85g4A8HKQf3eEKTCNpjrahNXkuiKvmZRyl1WHe
4TcCwLbw4yRqpzVcYtjM71afE7rWNbGbucQ/RwkB9URBXwZ8JhfWaEeUQ5uZae24
ZfKF7s+cpkydjJ4AeU0HoBUMN8ZmifcGrQznP2ppZjTFG46f2i2iO8rRVVwD0X98
XXSDLpyyu7tn7lypV8bTqv+PkF4v6OsqYKUm02WogUSt4dJIDmfeDQrjNUrNf2vL
3owC/VAy3kFqeR1z8d/ZA6CmX7IFcBOddVpIDkW8RnYflF/aSjrp6oUO0oL9Xk1e
LmtuOW4v00LFqKVj5rcZ72rcjGkKXvBGilWO6tzlymq2zv+R+pSRWWGUhOw+EZvr
voYXz7nkK6G/EfDIGmhmAR4qFBkUXUBmTNdonz8wTbT9AGhhTm/YZRGv+2vRDVEH
xKWC2QLKY3EG8arFozCZxmJIAjcrzHUoxrPLkGV9WZcYsALDxGmioMlbttdEbnpC
QQ5tvy6xnqmRbBAf88EZIsoNhWu9d8iqTiWyFpjb6ltc9nfzjIS7BjgFSfKRl51R
Wt8NdE/lrQQ0m53E/lkWZzb6gNXMzKjCA4AC2fJz97Fq6osO7uDtOcehZHTC4jz+
lU1HIy3sUKEMT0TLFgzAzk3Ni1AYneuryxrsE6DtaCYS/exqv7kQpQosCihyBPCX
ulvR7gv3wCus0FCwlZ58La0ktTHTcRy/a1Yel3LxNZmzNQLur3m661Lh0gdjkwn9
loETTOpIHD3U7GwPyyiP2Pk50oVOX+8bg6/qAINAfMPpki1Ak3ic1tqnoGifa/XI
WkFELfrkStVY4XXf6ogNfO8Pt49BTfT5Gv0WU7GTmp9YoDH3lflZsXCDaCDudWVq
wC8l5voaoWuvjWBQmkjrwgbIYQtajkPpAprCxwMamC3Fyy3AarmPZMWTCh08s9u9
DsKwJivZKLzkEiiHAavrl7dk5komIgMUorkFiLyAJOx1UdbSeSNIp6P+4s8u9x0Q
1RGPqpKPrpWbZBu6YbjhVVsdjIOAV1eAn/+YYh+aARiIPRs5xixc+KyELFUk6w2y
G/1dLfSojHiHlYnO9vgB5JTf0EEeSppk/YgPvBCcxppYxsG5dfZ6cp2AUK5GeLxS
Xz5FFrzT/dz1P8a1T3WM7B26AEblBfIF76HjgjJHGrn0dBN50qtyx4nI659WhHUU
rSpaNRmdTABR4mJkZNdPReLSLTr+YSApr66GyVHOMrEd368GbXHho8uyRCB8ajTT
Wz/rjl6CLUBb2GPDZASxQ+myRBh3enJ+jBcKb8mHiIkJRVAHXiYvZ72Y/CBcXkAM
PmBDwteSwvCfDjtpbhaH7azj/pKcwOHVrW8DxtS+rfUJQ+wNNql6eaqxffIuFurS
fHP2Qp4Nw3ExE3QrYHDAsoQ8ECdR1m8cZH3GrwLNa8EEpM+oVQ26QTv8DiHrUosq
igqLzmG9dgHPqeKWTYblu1RH5ojvNwUXKzyLNwgD6eye+BHf9xm3tnz82zkD3VgG
Rd72qN10JRPuUCR+n8Zz8i/PPoHjNWACJws1G7fbczfshWMhcB+dU/o/YD/o74SA
dOty4luOJ4ymoiJvrKacsFMK3QzRb6N+KEgHkvxqLH8aneRaH/FpVAJl3wnS8Usy
GWw9nRR1GTtT2pOPXsbCCoI1jRyHjyqQGmRN6j8qPDyyCZBEVzGYTP/07uUJxhqm
Vhe8k6mBNsjo1dR0ZfYuHnTWNbn5EuIayiDCAQAp1UQkdkHLToTgD0AWTrBQfqFX
+hekpnTJJBAa3MihO9mwcT4tWyVJvBvfes0m2N22DLOx0xLfurkQ10HIy6ksuVtm
Pr2ekmDox+6nr3g0ZwP6L6v+EasSUlEXYr5B9+kBcxMlFe1+Wly+E4Rc7wQT/0v2
krn665GR82IHzL4QEwNlSTn9rUKmAjLBIQhPhcIcSSPY/u2KIFQbqHGs6J5Qhj3i
ECl3EHYHMnqtu8J1JTsPSfP8pn5d6a/tzTR5XR8diBcvA9sohblshM3AVMogO5zN
6vmpsnprcY4dnDBB6+qiuilWBPjd3YWjd8vYAbZmoA270E4a45wN5VN0picaZUum
`pragma protect end_protected
