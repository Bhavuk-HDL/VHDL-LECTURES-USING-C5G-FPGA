// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:39:03 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
J5FEGucvIY+EnXYy6wkOZ65XwOGACSpLP2zy9r//gKHJ84np39ZuiVwTK6796y3N
QJLzPqTSw5uAcdDi0LhSbbG0hUK+ao4ZzRAVIfmlpTaS1+p06CcXc+74zMcKGJCR
E24qdiAEpJO8UnebMEmwNcBatTBBt8HtY73V1EvjCu0=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 48384)
X1j9sK/33DmveZhlak6pAA6mutIJdkAG9VnqPXPSEteaEVhmvGyuUR4xweKqxlEs
W/jrNQkkemjTYwtu3wQ4LkHnWiG7IX5r+O6MPdf5XsdK14oQi7SUfoCNNz+XHC5U
z0yFu4cSCLLgrIdVQLubmkItluvVomkww/p6vL2oXI9MU5II3GCtr9PcwaBg289o
odVjg01JwQtrIic5DGQ6XvqV5VfJLDjhfmaMkTeo7bHQCeWfw7IsWLCO/JMCkYN9
GASn3eZlf2CjGlDY1AUe461FeUvqB0Fr4Ha0/Z4bRdxO2GPbwLQH8zoKi6vXtFqH
kApSu8uX1awppSQAYUdoMcx/icz2fVfxCiMsbZyHbbmWhD2vImCBJnV/y4MBtake
Lxmp2kVpENkiKTH27NNLSwSsQi4lZuvr+xAhdbkXijJyeUUo8zTOQ1MXUIuygQnE
N/RqBKG+Q6PRi0CoPNwBlzjFeNteJKv/tqyo+fC/YZnIHNMmpD5IY1v6mxVqMBHH
ipAz96Ou+kVeXXqJFJpqkQuDWdNoTtpxqtsH4TD9xO5zVemuM+AXUxZcSiR2PICY
YXVrZhJyohJIIvv1+2mpoNk79jrix6VLpFebD7qzrbaObTyFAqDz/JDC/89nk/hL
5IZgoeWwyGRah+WR94mYOIO2Gv2baxgl5kvBHp5k4f/7lf/lrcCw658yRnB9A5e3
agAKZ2VpC1O9Od8T4W/KnV0b1AGt5IYpKhWFWrR/UeaEBN+4CV1JIfFiY7/rD0JR
YLIDvefaX45nulq1Bm4jHSWStGYzpwgCiNNgm49gb5t9orarX/Fe2hZn2Ogx8UrV
L+Dz7MZvx8FS3NKYrUKAKoNLgVBDpbBADeRld690Mtm8QLbbfAs+6TTWIg7VOspq
MGbn/rykiLd8KXzyL2jVgSnUyJ7/VNEEKUWiyo9quFXuAPbOrKSpwh5oP1PmHxiH
PE8UQfbgqGaMRBrKmZsfGtfUQFiu7+iNKrN/t5A23LbdM3AslLI9ZCx5W0poQLlz
A64IcEvQ7Mp0dwmJzrsLmvKa9tXJu3IduAWKQyc1JeMFEXVGJfCOKLC6y9hMAl6P
xi9lNEZAbMXXDhiVZxy55qDS3aEx9ncD6ucXk2TwxfArqB7FywDwEO/VUz8HeDcT
1PSsR3ck462zIWheU+phhC8QeesGsYedCzoNaHgxz34gNV+C3rnjEtzjk9CXHAiQ
pRDpEDf7ejWMc30Hdqp3xebpiX+M5d6GdXZ4J0iwwfggSzEXnPux+M/ljZoQ87/6
xSUEC3/j4OhG/fCfN7vWZqJq/1lZDCAH3uggYqBCQ0zUPEi8JTtQB1MtWUnZ7LBW
+1z3H3yW7HTA3lNEA25VVlhAa11CDjOBC93Bo98xdAYWV6k4OxucJP4znboCCH5C
PqL3DvXmJv1HLdxLtGuwaKjhZJNDI7yGeBPDAuBhX+r4VoEyNlC+y5PfC6ecXG6R
SAZfUEAaTx181DHoqt+GLSRJbN8qDoNQrs9wSbrjZfNs75AqNzQ1TuIzwV8sgXcM
jltKf+4iCbbjqXEUDOd+IqYnzrYzOwBFNZxRfaC2zFsJE2KOKkBFuKqKafgHGwcP
djWgtdUlEAeBUwGpkqyyQ/IjlUb1ydUhF4HfF66e+KmooAiLOnB9zLHL0eU1rVbT
Gzjt3KufSyMvAm9U2Vr7m/5pPVffACDdGH8jjHEHUH4kh50wWJCkA1FvpqkIhEfD
N20DeNEKCE+xVVgg5UTqphSIbXM7+Ko0xNQ02jf0NnXSPPr2Nxb73YzyvCH3JtH8
4Nu0QKLL1ErDZk477X3WRgTU6hTrmULqWlF3xbmR7Ti/VRTLPU5HGUinTAbLCMvk
2aicLY9UHaCWm7dOIEEOz3JOOG3SsnGB3lRbjBptGtMBhqGHR77kCtfLIxd2xTHA
kKe/EsG8oe4EJVN5L98yXVW8xZ2WEXLuPsAJPSs2zK4rmwI10y5iByuYsXVSa8jE
Nx6l9VI1SR/9mjkflVyEOc5Ppb3A7xr+tuw/hEWSo3UopnFlwxdU57VPg0ULicrN
W1fLbFmcj4ZBuJjHJ+4yluktBr5gwEFrZaaVVbePsIySQ6ZY3fuX25A8B3e5e6GE
S+KThmJ6yYDh41iWBREpKNtVctZ+X/XMF1Kfn4bPweqC5VcCkGovDv6ag3ievyza
myzdgv9emM+cU4y6mjrEzZWU2EaCO9ratWaYrs9p/t3CSe1233Ic0/QIgYF5s/kS
cu5j0iFth4tUpxqsT8Bz0meOKK2HcnHFsY5IX6x9/VcaxttEhpjtAVJDm5VW/MVx
EHhbnmIB3552UvUl2MDC7kfFgA+A2OKIWYHQTXh1pgaON14YhNbrpEq/OXcKLHTM
0Pcjn6DLLNnUYbft7eqq6q7qduDFY4Bl4tLhsuuZegApFkT/AoANlqpEarfbMzLQ
rSgBIu4WfAk4gYrwY7d7OcpK7gfDLwkYKCXDAH47E4BK/E+3ltsdHMq1zvLIpmDH
HLnnYEVwRiXo8iRkxaUUSK4BvDBISehb0QJGZdvNOOJZsMdaiwjHPOmGEhsTwY6R
i6UBIax3HaHRU6P+2/hpQV7We9MbNOojbTO9biPe2tl7UISMyWjBvWWsdL/WIWHy
6QYSlqeSsU2rqOYpPS/0Jt32oJvZ44/9zRfGMJFyGvhW/PfPY0uVNbMaMYqzgAaH
X9m3AUjDi67wRJMh+6v4GoYCgWzakldZYeJ1yF9IL4Woa7JJJCU0lA7zFhTDBw2x
3E5/FtzjvIsLS+W2S8hPbl3yNk7Al55DfpSBDhgPPGT2X2YizvP03PmtSLbvFT07
ZXCBF3n6PBWwN3S0RSnBE14kul25TvqeWYOhF+hRLgAaoFqGy3MPZvqDoXWLXzD0
+OZ4/5SVx8mcYdYCzhuEbijXOcG7tmzcK/ztGpriS6vAwGFK+nduASGlQFYh8lmp
4oM/cvYMJQ/sphUhFlFkKH0arAYkr2LiPA/P2n0LhBoXNArrp6aOLMVnwZRjoo8e
m2sRHg/MHfJ0oy9GeMwS1My4SVJD/ZB5/BfZOlbx1EmyHRyKX9sSbMeHhQCuLCaR
DApDdupJcDhVPRailGNrX+CzOz5qwBICcDsrlbGnXXdZF3pqSgQ8KGlDl1fYXNwK
R1IiAfL6uff5d2nrgU0xU7AfAMB9MEMQEO4N7c9P55GEEtWI0rgRNMFJ1agvd0HT
C6f7TLwfwt4VXDhjQKzqM5b7tcHUCqJTobZHBk94/XuT0IixR/WXlmYLEeh32qdI
v+30e0kFa0swGRaDBSB57c+uqytlqy780N7gjWoEXlb15WkIGdf0uvaCDX/v8gL9
FxpfoSnMLtnUuAHPp4d9xUNIETLe6sb7lVxisF9fdtl90jYf00AMWaso4EtJ6Byg
8oNkcaZBL0xDbyj8D2wP4q98s98lGP+MrQxnbWNeu/UaDOSg08lXiyzi+9MIqI3J
C/ATMP8JTV4u4fRoov1Fj7nTIyyr9kg0ffQUQRL9GUGSKbjIXGkEdPjGbLoaJXgy
wKzLq/aus5fdxRWvPmxNtH4MkwQSQjU+KjZfnzLODeza7jnJYAR98KBs8UZx+XOl
m4sIWQ8alwUVWVAA8by+np1ntvKHr6jF+U+UhrmsmZQkBq81QxvxZ6e2SrxuSfyS
nzobZKRdXb3f4WpG1LMWhVTDlMQaucdu3ulCoEiPCrtHd6I913qwAJtDkAxSZDqK
lqQMfg+nnQBF/99lTi85dR7Dp7jWIIGr7D5e6gSXd8kpJpy1lebX30OHdjWn/zzn
c+4MpHoiNG70e/pDQATzHSwwHmvozuGXnIfR9C4LlXy7u6NEfZCOYX13nBMkTvRG
HEjm1lgBXdqA6TYbRIyk1AY9dBGIKQjd9g5ORM8ofs1miprnO/UAIpwPrTB8DGGt
7YsKh7AVFbmUNdULscSt+IiNsMWZ5SGcxCOwtQT+tVDV1fwYuVqL825oa8JwAoEB
1PLJsRAK6iAbemoG98JuqBuoROM3mnCV/N8ibv1DgrFMZdn8Zaab+AmFKEaqZHwk
E366yUC/dxTa/Oh0yOsEgXfDWvpohexeSPLPGlBlSiw9NudFf4U/r4hMZz9Tf0FL
As4FpMRPHKdcU1tdvxWFd6ZL5oQt6cX+adI49TyCm1/1MsMjQPqgTqe+2p3lqKfz
RFTb2T84kmNzfklP1BWd0EhJQwVQvhaJjd/FZDwEmTatNCvkJ7REH84893jkOIg5
es6KImtunKcnvUuqp0o8GN83KpDZzuDBzV48rKqfSLqudg3f3PweP6WaVz1aYIxz
KfZUFnSKypILr4GE0l7NJhJScq5Cy430fOcW056nbq6BkXHZLQGY8BSFMmWs5N0r
gutCPTVKJ+8mioklRNcoFZSg683CwrLpx8yyOj7ba1MSHNdTbSipSNSr6qG4AYfo
RHvI9CMTISnbYN26R01x6t2p5FSRMEZliyUlt63gvq4qoWUZDGAEThkBArmngqC7
8mTD86zkUVz+yzjPGP99UFWyNfYgfgWkuCbjK5fsRwyX9oyNBTQQw8qTfWbMu/ue
E2cnZ59G87NCnf2/0h1wSazx/HIDf5tBIQpsDDWRw/uqFv9PPuOZx0arriL3qZcQ
lyTJ4q++lEvfn94rewR6aWte7SLoQC3gkpvd/r5Mi81K9QVYbtWs4wcbfzJU/mrd
435iBgnPpnO2At/lP5pVZD+/Hpuz7U0Olb5q0R18asB6hMTHewWstDL8LXMsGnny
CYFRryJdHNctzGJHeeILtR3/2h4booh8h6RyXyW/jQbrqbhYD27UUSclRoGn/uBt
5n95adGgllaxSRCDkVkVxiS7ygtBSrKtNBMYsPk381CVlBUaVO46by97X3ZaBAhH
6Fzmo27WmiuoNaHKTR5q8ZZbVyW2wDiBjMfwaTqBXcU04IzKwzQlAwgmEg603koj
HMngVyfRTPoEfCBL88XqTLTPWXUlK/yWHYNCD7cIh3wZvtjiTjwZ13B26BjWykC4
mM/UDEXdj5YnklICyannAF1dZLsxxwYSedjf2TLJ0mcG76SI/eMoPkkNDLJDLJFO
0kpDGNJzVrrnSqtSfMzBk+5CPiJc1PC2zsk9gIrfq8loGyDi0NxMWBDlwVdoWZ9M
8a7trDWU3GKQ5ig3a0uB4Isz29uk8f8cFaWZb746h3Oh1+QDqNo0dxi27jzz6QQz
Wz7J+kyAPI8xQtgD3RpVl0/SgmmLO/PYi12ITz+64nFulSqOr0NxrbnpcMnFeWCo
r5ZhdkSU7YoTDAqBNMGlqY4ASS+jf26gAC0WxV+MJ3Bhm2WtZ43ZWvjP5f/FYFsO
FcgNbIOEH9wise93jYTIR1q8iHpb63ub9zWZYI+OSOZ1qzAeAz0d3uXXQIL1j+Fk
fqnZNV+HvwrOaDk63vS2Muy2NLcpglP1pmmNRf6t8tgTTVU8KT693EyqhQNNcNuE
tyLRqjUYYLeU8UFaIg11oslo1s4CAAQXckKSXUJEYecroGr8CtZng/ws0Oatv6xm
bEtq+qudHQoYyvmJmJpmCtdSOlcS3suf5/4q7NAqZCNLKfRA2truHAO6u83QomSl
yPrDyWQy16/Q81t2ezJB91LzzomI5eHKuqGg3bNN0MDz4cUAdqD6ZtljDfCmOQjU
28IR9RSAC3bnv1byqDsgSpzj5F29DuBe07+Kka+XRSHLors7RSXnPOoifWHQ41UW
Y3HIXP3Y9YxKyeC+M3mf3Mw62CaSqqyf5FJlfXjE3mM9WsgDd9R4r1kDN42WsSYf
FBRXrTnzfG6AdEZ8J9gzXNDTkL245OO3x7Ja7hBd8WrhuvBTc4qnJ1tAK2ktQGOT
YOOAPU/9dqyRkHsDpWOjK3VabCeeAie4OGqKdNzFjQUQFM3h9JlH86in++dP4yua
RtFT7zNZTTA15XETxls+9p46eMucqw6vykHaFjUtNYJwEVJFSHB4OYMu40Q4RGRP
YogYFFVvMgfxtE2Mx/vRRMFWzrI4kOJcKak3lMH8Obw5EALzN5pn/Ln5fHvFu5X+
ztyYme9AOHnIvYRFW3FgoB1YQS8SUojpNBTATTz71jkUuoFl0q6vkTGKEYc5nb9L
SfLlNmNnUwteD+pYtMv2S2n+6QnVz6VgHuDtuj9l3MrPpOyRjxmrIvjGcV6pJApL
XTCUT0S6LxBcTZq2cg522IVaPDLimHL0i/ofKn7R4+mWKB4BMfBY4NWXoH2udxoy
Sl4PS2/oyNI2wlJevGsLcHRUR0eC30i5Yn2+PvJcvD3HouALPtSx+ruGrPEEQTjD
sfiETq9iWP6EHlA6ycOyKaAHC3oiR4sH59pLexI6U06KBJ1orEwo6G/Psec3Ii/3
TMLvYSi4UsULSVnTiEw4YQpn7ibJttPgaFtwuBhvbOIyqHXNR7WWn4ufA8RuAXcb
qdpf6kG6JGNuf8NqRWTtMLAUiZr7+z8InLzcpI8X3t2re/pAwino/R3F2j+pHmZK
fd+ImNGnKTsqwKqx3FU0rStvmJbpjHrhdhYsMRe0F9AC6SnzRjjQ8kTtO93IJYGw
+Bg19EPAQZaV9Le5N0hGIAyTvW0NA4eUtzlnfByKLHx5RtHfN9A2CVOta9N76lm8
gNTv3568HsHOE8zbhpbU/Rkusj5XwXPf+p1x2uxeDxlkGGWbAeEkwsoZKSvTTrOh
K0SF3sIhn7+9k6QHM+mcGj8bcV4ICSgzpbz6wYv/MT/y0uPbQj2zDWdsHT0p0iHG
fF7IMfLlemdsniVY12uRueR5wwEczCUdYgOqzV9zXTKccIB90qrrqdBDAlPrHvcU
X6KAZqnkTQC2zbpOWYMyeCpTOLSUJxuNSh7V7lv879auERTmdv3Khkc4Ro1UCa7U
ytTgY2B/PIoAnUjUB8zRn1w9FikTJOGTtQuR939/gIIBVknBtc2u54qyGoPDrGux
oOqPQYdMrLWSdQsYu7YMiSQ9aoo2KM4SnEc6Lso/xCpo2WQ0dulSUkDNZFNe1W5W
n/CnzMjoRuiulDcVC8ouKdOTaXUelDTE/o3EjeZCETNzulSKM6YWsvwgeFt1l847
E9ZgUybQ43yQ9gszBeNb8DR5fw6w0KUEIg/woSGFxcgN8ry57yA6zZznjm6bAd3p
71yIpRsIc6KFxqFoeVYK6F8mGfvyWojyDR85GAVEKJZ7ybSGuPY7uzq7MhPdOLAM
Y1AOHb3d7HtXIjJn9b0nkbX4Ulw0+QDZPvy1FuA2Q9iSFbzEAIy44CCe1Xpf9gUw
dzTzbWWgHWOiFJDCRx30GyMBG4GrLzwZwcqVS/YNDSt3k9oazHA9sHDAqOacASc2
yvwl3BZ2kzl5LoNnmJ8mPbtePSpoayjuiC2E6YrrrMjozsL6ni9JUBvvroDiEddU
KIJZCgQXXNqLHY/cblpVpASDe5ptosAIhQGTy1JmTGY6lEaRniADM9wYUfastDra
4+P9xLkGfqwVIRlcRLSN2tBUQmbjhKZVwZoHVMVR0L7fVSxvHxptfokDrK4r0ptP
cwjE7KCzAllDr8atjX7nGYPf3YoLl6mn7chXO5EKdthQbnSHkEb0Lg20/0wtIjti
qeJualWyRzo9KmDTkcxpVQ7BhlrYoZgiynZ60wDbRkVE6Adajh65pwrkdewS+ahP
1Q7PSWLnwV//j5eRiHf2/TgRQ7lpNqzVzCv/8lgMZqquKIGKjzmOu1DePxqzFya9
RIgNrPek+2ud+iyPa09MGJMvvjx7gBZ+7JivDwdfS79vB4Yxumys0N28p7xVNbwF
r/CXTjqP6ghSiXyqZSY8wpUcSIHGRFN0uenqkN0bQNLQzghbQCST5sxv9cyWPHDE
dKgt9kCdiH+XUqXjXpzBLJBElGhB+GmhIEY27ZYGWlbDkJG6JZ6qtQRJpv7YTcdR
GAopUuMigvyW88OJUwNWMuXcDCpxomCtQJfXA241IdPmmlY3oVAAF4R1kUMv95Z8
MLcF6NZQCl3i+t4CN6vWNP8tXZ2i+Qyd5GS5rywI+lcBjfMWc1hqGeYgADMNBbge
+KkPHS87/atiPmXKx+tdHt7DpVS743s9r0y4kMelh5ZzJdDlulYcpbupWazg1lMS
1OWq+5zIq2hoq+gFOYW9g/RG5KeZRAviXklT0jakV+F0eSdwZzy0LEgJ6ARJ/S9Z
YvUTw5+btCt13rt7mffbpXggPG2DB4eMjx26GWid3Ep9XUl0E1c93oYcyEFEj5T7
io0dJh7ytofa45YZURwhstTA2nPiVsZr5vLxy5mzeRqx/kH4nyvC3+LIiiXtOdtV
gSS0wOsvgZDBlufSMgy64dhpfkGji7tb+/pIJTFNlW+pZ0a9oaYnI5iYlTs7LE51
BCRToWMqitL+E8yqhcDJmes+QMcci4StlL/AYXlHI72fPI43gN/TCnByI4TOxxqm
rN+iS4u8bplQP3lJge9eQvMLuySHK89CwDJpAX0o4n4RF0hawCoZbCIHjZR9LcRI
AgBT0v/zK3bf2TWfuxq2e4JY63F4rsKrlFLTql7Xvox+GkUrka4c8HABrSGCxkMx
zZkoWw4fCpWPnlOlCmkgyWCFUl+TxsS5VA8whHeERgvQxj8LvUOtTuIl2BlmwV44
1eAeNBSa07GgQpAOQlHfEwN1H/vRx8mRYywKY7BJDT1qCToi+Ggwaf7bR9BkrqcQ
SVPMMAaVUm5XNVY9yI4A45eTRzpRUG8Zy+cWL1COfXtveKBvySYBNERXUskwM4OQ
2cN7QqTnhiM/tdO5v3z1XWq+clxQrg50gXCsvlCW6gmYRmnsrHoXPCcQjaGLDzST
A70QsyRR8YVxH9+NQALzw4yHJsXYzt2/ZS5tsvUMO+uTcNWI7mFjbeotrmhVYFVi
nASCjNwWJmonw1FMnoZYwVeU/Du/1ZwxKe1rfMoC23v1DbunucZp/6P+tofnQsYZ
aCCAUNMxPt1g94/JcDiYovUjyEhaceew8Nx5iv+iTVPkz2WM3b6W/4xtda8vsZOg
ErGPc0hr1sd2Ya7rQ/xVmmyI9IHjQiXxAx3BV6N1QWLmgB5e65VOCU+BEJVE4AsZ
LmvC7k1M25bLrS5A7N4fWstMFjluq0QyZ84Q8WWGUSr04MhJNPJU8IYRsbU0hXfW
Hmdhf/NdaIKCN/91yqsCTGeDWsMQcWNd2a97i3b9GpaEi0LpDLTnmPoslPmP6mSJ
H7vz/HSU8a1ar2DnnocP396PcJizt+zyNW2BLLRU/sMoDraHyfOnBUPwi8CTlxzY
QIhKMB+JaHZzDlhBoXQDpZwzqMwjzHmZHUKC+ZMEfwp9/OjkH831TdyNxUXfzHdj
EQcFFJJihlMB4+Zz57PepACYK3wRGYIHJQukM+QTqZatxAJ6kkhN0vykKuuSsMGz
m2NBYR/uetjdugwNWrqKJgRE2cqju2hsFVnHdVF3htqgxDi4ouhEMg7w2sUypvy8
tR0DNyjG6k+GrbbHDxElImMP8w0xLRBxh6fUB0ti+5SRmxBWWOQpFEBkYGBlXCcJ
ZwmcnwpKBj/T6c/jRzIdVOBiCOcAqNSQRVMqYQPWzM8eINEc3Va21GNYzkOlMrv+
9izLMxH7N2yhkL83XFNgcOAwk3VW7fwrUtrrvtKfmtxK+M0WZvEfTkaJc1YRRQ46
gKO7LIDQmXBnVHIiGy9VAySIUE5cZFLDJcL1pL4/8XKek5yvpGPKFKUFxAgGLnWF
oZu5S6/8Dd7lRrCq7A50vhoJpApowKFlNHfmjWAiMT2FQqC0uSjfsFXGkD8yFF9a
FDbMMYlys+Dct9E2TP3RkUyNMUksDkhSa8zXR/5scwlbzgnfpSVsEIg0DaPcJfPp
+ekKkxYXrx197WvLejsiGOuKdZY2GVd7Tgd+gDzbThLMUzzsosaM+OrWSvnIkvTn
SUK2pMjwqN6PDQ+F7XRDpOPOQYKkBrrAdtTuSHbR6lQaB9D1oTsUc4Nma642in7c
Tb0dn4WDFkUoiI5r1Gk9QTGWM+1/eAusKQfAe4ckA5W5gHLI1VMwm8NTCSG54dDL
91fz5telrkdSoPNCm4y52QSrCLlZv6doqWEHfWrEsblJUA1aKJd+b/jcCT0W5s+H
MvqN1yf3Hkf6hj18X0NXhn6PVQbLwfqQ9AkjTh+gFsNJGhT1N4Aq8CFFnDx4Kpaj
Q3KS/WzL1N/gP85xI5wj5Uy5J+3hcHbeXhUgGTNe440LTlycB3z6oRcAm6BtU8Uy
c5wGXJ7MrXOEkEtb0ghjQSVZEkgJYsG1b3lfzDskd37EqN9kJ48CaQjgPT+dI/hC
n7lK0faCSb2cZzQKC1sh/dnyQ7ww4i+AT14OWmaTXCfssnwUMzNMo8qHkF/3+/hO
4B9Z8YXlWbbUP7BMfHIHThM6DGvIZriYPr3XYORMLlsRCvA4EIAh8gNZP5ZhDbjL
HGpHK6OpKFU0iqxIH9BpwnD4Ec88b+oBzHsolJIF3f9gsdJLOhIZVKwrE+Or17JS
FxOCFYthUZng1d5edPML+u5Cg4ueJIWnQ5NXfe56Z0XOgl8AWGLUA+05r1eTha5Z
k5zyd0r4D3+9ququ7HIh9/f9ovJWwQ/CR4U8LwpyI6P9tdyg8xwRkIlxecQu8HW2
Chz/k+Yf/PdiKyZYD41xhGxY5o6j8DEwLH5qOLQUoSlF90FhXLeIiYHyReml5/gU
akIt27jzMSYEmD0XWMU9m0Di6Foms1lFF3prwvjMHs8He4L8lQLCueew5+UNjxfA
b56ivHSKx+1F7jTwnJ2qAv8HtT3czoR5nt0GjqXqPKD+6mOOGZKIsbSaAqXq+DhC
bkCw1OK1BizFFbAjWDt87yJ4pn1o8Ckwv/2vXRZTweJrHBlXthe19LIS8LkWFWIY
PnEKayJvSXkrXhUvhO2bbTjNgOM44lyF/I5uDrV4Mu06qw0aeuxnvJhsQPdycAXN
OJ0RxsO/HzqTH1sSfhG1Q3f5mQUNPfB9QjnXzG3/tbDptOEb94mynINeJWIbJGKs
wyM9tVEV+tYaCGtp4IQepRcA8zZeOwlXCeQ5e1xMSkSsdEA9NLg3/rueco6sisWQ
yoDSqVEPBnpcDDzMYTrD6k0/YXwAZ9+o5LfYLFTf9kpgyP0fnJBX2VF1jyXUs0k/
9frFD9+bgHP42+5nY99R3V5H4gvau8pQzlSJDG5PZjHuAGFAWUmj8gdKqi+YM/2x
A0CF5Z4j3urYwKA6TieNbWARSQYNeYrsWuodgO8eLJ+2oOA9onz0Liil9ZCAczo1
WOD4g9dEgEryFnBsFRn4ZbdyRcz6NHx7DSOBK742TzWuZVZDmQEXq1yepZLNW37k
9WEA9gl0SMynf84q2bnCWJMP7RIDz42/h8pyoch23RbcOuYFzxC2q/dfcgQEYae7
0IqxmMNasPQqetohZHlCW2xczK+1FPNMx3CFJ9OH4w9QykLFPq5+kC9JEV4amq5j
ziQYKHXLQgKLqS6xRHLS3O7G4CCfMoTRW+1iEtwM2ZiWVLkqxXRG5Rzf4h5PJgM6
POkv6rijq6Sp+MyNVXbRp4Rme/8IUgDTdRI1uyHYsDs/DOqF0+mzNmm8IoremI/Z
lgk2Yz6hc2+vzWiteDaD3O6E+zFHm/gFiv2NwzLTA1d68U1BGuNY297QvI5vh+RL
hy0ByHEp2jQtVEb6LCVsN9h3e/LehTaKbiQrUlz1k/86+xmKcBifzgNVUVR2q61A
6+nYSbQznCky305zAEvD16wALyByd/r+1tOOoAv2BP7kmsW+WX43s8R9JBiophH2
V54pil6OKEcXMuNQ3O8jKBDiDh6qdNSyOEohMeb6Y0JS2XvBAtZyy4cJxReU1ftT
uu6X+Iy9XWD3G66xzUfFWNy3EdTOJoGHkIZRjvJALtw+lQqP5RkQhyeyqhSeIQrg
5zQ2cuaxnGvRE8tDZW1Co5shZ5zWyzQaZUhX2JjF8fphU1FzSe9zRFjX7lO0O1G7
G/Fv0V+fYF8f4t9LgyCUWK/u+fASEEIxM0xIdVu2jxr6lg0Tu8vgZdFqF3uXvx5V
S28rRa3WnopNceg0UFZhd3GZmSGEffMG/sEmoq70iLzMptsltLtQvm9eCksxjc2d
4wHBR3R0Ay2Tr2GmLdfvpXDy+LLW2nlpeHx2A4nXbTYFz9gXDTPqtvPaVEUjZFrm
Ue2y9gyb16ahWDeudnoaooFUAF1NIl47xZH4FjXj99SmCbZv5Vb8oyt8HWr2kGt3
b14BCchcV80roY0YpUUUEC0K2/bttrqkZ+pnUP2sHAKcg2GBk5eLQ05nHnh6Ji/2
ws2E+W296VJmpNa9lR8df9dt5XYjFzZ7Z02KvhWaZoxl7r4JRUsoe2Vj+VvV/BOB
XFWgToMPqZu6LlGJ0ENJG2Xr89tw4hwiBzFANfjCo7U1Ar/b3NVnSOcR2CLoIMja
jnQe8NBb5/cakYFNuDC9tK1F/yf6p8th+dymMxsb9Ntm8z0+FRsdsnN6TlbkpHZ7
nZTMgsGkbz8I6lz8KiUgdsF193UsFeua3PJggl5RVZnw1JvhOwimn0S18xDHV9Y2
ZQiimbbGy6PCxk0DTaASNN+A2KEYzsZ75wBuaEm1zf3WLsV2UYHa4rncbCKiDcQ1
SLFc6lC+hz9/cN3B2gEKI96wTJTofjXDFSyQI/i0lDfayNeZnN5a5sHTC/NyFmUb
sO2RCWZSyKxDbnGuVkjkqXFpkjt3ruNOrYRmqO2Vw75ZTXdlWkdjW2Wv9NfApAnK
S5vrlX5QE+Fy7UvMW71TsptRZpJfY1nYI/2/g0HbS5r+Lg0UbKT0wtV79yFwi9g7
vRP5CIwxn8zDxbP4kqEceZ16oDUjaj1EVD/df3puKPny1UEKr8Lf232QQ7CfmbCo
5BAv+jKcNGnN1AIHNFIywGtuQeLlL/4Ihof2An1O7FcSX8FNzb/te8lhhVrLI8s4
hjT1emJmjgqoRG5zqWJTkIfbsjiYhmopCol95soRj5jRHrcYTFb7XwfYxvKaDRYo
//QuT53InfAdqWee8uN7fcaCs89/ZX4HwA6Ihu8jnDwIpZGj8t8tU4p4JknQzYIC
R8iLWfmeo3eQNtjpaKmBk5wbkLtGi9bU2zNfSp2pRg/20/jhoHW/sFfs9AOtUq+s
snd1tBQa6dy+qxxD4L3DDokbe/Fnb7qFOQPb0O9uBmM70+n9s7g2fevb78B5Z7IP
sM1pZR+RUfKZov07L4ZB9L7GfZSYmHRz5QrYRL9W5KFQww4cGJ5Tj9YFi9z7qb0l
yZgTB2zGV0CNVyAxWX8OolQQcW1oEC+m8tb6MvPxpdgOAIsrXOVhoVYCVJ0fDfkC
HM8Wo/hLzZtLCHsQRjyuXnJAlmgKnSepjqugJ60yEs8Gi1h5L33+/o0LkalINHTh
BkcO7E28rWiaQPm/nuwSRSwC2zUZWAPYImhgVdm6Ps37GBJmsVx9cOkwkxnjgXRX
kr03+8pob0ALFFYug6b1C9S5FgIZtWnvdYOe+JweVDv139B4jyhWwI+BooRAbNrA
p8RPG4aK0nn90zDhhU+kjRXdw/uppripb5/YOxZbcFHzx6IMVvVACEjcc0AY0ZHu
mv2OD5cSrSMCOwVFr+F86UBL1zFUzLchr9+/NFteosqSrckC6e7+VU8iCjpa+L/A
SmqSti+aEE8AVjqsOVQDjJJdlK8XaPlHDlRi7Nyonvr5WaykB1qOfY36I1bkqBrR
z4E1BkGAF1usHQq3rzmP4AVLaqp8jkmsCyLUwgPzaMYyEPsC3zlhrhflvr94s4Mh
200rAcTdcqR4xYvo+aNqISrmK0zVlTzPmDSu705hnA4iNhGUNWyM9GZoEL6GzJss
Xy2kkLYg2eEIZa/bSx9eCARMff5KnNHSNBG7+wasVYkx9Iku4RzHMht+YmJsH9Ao
3TegNly1RRQ6nL1XC9wtKcei8/kYBuZLPBW0iGouIQln+R4ckETGRdDf7w4JVfQo
2YTfpitms8wwFiqbkNNeXnD6VcwYL2yJQVkttUCSOwmOvQHqvN5/ntp4sy4jaaBp
N4aEqDrZmXbwDT5lkZAdOcqrp3AtpAFiz5xDx5VskPKyRSt9eBFQMe9igNNtAGBy
IFmUlLv8HcmeUpXAAG9CuTpW5Znjgtzjq8j4pY0+fgsp08FrlRiuQoFC9QGP/pZK
esx91d8eldR6JE2eTyJu9LQ5F/SNYDYEbKj5KkrgV7AtBqzuGfqhVC7xahXT52OD
KmxMcT0qtLcR20r8H0lc+wNuNQo8XdT0+oR5be3S2RqcYqTMMaC+PqaI3/zRGpiR
OpgaPAAlMR5n+XgUpPyULA7s8J42U/E5X2Ytugq1861fiPiRjR6ufAdCucpHKrj6
1hTSjo/NxdIQH9GzvA1LzlDOsYFUjUZCKL7aj/TfFZf7kVoWmnEqcL2gsefY59mK
HnaEnMwHGJmwRCNVlsmWYj/ngb/XceoRlX29ExlHFt1vN1YStz1t/oZ9D0Qc9W8W
XOtQlP6GnzUvlLtP8ZHMYpvze18TX0shFagkKa66bmh2QUD2nA4jfkN8Htz+QHHT
coTazKx2WfOpNh2YgNxDonb4v10MrVylOFSnjU9LlIsCih1+3DCs6Z2gwQQ/mJAb
iqQqEqG9L6S962lSJ6SVGDSK/3X2sfURGmhvV6LPwNnAzXCUvhsA16irZNlyYwMP
lB9UcGiZ58MNVLtyYA/ODZn/P5sE4ydWPCHpe/JDpyo9OpKG1hhIeMLCTTYNviac
ToghiT1GyxRMV3SwjW6xhV0yAMkWEV/lPaWFjXnxfqCMb6gD/eZeEwP2MXaKdVhg
uvOSpMF2qCkNAPmaUHovWezUrHHbkKl2GFJO2jj1J28oyUgGwVgH1iU7XuxoJfHO
ZH5lS2oJ2xrNMQBCQPVw4XEfHqRkgiFy95Y744zahMAmNI6lvEDuUIqAC12GpMw+
tB0JTCHjgerb/xdT0efNxWwwPFgWZNEPG+qGMq+UmYs+QTPIzNk+y4NmpGk6uboe
y5T/lYzxCaO09BtLK3nZSwizzQdvzmRlTuV5aQSid3pa4h97VOWZ3tYnSfI2w1Fp
dOUqXwrBlmCtVkSMLUeoBVkjxt2pRwG+rmMjc97ZTA1HY24H6dUSaFr3JYhLz2xP
ZnAnOUeeZt1jWufneQq+LXSnyVTuP4w9k3/adq1OLDAu5nfkGBq4bMbvyZir+loQ
lca+pyRl/fxHQuaGA3oSJn+x8Q/oYlTQiZIfUNh627UziC4b2SzIBiJEY7830n3C
3p7GSvVrzur5R0A0TnTCyIqduxwS8BJHPMurQ3mRz3PeHFUC3GKaryXZftMhUviY
8Cx8xEP9fxg8gQUT8aUZJEx0Rlyh9k+nAvtGUQJExCIbQDrIqGZfFcN3K0M8pb+Q
pn94s6V9NZd2gCe1LrPObMh6uTkwI186ZFd/6sk1lCg6OA3lPgyLu9Cy6aqA0et0
AqSmnb0T7pe6/XO9end+GdFkjN0tCSZcPGbv2fB7Y96ykonCfiiIP1pk9v1WZK5b
2t7kHKdcgLyI5PPycSKneix0ObrVc+2jgLk4wlMF+qqULwovBbMrUhR8TAL9BiZS
OH08XOb1HNy9ndHB4hS11kMA3gk7D1NVl1N4U+kmch7tg7qQ/Fz9PLbN3Vgrqr7B
rMMPsom7xTMA9jDcnV325D7eDIbZJ4ekfTfQ2VvN/pEK85S3HgyTKcrsGEMNYnzK
537q14N2hu/TSX8vtt5djbyxE+Fzln4NzkSpnKxubf2SAv55PcuY2REKkBO6IgC7
e496UJij8CpxWCip+l98pFJdyQnIDoEAR5k6tZkDo0ghtAYpOBUhLVLLZhdeFtHg
44wPfdZWmGrHYtCCPEyT6jifxm9GybhXGsp6LWOpQhpFAyrgXsb9PlFQOqeq2F69
M8TaU3Do+oaw7qGvfH9GClvIskCh5bH2nYx2u4Hj7inoZEIUvSN3Tp2zLjyb2xyn
6ZI1dyRTVWwzsmA+wLtmO13SxEhYOTkP2WFmi+gabmBPKltt/rpqcGq6okufxX3W
r7MnKUJF/mbtdF9DM7xa0f2HmyJA/x5HyUCnR5CCk/WG/n5DDlpcP+mrPOUS8jGc
I5q+3wiaI5MOunFmP3o9rqTs0PeQ2+oyMvTTeJ2tbQbRsLxWHQ1q752qpTfmO9T2
zVRWw399P+bkCnjaJKQ4Xy1xK6Vu3bCxLI+mc+gZiFtRPyxF1orxnNApgaGC16rJ
sdEW0BrzMUD+cSm+BMzl9ij9oxjFh4lTV+PuYEnZrjpQAnVKv8CkueK2vQmzz55B
RroMSiQLQplyDt7vBOkDr22IegLEJbHPtHsj7oThIVXtGhoy83thvyqSKm17mHI+
SP3e+TPgL5zzakPL8QxjUgf32wqdA8C+jygDwDegpIffzNyUuw0g1ldHB+o7MsxO
mp9ok86mHEHerHw4A/2qChoPSaBmYo+r3NhIRGZsFUQCteyffOK6lU7Xg7/Qq8dY
/UInXo1xBtZ73hUIC4ew7MsPNZvZWjVqCSePETtsmqIO8UVQvMGtPWcB6hub7AnC
nmTJfOIgIzEarPFT2Wqj3Ox2nbOsATXRbW638uMa8xejvxdYEVJHxzKWPfwHfkPT
Uv3huTNOx6sGVTN2H1184nkvt3Xyg02EReN/Apeh8cslDBfM7nbEYkG4w5Grk+Y7
2yM+jqATLGWy4X/YWjBBm6lHnVvFq4rgYxoAdN7C5ezdOl5dkzxvodvH6Bloz1mt
VlhM0pQmMDHIOuvlKd5mhF8dXbs3MxRkpQbsdNqxsdffqYx+IuducL5Csuz8jIR1
T/c9YHjuN/+YQEf7Cvp7BE88s7DJ9IwyKEJ4ox1vMfd4Of7aMcWFl8TyYPviqabL
5UQ3RVhaoMCEAbEhZBX6CyS6CyZ+Gp9+xShGDSi0GDjSHWPuxONNV2UvBmURrjpR
BtWnQ9pjiBx3tnjZgcZYrnPRMsWC2D3J7RX0go1inSops7pZMwtRfRQLZYa5MDYC
NXBesvPjIfNNyxJlyJdW2Wk1xg5QUx5J5JNnlKDuNYqzCMUR/TENeVwizspc8YE5
vStSSaxTVC7K0Ned1uR2SQlv2t1ZCq5Lx83wybPAG+mKU4qRJ+G+hFb+0yVoSc/8
62NCYF1WDJHXJawyiGoryaDvAewPgNdSFuICQ5UsF0xGkFlJUYZD+p8ghz3ceayn
5l6jw31ix/vqW0huHVg4evIZsfiXmSN6Zs55vgPJ9HVPCf1Gq1D0NC1dBRYif+Rd
FRR2sBwLjTWfwy9mJonV/iLjW2cCVLBVlNlKa2xE5MYkS1YEMXZdW7wTadE3pUjt
rLUpYMQCTVDm0m1WqFycht3C+1mzwg+OzTt97d+feV7FdeosjIDQTPITTXByUnMg
uz0ZEWUWAK0usZrqk73QsZrQ4q//Z9ORO6WfO10c/A+neO3yAcFVMXSu9tD0fY1V
rUOJDqdwDNpTVUPIm6kz1h9P0nW4QpnNVXRNtRE6s7r7KlDx4/5sn4jgIcAN8tio
YppEmh+2PVzfo3gIfxsB7wvnYJYfaj06NFwFajJPvt7mA9DNpyJkWuO8lJP+bMzW
hSOzKx3zpYGdiPor0FQMN8Fu+DWB5hoEB9l6EqMD9WTVbU89ItQRiXLcI/xARDJL
2gizbfAMqiglYyNxQcQEAF3c8SmNCwffzOLVBU9hk+Vk2k+wdOoMmNlBf3w/PT3p
C839d0yoSAOT/iPK8tOcEH1gXb1T5EdwtMg0BNQPkSpaAUEEduIIzSKIPVu7oBc4
ga7sJSqidCdpGhcScms4okcMK/q1oCRfFTnFv3zzzol6d/gorJl6reaM8HNW3Rrg
mEiO3twnJ+4CabRqIZoDY4bbTc0uko8ibcMDlB2vycYr6dS2JzEw+O+t4CbDhcfa
rjua4AiKWuDMhGEz9oFnPhGk07SWu06VEyVNWbymQjSHUCogNejiGdpveVhbLexW
jVQIfPcoVSzmGMmE6qc1n+IhfeeEiR7/7XAgEElJR5ya6Dp/V0QdySXPXdxB5PsO
qa/07bc+Gaqay4CmGvCb9TTk9FYhUoepRTipz/cj08BfYIiilLTas5ZPryedEfh4
IGUTo3m/mFCzMHgm3yIiTZrHv64emOZm8ELNgSKyXzDXx/oJDlxK3WBPbZ4S9WHL
aIjHEtn8SqzPmTaz0uCw0raFeDXFXmtC791c4FabwghUu+/60V0YUKikbEJw4Gd5
EWIHJlDhWhauUIW+HEgKe8Cs5Kk89aWyNV7eiATtwIqV4FxauGhOvb7JHAcsKlzg
kUCG3JKxck3wYTx+xI1EqvatYI4M/H9wWRo6jirTxv4heRSczGA1E8hEtFrhHlm/
ni/uvXHVO4B3de8p2oNTOry3YQqpXUDhau47ltuXNmlw2Sti99Xx7i81ISW092uh
HZqqbZv1ypnMu7eRURAsSglLBocYxVZ4n86DFIH6HQYRsryRl0oc42v+s/n/lSP4
DyqMVlVEwRm4fqF8lhEDPAKGAIayNdSduUm2l3qHDIlbvtiChmBNfIA1jR0MhrXc
BHZGUu9xr9toKgj3F0WFghae36DWDv3Wb9eGE+PTX/v6AWyDUu6tYrd0ZBdZKK50
w28yxhwmpRFelphh07Xu/lKKSbOkpWOVf2Hj4exiT45Snq7z2ixyWXiPdG2XY1sA
VW/vsUpq6aw07dGccWqv8CEto34xpIAc0BBdHBYmpuUkQs4WcCb/8i9beq8SVFy4
seRxdl5td15fByLKEtAtWk2RiX2YX/DDCS/k/WwUIZvWBeoXZUi4eXx/pIKY/sFA
YBSd/gvTI49+trmVyEQTBuYqxL0Ak6HMGTnUMelXMxtAGVBi13/diBleKIos2F9x
dGuHpug6e1iHX1l2k5ll0wZoYgoL6gSc5EG8SP5wOUCLSZV+wPheVYL1iVon7qt9
ShbkuLMOTRxBuJae8DKJC1xGOjgz1G5iZWE7NuSt1QruANO+lkPtI6fUtvw84K7R
PcLnzq+2SLtW4dXyJrsTL5T0hlYrch6LGFbYXmlWxMlujPTp94ll8q5H45AoHmpz
ylyu8rTy4kD1N5aQ3QKxgZvp78kxjyx0QOGBkYG1c0n2pxmsnahKwy3rOgJxCeEs
+Hm8uUNCReHggHZYpQS/8JFBfc2jV+7ygoPdcqhMyqyZ5fKYXXbKs9sxzuEyF8Oz
DfvPT8x/91F9XL2/nwV6S73OPMOz0941YsJYWdePG4840DIzTKF3buErpDWOrO0j
GTIck44JtvRYMdGBdSTJfpjKA5tPvi7n008oxVxvkYhmgpXBLMMaGXFcew6ynFUE
7rkYX1g231bCxscJyD926KU12xQBH+XmAaj5gSAzrmqNZ1hpsF+5HP9dEH687Mvb
5dwVDj/bmnwSl4N1OPDv2iJkgMWmqSjFJV/0DIs34GrZ9XQW64AJPdsDymbc9+5c
zjOeDePa0v4kU5eJAke3pFSq+dq78GtfHwzgzEpDHvmjd7Rh9cETMAsjU3Ulqcm1
e9Rgr8NBPi9ylvq9XdUa5/cprUkvU/KlL4J+HaamqvkuikvniG2n/ZhQJyA1kt+w
HMhoeaxSDuvKEssfvdVnMquAM8GkHtq5gQ8CvzRcCxLoSwiLrP0hfm2zMRizJbTJ
aVPOxe6ZVKludXJ1KjKYXnwflSFbQruUPufRRTV8WC6laay7zjMaAtgd34rU12rq
sJHeZfusv+jel0n6nAhIFI02GRKfxnc9S8Z7nkNs923aRdrFtxr3k5JPfGYf595z
4i5fUc3k90pOG8EsmBZeXUP0xznJm+nyQWxYSlkuhtOSUAwsuwXJLF8emCD8kVql
5eTItENFsKLZLYK0/K3ppYnUmuXIczvTjWa1DZ8NIqSPpytSyzaRQrVttEjyQ9pV
5LBdPf7H5GVa2yJ0qYPTrv+F5N+t1i0F8XqvhCPXPMGcTAZbUr4AljnsCJzpH6C1
6eDKp9VQV5p5kHgTNRsL9n6TaUqw4sMHpZslUwlmrqwPsdVBEk7IfE0LkKwxtvhd
j9Yj9C6p61efAVGiQFtUDRf4dGJJTtUwBK59aEyubP40bjp0ntgkLGX5slQLCL/U
+FMcO4YiCGquaAGRzO9iSo+bXxT7guzKASSDZT07Q0E/O8G+9734QxhW0Oo2kmNM
wrA6xK4Z9R7xArh77A2pgQxz91uToPcbifx5OhcL/qpbWuW7PP9UaJ2DeKcg7Up5
3bok2ZzOm3VZbTzRCCRKd6cb1V8RUVdVzeze3st5GW+9v4chor9G8JWXkV81BuUk
hWWoKg9Vvn/RU7uDI641H0DlOSnmipdJADDE+3XfKn5pRqdurWos76IiqjawPlZ0
nXJh8Cxu1Pfy9Z8UEqlhHHq1bfVP2hgVFYRnHbTsWNCLO5o8IzPqLPO6M3nf8ysy
gaSSL49q8R+m7jzphj4cUUwNberrIPD+mDXLAGA73f1gB1v8OZR+cYZASYPVkFXN
6mit1xHvUdnWuvbJmwQKJ0mG1wo0MGl1hG6Yug5mwc9/T7vpATP1W6cU6CBmLoEU
gz27e8rcHh0Rp0i+Q4qAAS34dopi/IpOcFqkCVTIZX/igIE/am3lhfmEeOLFcAvz
BgFPgOtR4dsNRFgP5VCenfFspt8z7eRpvhy2TN/aDbELpyYRoSMpb/EMsBlM8QAg
H4b/cV6/Jft26bp0voMx5jum07d0Rq/sfZgo00cr6gGSACtx8nFggrRKrbtewge/
ZfDPNLbrs0ykRv6r3znrTAcwl54ttEz7ffO/mFOcfMfnLRAIJ+u5aGRnWg0aqm6a
+R7EZlSWQkghuCFTUTrKjngfmaRmRGXEIC24ajH/XXRTUJJh/mhnHd6S/74/HHyU
Be396lV9VkU4ODT2EX+PUUvEhyJsZDtGF24j0KiLCTbRn5hCCrq9PL6f7+BN20z9
Or3pSZHuZ540rZkY1lg+PBIyDoqA/Su6yq0E+dqkHz9ODyGaZ9chRVbaCEfCzccp
1WCAaYd9/mCDy4H5Knqv7BKGq2i9iLaZDeWQiLWayr36L7Hx6iZi/h8rYzJ7W5D4
m5YRhNmetyO1d6SktMcT2zQj8x8utOXSFj/goPWZwu4O2RosTvM6t7AjARhOagAV
4Fcu0ythOMP2R3VuqZsbk7XvsD/aevQiZxoSYPxmeUJJEFey3XrzbuDsfrABsQoI
Mk2FwwFJZZ0H9xUIQbXh8fuVW1JTDaNvw/Mbd+56TdLSXvrP1RagqWyRiRwD1i/p
Na0vWc+ouLgaQuJRx4c1UgvQm1Dg4wwaTmr3CmVJast3Tadjp2LM+lmdgxB6v+Yh
tBoFc4nFZ42Nj+2k6EBdidY1s9NDj/O04Vl4b0rdTtM9WO8OGuG5NTCHu0xIMRpA
pZwthEDRlEjJx8RZ4PsXe+/eky0G+Fnu1tcthpfXkxXETuOy6RTElTQD7hEu4OWh
GLj8ba1Q4UPlan6JzhOIcVWspzb5rTxgmiqeFk9Bp5RY61TNjySTx4Hnav9TBtDI
KOeH6yNoKhjGGyXPVFEWIaTLS3uzK52LEzqCWDA987yd9JE4Nz5vDhvr+ufBpVgY
b0pRHpmoO49wc2L16biWQVXLx030Fv9WP7RGI1gZ+sOy/+y7XQjAtAQgOH3uTzEH
dNeR7SCxo/7BYV3I5jQs+UhuuvOH8ZtBR1YlVU/cyEgo3NmZ9MxRY6MiiMlyRXhg
B/Yc9dLpuRyQeoZ/G8VH2sPCkKL09rZ9Uu9MyIk499qByUZ+j3CoiGzZsWENK9jv
jzFdzjW4+GhVQRzluFWym+WhHvb8pUnUX/qVplxtgG5Nvy+yaBceMOLYV4Hzu1B2
Tn0IlSCeqUTWTCeyQ9s0ZOxl8nNu1u29Uy9D7JXUR7EXb5J91FF2YPacyMh1tP7f
zibAz6AnuK1KAunDxh/2f1amIgWvmZ1HeVFuhdZpHhGMzIE6c6V1dyyHIqKLnxRW
J7nB3Eqkia/rTQAl2Uc9MsEDaR3+vsny8pTZWzA3CuWN5p32uX07JMfKhid1KFVh
K0kILgC+nC+p/7ZD8L2kFj1u1djXVkG3cJlh7FLHeUmEkEljMzFoOlp2pZv+I+hU
iQSEFJErJRhkNf6cGprWVlfRC2j5mfDn1/MEsnM8wJx23z72wb99PB+JmFVMqU61
ULMhjwjZuXIO2epRCoOq2cup4zPT9ni9MmIVPZQvT7D1AFKrgmsKPVf46QpGPg6s
kbUrCedjPLDX0/0SbX3mStFrBjvQ7GrWqh8RlqvXjhnGPp+tAA7AL8cDQZ2W1yRv
5ZSrUH+LQV98ZiwsALDgmEghlozGDhhqRqiMg++FCIn3skFuHXPYxcRoTVHpuyHU
rVG5PWgMVeTCX/oKuoZvLl8joV5xdZWxW7pgAHwSC3MG5MUzVDoGW/YWjVlGsLMF
o/Y3IRBrDlTHVjeVAhG3TpR9TUHwpCVcmtCweZVdqtPlFzAy1oMGDdA3VbPQb5Kg
Ob4phRhKE1Qiih77bic4vRQiSifIOj8ameJYkFUttvatTOfSWSXb4sE669FHjNfR
EPmcar612vvg4ajAGI21lLbPaGvJlWGnF+GMGpLgflue9t5xeVp2aepkEGqRafXm
iRjyApAAQtVKq1T20PBifOgKLMRjHVQiaiQM4oOgIJ7E36p4YncK/QGUs3lgWepQ
kXuOTJURf/TN/RSbe4496bI9zGCdGFEToI/8yZnWJL7fiAWACaJR8PwZokvHp/2B
uZqQhBmdnWyMhtGKBFP4pt4JwSmZrMK4SCRRvKsLNw/4Gh81E2XpFmbFUOsP9yBx
u9+oyK4SeNGQ3WU1M+KC6R3YlPpPSHvoL3bDv2vs7gBfrYx4I129/fN3B1NPfEt7
0oaOTzcIObV2eByqH1TRIC8f6FRDhOX8RY0qJ3AxOWN6H/o8sXuaKnWDFk9N5vEt
iAaA/rirwHoXmV5QKun010vYKPE773n/Eb1RJCW5fWEdcp//PZaJMhmB2D/GVNIW
6UXkT7nY7BtxNo2s/1EnR0FWd79a+D/zoSuavWnGBSHnzyygrD1il+WCFJWjV9KB
wGUsO15Ub0cCnIrPrlG2jMQhqfy/GsCMJ9TDXHnwC9SThMDgpi4TcRi6TCwaikxh
fJ5rL2f6h2DnWel0bJnLoZ8eMS9MqpYTwfuXlE8/PoS1Cp/HCrfbh1bFsMXWwDux
JrkdpimU3BGyJaOVl1hspjxvsISIeFko2ilV6tjrKsczoCj6BNB5F2TyKHlIu6vz
VIFbvOtcSBoAYQbPvOwRZKC/BFK235XQs+EtZ6Ehw9Kd8IJYDSvLHHBIzWN1hpyV
1o9aBPbqvkLY0p5Z4etkNbht95QofKxE2Fe39vl8zl7lVHukLO6G5Yc5waenF/iz
z6ygl8f/tESrjL5ZM15e+d8TLkpGI4ti3GlZjDl4tuqmJBgEuQw2Arwz/Cv0zvvW
4fBTeTMMDmYW5EoiRZbymwByrktEVTWuKQTEGFtft9jnummQmGtZWgos72Nib9YG
ZniSB3U+Z1yD7I30pMVTPON8ennP1vQFwxhP6goX6dA2U55/891vqjftFYYffh1B
yVgpPbdQ2ZEaySW0aVP0LjYsC6wYRi50OLHONkCxRGuduxliOSk/EBOs7KLlT0yn
l/yrnpWmMcBAHNtupQlCjKhkzU3x2fCIOquvQG7dRFrhJGUPtDppe3IeAFNrsFwC
5Z02edXosSWqoEan7VKUCWPYo93i5fIPFkZ2fm01DaLXejBCy/GvMzvSFx+OSKie
JyoaJ4MnezdI1n+Ji71mEYtDWadyXgf+Nm6DQP8qsbwRuCSV/8MRfQZL71MM0ppd
fTAclQXrsYXeENTq4zDDjS4VCFi9E0VW1bqrltZUebTWUeAg4OQu6W7jZ1eOuh/L
KwGocz3/7tUwGcohO0cBp+j7LF7ZwYSHju+BeU7AATISXH9nBqHuaAGkBvKPMlsZ
PKCx0J6XXqEBqMrgCkp7KNR+gH9KnTYJ2/aLpZ5CgyZ36XTccWHtN3/WTWyb5DMg
38GrhtqzDoMcJFplRFx0y0BqUPX7x6RN5YmHvINXhUBQE/VAehcFy3dkn/PJ8b5E
NJc5aYcbvf+ng/erg/x5Kpt6P0iWJ0tCtuHMvGpiJqAtOjmg/8vc6Wvu0VX101BD
KaeVVDkhDrHKQexIFvi/jnSK4vsZVA5ZNBZiqCXuq5ZsaedTGjlI4gsYN6V+YFCH
57aHoobHWsIVs7FfboNpXv6r/cVD2VbL0xYQIGnzq+LvwaelbZcQG9tqDXROVsw1
/zezXtIsBxL3CXEBBs6IciywAkwfFV8UjgHW5/0Vz5jTpluMNClHx1a+OjLI6YCk
YrpKw6PkZZOSmkLm0qqz69YIGH7/Pt8ZtsLwgDQSW7udwPUXF/3ZVm4RXo6Kc2DZ
ofiV7L+eufmovCznUqBVzIOHXP1sCIcjpXxqSCH3YW2djwf/EOxDy7Fn1MZbg3z2
L0HjA8tQ76G4M1vQ9c6A9JRCpuwJcmFD7YixSjCuIXMXXrzHQRdzmmE+y0nIXfFm
LsuiKnvytFqoG44HmU6lnIrBSIuy6SzFc1xjupQJeKrNhk7jFO6yz+mtxA+w/NwO
eBWV66Uc68O+udGah8m6j9xHDgFNR47m7BYH5Df/IQ9llQzqpfHa8HyZATmYKv2o
qiqpEwd3iWbJnErqS6lytvr3/9gNVx5Ohmv05XHhwfSMPOToj+4QhLPhHQwskB2B
VG991xzH1zX+Km/SWE6hUecgnu7WgC+2nVG3Z1Erk6EEhkneuYs96Y+tl0gbCUtt
nE33rRm0pTlZzYfy+XrPBsWay+lvZdnWqproK+GoJMQzJeAYJErP5II+SXfk07kI
FC/412B1nz1+bAnzi1YDsotoRNEAaXKnSm0p/QLr/8yV/zAV3Q0PbymoZB+lrQSL
tPhCsNJg3Zr9GSwB977bNFRYO1Jul3h5QyQR1Ig1oM6PLdkpkZJLiRwUBcRlenEF
y8ifudaXmUK/jBFAzY6SlAInR+RByWv2m+Ro+4WFdIZcvHlw/h7znVwMsICHiIjA
EqWk+6Q6pSAjH1vlD2olmifuJUN9ahPtqUZWKUlxNWK6RZbcIBe0TxBRsG6Na8Kc
p9Nxu33PuMuh6QAOIjZKSHB6caYH3/n5SQDI1CSrRWuCp6O2MDHdKgRWQynyjXcs
7Zv0Tkznb/xiRmj3NWSqoZIVzv3gn0okOn+g+e+8Z6pGLqHE6YMwAbU01pojttJx
a78mNhJ4/nSbveRGd/UbDr5t0X3bGhDJMq1D6IQEJq8mIHVh8XzCxkfK77dQq7SS
Y+YBTqtI08ycX1munIHWMxPucGQz0YBhw8UgAp94jkwKDPK4cZ6oO6yZtMDhX3uQ
XmR/G6RwFXcnBOIcZ7Dc+NdzU7HzSt8J1rXWN3MLXxwW2rAVgmrJvWd2bkvj43n4
wDv6cihuTJ0SmWf3vA61Il4/c1U/tGWf2Upek5p2cFiXsU2+dDDr+jaMd28OGict
tba2S5bWHQ3lnYgPT7kLTIyv4W+PbQxyXzWPkH0NimfBZNGiya7YJ7BVZIk8LJMr
sAVxFZxNklX7ocQDzem166c5Rko6wquQ748rM1KYGwsVo1rsbx6kIAWVe2hdKpRo
JYLbHut0FSymImrD4v9MBRx1Cw8Sp+CGDN1MZbqby49yN+AVt7352hDZ9gm/cFr7
tYU6uf1lQ2jCnK2vyzQ1kksD0hTVumMGkCsZ4uYekvGPZXQ+dsupNr47FidLfD5O
fKnZ+CUfrcgRFfIJYxoZYTRCQQNk4tR5CjIQI0eCgwhgdXTzZbl5llhaBD8Zp8S4
zU8yiEr+O/fH5YmpjMjDSmjNDB+NAhKBp2G0TCVNCCZGIm0Th36C8BPR7xyGRgcn
JC9NkJxKs6vYG/oiRt6EQQ+/LEWgOmVv4TnJ2l+RpObJ9S5cDgTF82KioX3FA5L8
WVKhhsKWViDTZ66BtgBifXdAl9CrNUl0vkmXePnTDtVh46qoIAvP/jilS3m4LJ8R
fJkq5enVx7glp55b7G9S+W9LFggVJm3d+qXgKw/s/AMVpc3oovA7dM31AVcu6fqR
xDKkZsWvVjl8zqYAtA5eIoLEk39ShYZkCOf89uzeHOZVDacGgdC69MImpzDAIH97
vZuM40uu6oBoX+rpeiGb3uoIhmPZZKdBSOdlj0A3JkwBLvGQu3AyahiYkAUTU5g6
w5zFbZtvz7tmbsACFDa7WtNQwTkNLiBeGhMSE+43cERjFwtpI/23NPuv4bzmq6Wz
6Rr+6wo4EdF6/PaOAlM5RGMg6Jy94zrkXg7wdIf9YzGLyd8AzRPJjwAhcTG2ZH+t
1GtvRrtuFhiBVjs5jpAKPgBqfprxvXrNCPVc0YYZcuJHsb91fxJzopa5GOXlD0Ul
u3r2PLMDfsdkC2STF/japganSbgAj7dZDN4Iyx+Q7z1zibmYg1iuXH9JWLV5gKTd
dQaxwZKe6NZrBY26fg8iXsc5JX4Y4AyLfmcCOH7XLuRAhIkCww4kqY/jVvo9oa9S
55q8OSuLy79FuyMQzZxpAXBD5I5CB6syvpx5WUiH7o9nrmIvBNH+BmAmqrocl2Pj
DUBwEtXy+GpzzIwAQikv2/ihwUGMUH3n9K6vQrpjJoX2JDTosyD6TCzjzGOC+Dh6
eAyCGoiF1Bjsf+fJBaKL81zs4CgKCPdmutJ9Bm5sn7fcNEEQdzk9NFiJ5PclYB0D
Hf8YGtT9GRgULRq5O5QrpqALXB71QHGgqmtp5G7b82DBRWPTZ5gKmxlgeUoqaNvw
cgU13H3ovSS4tu9AL7sJfmMWem1B2LuWbgIY1VdmE2hkNL8N5CK40nXJi8aUY88L
1S+eFZE45gIRJOrVQsugrDe0yAG020K4zG8V8mAB/urmcpB7F7JOv1S419iZA1DF
pNL2lzc2HH21j4c3z3JDp2/VmukjCcRDYEBeQhoiuthJAGs2hy5zAjGwlfcL8yzM
KDs4iyke9L0iDQMVFa7DYgeyyE84YfliZG0TKdqyP3lOBIYL2uBXGD3lHhn/XPh3
09J8aI1W9cXygke4VeCBsIZ2v0CFZvx0ENgunleJlGNbBDyrBWKWkpcpKzHXybYu
Wff3l4CsJGj6eaDw7Ftm8sHPpIrCh61a4o/IpD/MU9+rHrv/uAgYL4qDEMYDFFgk
XnaUAGPbgtlaC/2mNLsoWGbOao6HHu5gWCOjYkmJPBM/hlul/EbGZQsyneYcV1f8
o/9NLrM82WAb3Y7Qd0pOx/nxnZG2Z9vpe+9T879tN9NmyX5syIIGjBFC6drpR392
dE3R8DdhAYJS8pNbBmaY5QLTB1i5MaCzF9R05m0KB6Uw/b/WB1DQjmwxAKsJCn3A
w/m53jUD20ZlBzpAjIEqSTWeg1Ra8ICD+EXItqlVl/8WCKhw+hPAGcR8TKYvMqtw
UYSJ9fBgj3OR29xOS3F9AEizlgBivPRwgWB8nPgPHULHz9JtM2VELl5JEKzviPPg
JKceYEYSiZiEKjR4HAnMmd3wqxU0yfgSJuphERBhpDEWrwOICClrf7P+7SK/Q7rB
mQGf1NZprJuFPOrm9BEmrmChKcnQ8li6D6azxyc7Pv2ryITKux8ASRTgYXG+vbVG
SYW4/yPpVXzJevpS+fVMBSQujiz+YwZEb+ubr1O0xG8GVIs/VU+RIdoAYOqmJEyt
RMVslbjSlwuuRQPmDXgv3W8YXWiVVwRa6CkIoQMqrzQIUEkOEUIVVPExjrcQhPMa
jvE2rm4YGY28L8xNyRsgabcq8QgBMH/lwuNxN4IsJWFcSvGJSLX1eEvChcQdb6VO
DIrMPC0oWz7rvuUpQD+wwe2QN7GryjNjMnFJR9Tr8zc6mGFQJbVssAQe9irlbDsS
fHtGWl3i1IOQxxD6n/wuBCdX/mP+pZKyyB/mm5duZeQrwFChBIOWbMqYsDOcNTDp
otYqfrVpNi59aOIJDkl2fMD+Ahla3oGi2B2AfIFvEwx5H4He1m7qweE02PP6L1gw
kYZX2XJjZw3/jjToOclbiuZb94i2Zx9onjbzOGtLsAM8msJdChrsmaNT5g2u91dd
nEfZpRVq317a8EG8RGel346aPEYl6xsdHcFcSYUL2qpGwn4QFjN9VUmj/1Nbm9Pn
Zv2upn2ijWOV7IVolCSJMhISpxsWcleiFyxBHui47PJsv2vQgweUmyQwAiOEfKJO
fdQOmEmaRSor2RsXv5QYoPR8/HXF7oi6oohiXYtohbsySZlGbzKapwzVmQwqisvK
FZ7b2XF6KRNNT22O40bXnXRnz4o0sP+IdpnQlybPrucnD1d+N5Y8HvHuKyvSvA31
nAX/DVEN7ulfx6yPIz8BA1LvxxiJ2oSIi3mLjjVGWBtABvpbLSvOctydO4l2Ic7b
AiMLwOxEQIaEzTPD5Wjv+fFuqSaWoPh3chwKk075OGXwcJvwLKIUTwH/3jvu+Yj5
mpBOsP4h050UCqpzc9J+NgWerCDUiVMviodd78uqZ5PGwJsy+nN+WJL9dg8R+Asr
I5GDBB/DUfkFKWE8Fm0+9X/lMtsj8bHMGD9MGwJEUWvTf2mQlHJlLrbXENvivzSE
f1ab4H/TcrronMEwEH3PztbjnzOWV/JOp6T5GTQxS/UNK1qr/grtxBW4iLTtRx7R
8FVlE/k/OoX6JvV99KVIi40/igvbrkxW2VCBD0TfA/AiBT4pRTHLIQL2fCwpftEL
tiG3jSlqBOXCulyyM/Os0oE6SvfV6+ZL2Uynv+gg5oTaH87zNapfYVR/a/uSmbPr
uib34CZzePSlLtTLdi6u0LTisZCyGP/cEtmzDRIzmdiNxf6UZWqkbPJF1uc87r+t
r3soGwpja2gBE6zpZxIAxmQ52X3hY7jjcP++MsP5wziTeEh+e4BCImt0ygq45EFl
4Fu1jgmqENmYZ1tNNqyRTPQbh+vnQZRHK1FiYUINsx88mpZ0JN5fp2lBev8YPBa6
D779i8R0KdZnE8n2x4w+hIBAo4aMKD1WUKZb89iFrfqvkAQQiHzMw/tdqQ0IlyqS
FsB3+1MuWmPE/Sw3ux6f+aFIbwYTF26F3clLikX1VlUzL7fSMCCqwps8hYt50hUe
pvvc3Hfk+kEZM7MzY67fSE4HJCNOCZ2adfGISQWGu11JmAZ+NAYplIPMXYNOv0Il
SlUwb+WroZXH0kwB4hx6mudLuY84rrSLu/cKeYM+ybcblcEnj2OHjyc9PWefOhgX
W3P3biFs0Ecuwo64dLpRUByS+jD162m09I9JgsI0c0omzfRRQgG4tePHg9szD3PB
hE9DrHGntAJ4NnoIWNQoEuwhVHwzTi9ONjtWQgAuBIgSkSQ6y8BzgNR12ZbIfWaM
rkfhfOxftTRlH7Sh8gzNcYqBkIidUzqsiTtaykB0CmcZxbNFF7vm/QJqHUJj105s
TSOZC1+kCyrn2m5g3XqoeYwWFfOvcAjpFJrlAHWBCSvZmi88Cf9WReQhfa+PNztn
a45Ud7vjJUVd2ZAsuom/4CLumcIBooHfX8bcG01amlHXN++jvnlLq6EV6eVgUllo
xV62J6bwMA5GfwIoxQbQ1BZfMo4dHngyUOMCia5juytOUdgqwZENBEYyIwEWWGF5
d1sJD9DeZi5f7onzwyEn1v31JBGW/4j7iEuTkrLBHT4Qn9+fkYpmf4TaIiWT0UDw
7EiugpkhnCQssT0bFSUuU40KDyMr68HyPol7ProNY+PDUjZwrouHklERsKPPL7YQ
wtamUV47kB2BPwoLSA3YEhd8WwSqCV7KU9TVTwtsgVpb0Wk40W1szX6YwKaF0uDf
9A8c1atvVF8cLKTacBPruRKsnkRepiVYJ7d9t3+OF6CBQgExS1CdU1uRhY5LUBLr
+k5Atsf1v5FaNm/dc3r6rSreHsS2n5rFLzFvGjNdl09QOpj9HJsjOYMyWWLROga4
fcVMnjx9/jacayynNVansP5UGYFnti5DqbiW35BIVxoqWaRZZmVmph1MvXAWQk61
xWMsTpMef8DS4M9yV2LznvQS0v7C5F5U33RITeEV7cDAUxdUNJ48tSsa3SjTsPKF
JXm1d0I6VD3oyXsJTKxFG9Txu6H3jLDalD2Achc3SxWtvHljfpMoxl+vQE3xyJfN
JPHEdqLjk74nnkAMWnFTiua6JOMfn+PFaEV45bZ9TixiWCR9TaaHsYAn1lPNdfeK
ehkfN6/CBm3ZPhsc5mQWkCFvlx03PqC5S2R8jppZjl1uAtu7bp28MZHuwWjiAiOg
MVB/DTPWgLSWpQZk/UOAUAeiHT+ANYTxF70EjbU3QOYqc6D3P8HnJB9TKPHKVmt/
ucQTfnzeYBowycURd9jng5HT2LqHp5LtFgkPTDWuzA1ozN8RCMOt2NiVM+3FWWX4
3Op857PrJhuYc+scfBTJsN8TW6yv54hN5CB7oz+9x5ldv8IdAjxDo79cMmMdaEDL
N24hJxnmPrMGfhCRX8lAB4ET1toYEZxxrruLTY3fXiX+LnbzvYXI+/E1DBehf/L5
tCwETCe2jKEsj+NDrRWyGkCf7rMo0SW8jPW6Gn54udfpXQ2/hBqyzp1JVetrzHgB
S5SGzjUBdHrzYOEzD//LS6I1pmKUYDBffNtvCfV7gDOA1QCs4M2He5wenmmPyd5O
xvQK70CzJ82mDMaNafSkSLzfmndcHcHwi56oJnQkMgRXcaIuGPG+KOayZn9ch/s3
GS41T/Qp6yw9TsfA0uI9FvUIT9XoWAldzv35tZFbfp5TRabkS5sP3sBFh8iAi8U8
KBBUVQe3KGHfNTXQ/Rdq7VpurRn1OYNPIXQHyTJPy65zrs5pABzGAEsSs5V0bwVL
4rdICYlmggakvmAg1q3ZH6kUg1Q3jjrq4JlBE+JVubPhsQBiWU7FRXmbEuhdi8yS
4w3LdbafpX9XCCOchjqSEktt8HGRgzc5jYZyC7psa5EUSJ/JrIwdRY9ba9lmopEp
/KC1Pa+vtZJwp33drzIDjA1yURdXbUUyA12wZJu7WgOTsMQvjsKUBeZr/T+7wQXe
v62k3dvAbsLa+LH8SzAY9ppXjd4OKIM9SI+rXrV9EqizhUsUtFPD1lT7zfcFpxag
eO3DGH2o6Mr4lcd9tY7cED8Z0bqrSZR+WHZ9v9NxyZmx9WM/nTgcrBJ3noy50LxB
H/61uS9MzO7HhnWxB2s404qujPqvGB1hOWvgGmP1+o917AwjfvLpC7wn3XcFZv+4
6JciuuECIVqBrB1gjFMymrkCOunW9WCwsEF3ZgLhu76eKUw5077Stf9OC9xnqjJI
jd/fTj4byWiAFOgsImexNiRICiZBvtmKwy81TtTj8Pd7dPMi+BMpUU8vUN4Bkxkz
BZB+i2ikyMuX6An2KppCJak/Dt1VSNZ/OMUlH9fC3kZhS48N0P/CW03SnawI1SxF
gZcf2PAMvcXh1zUr9ZKYduYxb6+BbMBIC1ojcbvgmOP44SC7ZSbjKX7HFyN9zA5M
xcg5Kp+8Z7XG3DKkKhURw0X/aEJ74nOcrLsXKvzC6UuvekE5K0EicGK15kSaZLcF
TCVG3EBWF9dbmyyuBEet4BajQjUKm5nTuEXo5gmBss6/6LXJXE7dWVIbxXOHpW5M
u7h7IdeE8QS2biegaRS43PEwjjTtFMx+O1EVkeWTefJemn7kLGIwP/OrMTAzifcl
R3Zzyax4+FWBMyqlqtc2CZCGvHyRYp5clg4uEGnZhoj9pZ9RLJo2rn4DT1etiyMh
t48PebgqibmYJXmodvYM2p+ECc0C9qheVLvo1EXgRAxg7Pzkv+aW3NWnXcL5Tu0Z
A1RQlrkEYgQMjDUIz9yaoZAPUWt7Q2WYB1pTFKinD/MVCEFYGVuLTui6QEXp18ry
SBx1sBhex2JCNoeLi67FdjxVNN1KM65xVpKRRxXwWA1df/nMHXLPKMPPfOp2kbrL
pjnJa6f7b8+6Pw5C+FTUYiyHf0ZrlEixhfTGMLTP1zzIN+fvFj5Xa/qrybnw7giw
HQAyCHPKhfsYqE1VwJHSQuF+B4ROfJMB6mfX44UIQtVGeRJJCRq2GzT1sOFUBnXi
LjSR/JdZHYrXMnbzHKew2Q4Lobv2irH1EvETGwgpFRr3obDLKOdPjHArZH0nHrVk
kUjTEYaCTjmYzgxmRSjtZQ1hkkv1DvcwtP1hHBXobv5ayAVvb9sACHRqrhVYLhFC
A8Ip7YBHYrxp/2IRbIfsvAWCKA2ypZVVwklbRnyXeOHRONNQJEhjaErBVjhnSlka
f0p05ffXrqaldRRuBNSjdeWmUd331YrkebMPOixn6v+BZcNdS/HztxYPvwH4wELD
pGlShfW+jt3t86Lzagu3ZotULtKFm+hyi6iRliGrghFQDBcjJd62F/jl68ONEngo
mGJYECq3ZLPQpGg70scSPA/j7nsCmiAHpgJeNAjfuEs95kpkgrBypSgDI5AkZsh5
9TmSIFJ1Yq2dQQHAC0k4bCpTUgzjVYKpeVNs+0zha/tm/f9ywPliw/0L8E2v8Zr1
/DnAs0KApQdBnqGJby+1yeDHG/7jMxB4flVQSffwMvAbYuEYu9Cktg8//j3YMMIi
4wWLioocj92BnTJ6AMoHZwh4xywVBv36QjrymBlwCXRG9V+jl1THtRB9Lr6tWgaf
5weN1e4M01eoIEBHhlp+s/XOFIUQTdXcKydSOB628Ym8267vf1keAZwkbaThVzqr
rYFi69yXQcwAq56jIJgyGsmKJJ9IoEDef4piwL0E0M3EGVLrYOnb6e6x8hQw3ZeB
7ksadHiYrZVgSiIoA2WYAm250c6pY0Wex1wRpnTtDf6YhIkCZMKq2NCnXiwpEBt4
kLYwTHvOhbn8zkMeC9ybIsqkSqEWF/+p/irgwKPFXjyyYifv7Dn0D8YkRWMt4+Ie
6X9bxznweb+0uaDUmLulsVg/P0rNncVTw4n6iN+Pa1zrBYl855lIiEFSkO7tTjky
NroKYHKpxGoX6Za6pNY8q8vWmCybAWquF7drLEudEsGClQ4znWr5Y/MCYAzic5rA
CUsJg8namCHGIQ8mj7l8qFGYAkbzgX1T/sjTlngwwH/ie5PJhkkzgOc5lBt8Ljx/
dJQVzPISwxv4mGgixlZ2B0+ZBE4HjBuPYYR8lG0IzabmYKDT7iAKOFZhgjEiaEvR
zRKa4bTE5EPWp1h0I67UAfhZlaXJVxa5h3weQIAapziGfm8Oaj6jjtB2izlS2MdR
CRrxRvCuztaQByRM4AbB7k1vhr9rnS2+u59yRbNLzHyFafvIcH/gwdIHWs8TE+sf
AAIUOBVhiltWf3dSIzwQKJWYdL1hBWsDLyGzY9DZUYtjllyiPPjkr92afYiSUE6l
cdAP52flUpSDc9gaKY3rRYcxUHxEw3BRlCtbBsoFH/2B5Jakdj3jX/R6bFWa5IWB
nR1HeA06tB5UglzOTg1TnJADXHDH79jKsdXOoAoCu/eNeTocwAeegFyEtvbunMZM
VN0Sq5yE4oDHP5p4m5TqFhRvPy2yh55OVzVtkSEusatkFARUJMiNLSM9i0mgwtOR
uBYF8P7UjqDu+JG9zb9FsjrAS9iq2eB0rssbQeA8ksltBEj+YcbIUIC6UnhMSziq
TpCGWFPlMOrGGLaNVwyKdoqXXVlLsgoIxf9NNw48PCeSYU5jiCWzPSGlyxH60bR6
1bc2mHfen2qoUTm6gsirtq5QCPO/jyTHmPX1sb1seSvx+Spx94nE83r0+EyihB7J
xqIA5wm8iDKX2gGcffmVs6mJYDGqHOdSob0bxvEv9bzTyodF5p8qfsNyC4y/0P68
c6jPssv+Cri9E4XUYA6DxSt/edokQX3roJ1B9JzdwCfd1W8Vc/jFMpzBLjgWWnMS
jMgvDQd1yQmcjXFL1g17aK/HJO2Dfe659yr4Px0xQCqZ4gMZGRu/C4E5OYPSZ4g+
BVfI8q5qKSNXqIw/YmIBTVn4qpo+FchXZ6DvAx4LiU4il3SjkpqvbWMVCztFobz/
te6N2/FaXN+ceBmbioqinVaekPgugezdbCpjPkySqB/OAENiS83JYXRTrW8NCqrj
jySxUEv3LgK2UbZm7xwtIJsVky3xHyNKmoUPFijm4RT9ui7328sg1PuFyl90KpfN
fdmdZKJMjZx5fexpW9HclYogLef9k8gLNKrINBqmiipgj5KHTqypUpdKoimi7I/m
jjNt8XePaV6w7fv20elJaPFktn+6/QAEYDY56EIzeGuY/pBpgQXomoLIKgYy1M3V
/MlTey9/P6IuWPCU/i+3iFNloFU4I1jGLS9BCmV3UZVkw5mab3D0QxFvrNscbPD5
oQZmwdOTsGmEgX7m8Yq35XHn5kAqglPw2wd+PWQWMbW5/jVtjwsozzyOkSqGvshH
Kd5xp3H3gxgDzM/m19XOwKLVVkOLZjJ1RBLdr07nQuio3Q7lXQj2Zvcoyd3CIBRZ
eKuU69+GcdT6SN+dUqhR9PNPHqxjygp0e6hHn3GqHNAsThGn6vHjzg2MWjpRtA/d
xnwr04tUDu4KD/HBWXx5iDV6Pdp+0HFeBKp8imObNnpEgoNgJU+ziIJdfDZCpgYM
zupdsQo7z06Av7HG9PWPW58iPeWeYIhzt9aDPED9uocfgWOwN4KmiAaHnP1VjB5I
4ABKls5ptRsn09lBnhKJvNLZ6rwu3V8saW9QFmhjxeov8tOuoQjMOG81csPxZ5q2
LiYxHZwguIm/4yIy2k8E0imflNVfO6XvyhVNBZ+l8F8ltptv618iZgvmyHkIyiI3
pF3s24n/fixTFY8fR8gPQdd8O1vvD7GvmRgwPLr9/OXqc0rpFA8tO0ur6sJ1cjbS
k43BfB0Cj6nzUFqvPEuCCE78AnP6/d6Ge2xZmwonkr+DZK21mUeww8rb4BBCSmY8
rUErRXVDvIffMrbakHgY6VVwEkcLkH+PTQhKYJ+QF5YK+8gynD8AW8nQy+HaH2fD
JyY3OTHkafAyGZsKzn86rWTNlqtsjNTky8pmZ90cIq1S0+cAzo9F5ofTqLxApYQP
YqHXiBs5mTHIO8W9uZ84BnIVk9EzzloAkicMUw8MTexSAQcbu3icC95cih78eURl
SgiPGJef5ggTMAuhDYlDuxo00lHtPeQMWcXfcPDVHq8mehrkqHCfjd6WbnobzbFT
PwKGKITqgZwHmPTjFAtV5KuS8IfPoxvjasP7I2VZgJOqYAU3SCTC5PZ0ml4EszGF
Q88ROf6RQzFVMOMrsjsZ3LZKaOu7xTDsCZ5/Jc1YMdGCHYoeIWYAvK4+1jm9O787
QUKzNTIVachJ0OKBGG5IEaB4BGEAgsiA7iITISBbAtcztc0VJ3AwLUHfMFbtFjfY
3EO9wc0NnP/fsPsiMcMKPZyanQmf8mCgM14U5CEbNogG31xmE/zSQHY2RPeFRWjT
MVojo2y+Llrkm1Zd/8CqXbIxfDpZ4V/7SW/iUb25kVYv/vzlV74Q0FT/ENpMmJ6l
dLQ7blAU5/1e7KB7diZrAiifS4zRdR/O8GQ24mqMF4E7L3kvoNvLYec6mWFewgzV
zk6WhD60xdGDCw0Xs5Dl7ujd4FM+VLFhR7sn/velOT14vlLKt9MB2ME2QzGgzsHl
sSMP5kcrsmJmhzdEHyCoTC/MGclzwcvw2hIcJLnlUItx4Zr6QeLL/33VDhaM1/OC
wI8N9A0+r4l/LO63tuOSb6zZI7ZsgVCmOMCkhlbbAxMl8CZtrY5vR5Lkrwm3T0OQ
Ju4cmhYSVfQNx7rBmwwy0JPzdyRI6JH9OUSZIAXnu5P4vatYbN/asM37WJQJenAU
87CSkCwY/ukmhJ+KBFe7gh/FoQFNrdlQY7dVytMA7uMDt1+2IDwFEOo2PvaMhl5/
3PujEaBxEvCiXcpP/qiykr56dIHuW7i7tqAfeMmFbmC2OfBILq6IPWnpSJWEW/ZS
uYTqWn0yIcFbkbIl0x0VI8GlmzH8nZ6Hc3AMSeBPc8uX2V6+PDNkV8VQfANkgNbk
dSigGQBt1C9hJLVlZSkvtlMPQZc2Zj0aAHCDyPWim7Vy6jAe8W/FHNRTIfVessX1
WqirV5UddS5hQ0tMAQ6lN1EU/Ka3MBY6X/46AK+8VRHnGZAcwGgnPOzgWN+H6sZ0
zrO6VMPu9BKMOoplYLW7ofK2eXqNU2qKPkGeL5R5dsh74boP8otXm6J+YAqPPTWl
YavZ+yh0HVbSPgPbn0YovWtp8i0n1LDDr/rcI4QcuEnXOh7BVQni4eiw6bO7pxb1
mTCkVx3D5fLeM7msOALtr/UDMKLwwWymF6bY3nqNIlEsybBuezgV+zKpvEes3sv8
kumVM1ODAOJ02HCRxWwngUgzYyapMAgHLUituTgJv5JNDdX6B3p7rRr/Fc74GWbF
Valk+4DVuoAe65pwKHB3YcamxTX+CA8mdiayvhKtSFRSFdZBLW9OV07GuBHFK4Z/
bJdpolTEHAdtVVRpuoiklZ+iKaojusM58d6IknVcSkuFdzoHc5kJmrOIrNryJLf4
wk2BT495fNzFFusSa7tp6AbsidSJabEaRuwbZZ61FPChSCEfQGFsTlcYukPRddX+
I7h01KO4ul6MjdTRrO5yJQkpMdhwEMyJKM8CAzhHYQjEr1jN4UDztYDphhiTl6ET
I7qnA/thao5S03MNBFufEOAuurdXO6dnpqAnG+IxTKHmWjYVtHPN+7OWG1xuDhq1
bpGG7r+NhS7HcEovrPEVG/WllSPclqbkazNrXYUK/DZ+WiFeBTo1M7DzN7WPIrSv
iRqiW0qxTG106vL7rZOp30o90cJbw33xv4XIzJzXNudhh2kjEjsfcMGJcO7XSkSM
ouKx5UZxnYiA64SvliVuutLgm0P7ay0nO423RnQ+Ohj0v10VG1mbbuTmZfNZKgZn
EaGBF3ahGi2jZh5qe+p/veIzzkujLiY63ciT6ud391tEJCCYWy/NzxNpPTbBXEb8
dK3PAZvxKoK8gMLiVAup/+ruRArH1i8ChvntXDQs6fyOQeCCSHTbjoQPr51567Pk
FLuwq669YYPnnmf2qFO6niheykWzcb95i2AKRYKeqUNYxKiKc3Lm+LwveAIGqvo+
IoynVRWdnFO+o4XgpOZrWuDMMpfIf9hGYjCnsisgmrSLtcEjpcTcxt4lybi6sHsq
W1PJB5PTprXvy2sWqqM8BUikCY3+au0psOIx+mpo555erJ5KE2hfCbZ/GHYl63S9
oFz33SNPIvDGW8UjtcMjFqoUkD00TkyA9PBIq7ZFHtCupsQaUeku6KZxGhQwn/br
+CbnzwrTIM+9moAD55IDI15JINEU+06pJYuF93VUEzD5P0vMD/MAlPNymI8BPeLK
12imgHNxKRN1vQhIooofk4lxNetS3/jM7EOw9+93Q/XA3jp1lAB6vnWcOQTZpeGh
xr4NAlfjg3zX4oZ/mpc3qiF+V49HE39cGPeVWdFderLHMuCoLkcfvpQlT46ddyXF
I/bskGFwjh4JIrNcuybu+bWfbXBekKwE5IRPv3pIQ0KKkKgBUe0iZ8YDnkEHtXvB
Iuji6iflaA2jdUTjSE3nUa54qBgGXpbS7Bdk6s8LPmgdLGwLtkfWBRv5YqKsLSYM
+THrN4g0ERYEDhv8SNeuqR3O8FvWXVNsux0K6Z0lkuZEibeEzIzjcgGqS1NP0lyr
IleDu6nt9GtN7Xuc7idrdF4k5BXLZvjRMJm/Gex77KnIw9ILBflCw6gEgYbyHaFR
s3FpH9x5rkxu8bqlYgP2ZA1kz8AF4x7aHpY7oW/AenqUdAfYg+nWuEkBkgcmx/ge
rZ/iv5ayTyqkG0jqDz8EL3sV0/TIYbmoxorUFdZkdMUoRF8pOwoarZ9X3AxPprIz
5XBLPRnnx0d7TqolqQ0J4wEpYYp4i2JIae8vVeAWvNsHs5ebS2/vCw1LSV9atRaj
EklZ9RWZhgZThDsbmAkmwCeZLMs944vSIw4pe1mfnVpdSB2IFyls4po27N4P4JXj
pUGLzZDccvDFTO6881C3wTI/W2AXNYK5qMc+fO9XpKY+GmMeXqUF/1oYZ2qNO6Wq
NQB22tIJDjiM3zdgjK5nJjZErhpAtPWsTjJWUbxjA5XtRqQoK4u+v0G3xqCt4E3U
VwmjPr4QvKdqTnQbTDKc0FNZ9877rQ2UR1D0jvwynCCcgG4ZXLFFaBuP2uk/T6Q+
yT53g3cJfWWoYy3KSHnm7OqED6QgFcrCsknx9z7SuUqJUWbUY3UAni/ZCFiBEeU3
MWN2pLiVCumll7y3Wr3JO46vusWAB0p3VGGgJ0v0NK3KsqiQNVlt5P+MI0EZrmHG
NYm6CC0fsW1CARTyamrXgsVod5V6wHMzROaNpBK0NXyQXL8mhOp2IBH/6POwAzqw
xUHXmN30yNySJ3wdQiJaUIbt0oxf3y/R8YpDSgA8zXiHKjkBzMXC4PjBD0aYS1B7
M2VjSTasFuqMvioeXmPQTrtBeVUoh8os/yRyMmnLJM314qD9uwe+dwYYK0Dt/Ljp
aeByZSCp6yLp5d+GCH+Fk8JhWJBqsSIj4WwW2f/giiB+AbKxje73055wA8ZnMKYt
OMzJKcRdCut9j/gMwaEgDPAy6IBpLR1U/a6DKg29pjiQSB0mGialnFq+enfnp0lK
KOxem4Xz9OqLwg/HKQVviOMCpfgskuIq+umvXxcAb3veSQv7oN6Cxs7cU8PCzSFc
OcuWePrBryNO/rKlFDpW8qq0r8BZYk2GOgFvE4LOMsfRaxYKqwyjkwvKk1PO2bMN
KBh3R31ecJ01YVLozNTz67TVvQK4UJzZo75jK28p6ou13S85nQyC9e5xR7hdwrk4
sCDYJMnzzD8MODKt8G3cYOYQLrIV4qjjlaeF0yXn/ts4P+P+1WM7syOabCvfIP87
NLUjGTU4JnhUm27Guar9Pyu5xaUhtJh/tnQHUQdewKQZcD9pJZykUrMF6MilsiBG
nqlM0iNzdhbYCDw5xeVB1rQY3pK9TlB9k6ET+E7qTJRzlUxde3DR7gkIs/2eGgyp
BCHIMD2FBhhyn//9Pip9IaO4VcKhA6/K2iFM4waZ3F69qLNW4P15AbF/FBMf0sMX
tS5JkKYQvHw5TfcSShiOp9diDYKJti0GsAuj+L0aYfzwBzAqTnufwvx/AIJ9hzlq
AVllm0C58V+YrH/IDlsrtpHu4TrnZvmmQjl/ONS37X1SUCD4oGlhHJVwVDhxvU5W
45+W3RmFog7MU/NADlEGGdqpZNL/9DcLrEwqh+9hAqqGssExhyaOWWIorEtzEGEN
XGyl55EXY9JYdNwFfZ6WHYAVoBRT/qVAbFm9s5/4ZUQ/NvjDd5sCljocVmx059/u
JOIwg40WN7l9BPfL1tHAuNEtGaWZ+ebDw+Q49Kiu6eb2YrKLsxdo3VudQVk2xqzq
2J8flZNrirPXsDLeworbm831+YyD4jPQ+S2bOphvbyOfzRhSBbNrC4iBN4FeXIEN
Eg9G8Ey4I5dVnsYewxM7OMHExYQ7fMrC5e0y83dBf60qGJ7lzzWQXUhFA4ijk07K
8jq7mORICIEdK4KHaFcTjcJbPjtKbq6kr1l+LBOq3tZcd904H3hn4Ss7Ox9yQz/e
qYuqOLmgSAIZ9K2la89ibwWjGUxlTWp+wkDyMilimFyzPraOWtc5r1oaZe7rzh1r
jTKL2PCivISsWi1ygMSZlOhbBCP8cmDqKDLnx/n3oLRFAIZ2U/9WMcaYzrBTipcX
Gem1mXsLd4wCtGJOT5iW7TMS8+KbPB1mr3NR+bdYq3yTxM3FCkk9BEXUtr5RB4sM
Dpt9S1A7+maKBLaeBfGtZ2oJ9MbQP1weqIepYfnaRjyrTUrnDGOlBQHBoDBKANdA
8Gp4PIJJ9V3JLoaUQ08uuFW+SZwSvQwqb6k9eRGV/vVCfCIuge447QBtbhIVWjH3
TyebnwV2+aDo2yj079e3VyUEUgSHqCvyOpKV1XJCQX18a6Qo9gXYidcCmngoiiMs
ksZvFGpXTnqPS9J+8v/qn/lbEZxz5hIpV2dIhzJ3kQnFW8NwcJEXqTS9ozM6QUCH
e5+sv6ImYz23PHjWOqMQx0U207Xtgx243d808UyNtLxtuzSa8kK0pPy1olNW6Jbp
k84lFmeWcquCppboWst1ZmKI26/qXZegpn5A4doFRe+mJyoNQW52ahvnnO8PNU7D
KeP+YkD/tMt5EmrkMErrTVGMNu84tbk3T1EeOkzHkT1m/eaqODQgmo69Zf5FRc/9
lyRWksTD2tMgOmz1yeiGU2UdOrLvLCDhYth608c92PgZ0x8Qe/AwXxg0Ckz/fMWR
/PHNo/jdZtmRZCgVS1pxpejONaqbQEO9qezL1QiycRZ/eEiFkMq319lxPjC2dVNj
0raAyw5M3AdkBGgDAhJAC7H54Tl+UJ0FV9DhUBQjfhAM5dwy6uIhSDPXKFdL/SGd
uWWujQcrw5nvxcQAsuOwh7wgyhgexiXBKz54LeFz/0EWrx1WN571SKkRrFg0lCOj
0or6FVSjhsqPXstT1hbhR1HouketwFRXVaAqPH/KL6AlzX7NuqmympGlUm48yXUj
2bcXqsQbSBjQIU1TTyewOJ5ws92mc5VZ7AOKqbxmG6gtcGfDctdsMhelvtkTLfwv
F8oUyOFU2BeeBqt4vjOhpQbMZey6beqKVbajmTMr9tcWou1/zZXH+TTc2OG3cJ/O
5OOR1eVBfUqMNsAYPzFH4w1I8cvq1s1bM50RGJlXzs1dQv6EyiXSfNDGFzB1Mkxa
LlQfQ8xMon82FYmRWplv5lx6HucrZTp2JK8NGADqholxHUKL23M9wTHUFFUIuvrb
lRHJLdtFkFK5KWdHo6NN8mJVt0zooXo7stOhl8wadgwjNuMnNNuHEl1e1ydZjdm2
P959NwhSI/R116TBa5OKcsTa//HclmaZ1GEVGJbqspxorn1DvZwC4n8qmq3oImG6
IjI/TT9by6ZpLjXCdiwYZ95ZbOO0YUN0PfuLUWYxa7LxbpJMeyG9F+KARS76aU3V
OAmqEWiXPmcNp+PHvu65KEXIrFqIFxyvQaRJTM/iHYUvep1XwbclogChhSjWbqft
dab/t514qPRTVvd3NQrdDNaHLMDt3WNR0zNXH9QCSaVfCZF3LVgtxRMlTMM1oWDn
mFmMM4QOQ+DuFdZtdK1e+VV8t7zQ42YECnzI2tjnItaCgn2hGySxJVEqvgCS3ZLm
A5y7uwAeXITWTIoUwotN0QJwAeVBX3EbXwwmO9T15MaitIC8OfAxLT0yA9QMzJDY
L+AbfICeKiiVTH4nIdW0OFkMvJoKbYnBmZ1qod1mn1RxQFPD1vQDV/sAgvZM59Qv
XNY3gZ46seD+6AocdRZ8jMvSSg24YHNR72BqOvV2wEcUX5QcSv5UIv3GtPonCZWp
jkIULAKYxHPPm20SBid+pTN0k609Moh+ex5T9JoD7v2sX2Ow8MVVsnxNepdCKrRi
v5tOwG1lWO2z561B0/xLyqivJU4LAswLNOKBpFNfqNufEKmena6EgJphEOKahGGv
nWE1hLIO9HCwGGVOv+JVCBd0aKkhC1KmqIbPhYnx1uEfwki/594sX4JAJbPwdRUL
C9YR1+tcCL/XVyHLp/Ky9IwF3le9YlLhu4lpukS0M8MFMPfSMbdyHuPqfXy3a7Xz
Zk8asKeP4K1XOMFVOXwBZ9hmqVSZH1yK+nfB7Nl4XvnjIaCzmYXfstrSiH1kmzav
Rb1//pRSFExiB2wgqtpVuTWHYXLZRfyQ0ckO22mD37Cyb/KeiPE2sHK7lEHh9sTj
ht7UgYsImMpsYAeRaK6lS3uS2aBb0BSVplywsnE5/4lZWDINi3l8u4FJR/S9yUV+
6IRGd66m0AyNi8+Du36ZL1/lQ+sX3llaRD3wx0joPky0sV8M14bg5sNxDmvPuo3p
3pUakYq9IuUcp7uNB5HxbLaL86C02t4QYfv72d9IiJ0pvXS8tsYw72rk3v3B0N1u
H1w2GtEsbp0zJaPYnuuo3EetFnw9j68q8J8v7lG6p3jDCrDMtH8JoEMQRxw9DDMU
Q8XGf43Kduqj4du829pLtfgrhnTYgf/+pXS4a3C5qArjoI4PG4tQesyOiQqPdJIq
So0TFS0ubfZaS6tNtiArUqTbl+ZKnY2voSmKErVv0Z7IWHCH/6SWDr3PZ5QpCyIi
iPh2YdTkL/kPa0wS7o/EKPRAnJvAuBJkkHuJciXY+0DgUcpZ7Sw6qMNA9esje3e1
ONLlDna9Mr6PPQ9Eb702ek0qc8K86kGcGis3v/V/AaRFGkoRnJKUccRT9y9Bqp2n
91nbKnLPu10nK2Zn+rOkRQNNeYRZ8snVzdEsvYVYnaQW7812Udsni8kgS0KYq5DR
jKuh0cKzEaudFe6S79h9V3juf2OXtwmdEhQlk6p8u/pFKf7lrHH9LMgUCwKwR8UO
8J875hM4n3vtUmlp9sFqpAnK1I0m/bgpjoiMqq2ITP8uW8EXxuCjAVinJ2nkRhjl
+3z/3qle8ray4UOicyG31MbPHcAvi8FqjisABbIqRMmlxCCoCz/W1CqUs7J2Ah63
1y4E9kQe9z83OFcKK0Pv1Vf7pzEVox3Ovz20GGu0PFyjiJRPbbIEPeTpsAgZ+JOK
7gz2YMO3O2OxsWVVWKvl7hxlgRLVtDgk2YPJIurw+AWCbaftPdo4G0E5poXIom7f
iUPxLYs4DvSBWZiqs7PX6iktwutNQPCn/v7TjK4vql6mkSeuFcufb43BdB8BuDg8
g9UttsUhdn8ccDrHXsYETtnLHszrpsgUjgmNLV3E+0RjpojMqkLFEgIG7RJdt2r0
UT5y8uUSephWkMLfD39oFM6FI/5LM+YZim7s+86n73M8X5V7huEjHfKcSjcfCFSA
6jr7r3FOU7GY8eju1UcwjxIWB2xHnUsBCUe8FU6Mg+9E19NbhWFjb8u7Xj0kIQZB
5v7wwdrt3zUR28UCRdllKNV669fuHqnOfvudqQIKUyUWRZ4cUX5FU56E+mRD1LJh
Kb0HZr4x+xtk+a0coLRjxYw7gHSWfiSUCyOekrP++hnzb3l5xxS2GeUkr4+X+5y2
YieRJRsW4XHEaZGKpNGLeEbiz5gdeYffpnBxYOT+7f8oi1jpHEbxS1G/vh6HppWg
t4gAuAx3QbmXFseqQHXim4Cmid45/COPLXXNTKf3eJdQbqNXdiMERK3FkN0h6Stt
lbF7KEbcjjVNShp78AxCVFrAa94SJWvY0gnJjPLrSd1YfK+ctgKnLSMalj019DGm
x+R2RwNxgAN4XystM89a2lvF6viJkCk6uENQEVvXaHvrUfDBZfcdFUTW8Y+p92JH
dd2eetre3Sfs6XGiNWgDQ2JAL3rgCHb17+IBuVYHMrLONpVJB9hlHt19ZoPwQtxk
rROBiSdnm+zbeN8Iz9R8H2dahuRvfVfmLKdxktapaoc9NciheEZFRkebgYg207Y1
Uaafv0b63I/r8uvCWjpFoTNFhfELEolHhddnbiTe6V0o48DqAJ2LuNKPceHz6K8Z
bN6S/ncDhtEB1+wWKOjNmE/Nlcy4mMK1FPglmpT8JgFqV/kvdrHugMNip7MZHGW0
aHLopBvvE4ENfuvKrmbTNpR3AZx/THOOc5RHDsoR6yN9uBNGFs5IYVEc4A76CDc5
+CCaZVT6+ARgHi4yoD6vWBqcEiy8Iv3qy5FoGOK7gZ0xdoiaXMaMfmsyY420oN65
N5OyUhhe4CJeq/DgDyqCdYgY7M8kGo++QFUb4hL1bZhW94mcimWnaxSkQy9g1p5u
odc3W9twiCJWq2evNAWg3ANORzsSJGUmNfsvYPc1lHPbcvJbR/71IS4wS/0mpe4R
fIzBousi6/csB+mvV3dH+rL/JMqcYEYtFSALTMVp9ZjdK9ax6WzUjdL9smVcKZNh
hn7PGRTcZxph6waf9sFlXUYYhI47maamO1SCP0cppRNJ0KYO/lY+oenXGOEM7SG1
0x18nsAno7ngByAEMpPKiMasCFFOtiGxnslNng+kuBiebDp6l4DcARRHPTUYZ95I
JYs2cd/rOL718Drwfp7iEskCO2LKjygn9QSA8nbPZJ/r+TvOxftvNvtkS0x8g7Nm
wupfz0i+M02N30IKvGD3TjUqVC0cpU2J3oaXSsle80ffFACL6JKrETQaaiCLQSNF
4/InL6cSdbuPK2V6jYnwJ8ZxWty9xuQ2HmNi9V0375WdXT9dbkaYEJWQA+jTUjYB
abqnkpjFTQ6KDCLvKRIDeOaQbrU3PoTzkG0CuQxH4fx70igw0ifcEaUriWxbofIS
i478W4vTFnB0f2/zdwHhHZAsZS45h8HfgblAO8NigcB4+48PN4OiZky9Yw7SBg0w
IZav26W1VR4+xZXEIve+OWPH4Costs9G6knFbcQQBBTJ+xvdwphZxLeU3VxxTWeC
9Upk8+NktV110sEunZLiDaUBuUo0BgHCTMp4DXyViqPt5UDUYjU5AiOA9iTe9Pva
5DlgUaUlJw+LnJnTUAffsuBmxHTf2KSdg5XMiY+nx3W6OdGZ0isjRUO40G3UkmTn
yEstTeorQ0WhnBIHqWsxg655DdEtmjmvhJ7f9T2DcqrvkKvIK5yp+yZxpXRac268
Z0O9OXwSyBneG23myJY0WHPCCMOKc+HJKXIquZG97lMmNq13tK9eHqJxQNw6HLOJ
XnS4CGAR6RyLJPi7shf00XGvbY4MbB18C9oj5hjvQXn/VbvJSfCidxYvAlUpU8u5
vJOzMNH4+vpNK2jtRFhbFdeBH82oZ6GPX8GtFwGCipk0Wj/Nz6+0XAh+IYKdu8iu
sm2rMoo5DScv001ob6xu/opjnUVDM5AezlRpzXgjxbBEiE+mCNwLGEbd9lR4ZEB1
SPdZ+W9XrzT7o/ytEn9rWrs9rN/Rvt6K1T1DRayymG+fCD60MfTV19RIb7ptzBd4
DWFng2gXW9ysKs1GZbLxxuH6EvpurdsM3L4zPGBNGcEEaHxmKk7UULavBnLqezxQ
yzriGzNNeXXMGUCvm5ijt9C7JoCkevjcxPmcobdT9lIl4U2sQhEx0B/0VXlDFG1k
cx5gM1Ev922RhDOk/oBhyUNBhUQQintzWJKn4jNvJI4CBJpw+x8f49gSLUukyzic
Kr246a/thwQYb+1glfkkWzm/a8KERz4XWQcZri+aKg+O836ap4+ZI6FwhQ6vVESq
Mnl8Zh+JHIRl4aytyaBoKlCPCMZhDQWIdyPcOL9SqWP/Tc3RAG8FdUE9m0QaeLvb
v22JGMHLQdp2OoXPwpMz2k+miGUdrP6ca6SV7afvLHFWEpqpiiGeG0UwBWR+WsvV
iYLCA4aSErRVrZpC4JuktHvlkeYqMKv/xn+DoWBU2LWZ84+7s9ccWiO/3aF5KIb3
ERH6k9HwiCpiC5XRgjOQW2GWaEwiWWeUooAbt5v6w2e6WyWtsKP93x4bhSC58Lbx
K3gamMydnukF3kIfN0+h1fJw4IIPDU5bI5zkLZ5pl/uSpOy93h5twbjkMVN+seem
l/Ai/JPs7grBAtj2peGZr5Vpj0vCtSTG6fs3Hfh5nKOofWQaGA7E2vb0ob0AsSIm
ZpN32hrjr8NHyRUOeqJVRWiqkxr0HbtgvA3BXDAHqXghmQ3ATZ5buMIpOBIliIBp
k1DsnsspdmmqFnvLETA3bfb045FgGXEz/eW3P6LpQ3JiwezEl6w9JYE93U/H4GEs
FZQRmXIrPRt8A/ZcW4eUNGWxkaqzoawfK7Yv+Q2kSFDNuiyrFdEyg0Z2wcQMMCeM
S8fMsKpOuPVink2CHxaAegnBneytoPl2ZwwavtP0Qocp/3ZPWmtGiQl+tAs3w8ba
9ftvda/vQCV4OcpTBwQv52csm7rbLJYnBulZ5eSOIrGXkd+CI8MOFMmWuj689+ql
sbzqV/fLm5t6F/x/2ffJM+EDEksPO3iNPVYxvqR9m9PbawpE63YOtNpDa2LWDvYC
DOtQr6qXpZR8LMcpqMccQVsQD99+Y5fjPSMme0d/agIiDKbsDpwf6yvI41UXPLZo
b5PNBtHts+/GFDJd+76j5bkC04AfH2K083qpAe6eLggvx75h80AUy2kWU4mnNa08
cvNXDFKULq1NMIyC7bTUytM4hfRGwfBm+pQoSVZ+Nm4M+EV/NfOnV3mUoQV43FjE
6tUPbgXNsttlDAeAswPYt5oXzwlJBqbRIg24szEbiKtTAda7D9w5lfU6UBUyria5
loBu28ptXletwsj9VWQiPrhynYun03HWuq16T4cliLVFlU5IryXzfRTNKLcWOoQd
t/8jF82d4L8S3BccXPFNu/SjA9MtBn9fhNFFSiuCtKW/w9x+ShSPtm+ykjIXlN3z
vP71MGMZzVHd5/H+mTVigpTzv/JOXfWEzOBb+3C9zsKUWLUeVmtaVZA7v4SF3nnP
LyA+n2AdV48/FbhTN4gVrbcCzd9Eh85AZh39YK0jRXWfY88TRhtXHksK4GTELa44
3/IVIUpx1SKn4bGH+tVWhEA+0pJQVrcQQZCH0OG0sU/ls+lMqLp8FOQhqxz0Xfst
e0iCPrInvVrh16hR+Qzjp4dXX2KnGsYKPR26HwuY/dijYnUAAP0X7Q4N3SE2fTYe
+kufrS+cZi6qI3uFPGvsufogrYuz3uG3IxypvC/6l6Rin3A5Y9B12RsiIL1lq4QX
cIB5DS7mL7abHXHL7OCenakXgE5tdaCv/Gfz2htwKWZHFFETf76wWU3Uwy+aDQiJ
C2SKO4h9zoqv1BHmWzQmEc5XpzULHznsLi3qh5cFXVH7XuJYbfszkFc4QZDgZREP
rhvFAH7Uem//wB+PAYkNqbOsSDVnFNWkRxpOGRpzIPNVqVS0yA7LdTVoAx1xvOTB
rJ2iotOhm1+571HSOByiT4itRjKfSAEH+wX90paupdFS6+pX75lAlZSp+wTeDbK/
Sz1olMXuhdhHJUPS1vCBEmb0v7cgko3iW7iW7KwYzAh9cv9mgHydC7ZAOajgjWXs
Fd1CR3zls0UYGVjkgcJzKFIy3zEEZI1cJm0YN9SoR0X73Hrxuzn+doRO+45Yy1Ui
cuDf6tcJGxNEcb4yOk9qntwDpNoPeFovMqKrGuWVAxndCkH7Flf+CMxS9TnUfsWg
RSRhbtXMUKjTO0K/QJQ8H7ZnfNURH7iwAGqgaQID8CWiuoN+wuZBgWYV08RAk+75
SIkNvouVg9sExaoPcXyfWpSCeYZFEV1D1jShFZ7peFMiP3Mu+8sFluDU1nZpuWN3
HfkqP9ng6K/zFtc9Da1RXHchjBLsHdZ+yYcKg2ZGWpsaFd4r9KIX/iCiq5YFpMPz
O0Hik64lHprSsBYPaMvRq5i7rCYWXHORsrce6rYdCfGpGdRRLEQvjBmZi1vZS2q7
44hGk3ugVXutfiTIoLXGGW35oRrV5JqzICg3llVR1rloAZTNsU1ERMY7jl6ywFac
WvRRYksx7R73QHw95WYZwZiWpjpGuwOsutN56RCb3+QUxmbHQtpij/VZOppEvGtO
GcrdiTLWc0JDzy8ufzx0IrccpRpQv5xYJGlTTTZB1uvEQ5B56afq6xwnxQ0AeQtu
zf2W8pYLWKIdVtDW/GXAJ/F2nNBWOLBN1TTwluz7/ai9c14/U/6Qoyd91O/BpRjL
Lpj3BErQlMAYbxEAoHXWMdPD+aNgyq1CKJaYh/i7BWGkq04yd45foM48t16c7K+g
zrGCtXg/s4JvOpUQ69KH71qbxBLzb0/ivMOPVqFG75Fnv863gACLhB6bT8N1bLhB
Xuu5UNReekDk5ui643nfnGE9eQG7Mac4A1W7kk5Jd12YYQaYvyj4wjyvSikrUoC3
LNKMU9iM2SXrn1JTrHG1tqicqeLz1y9TsTYuIYvy2UvIZu9TtGgcz2N//FHog5J3
IpVfhSiF4oDO9Ae+TV7dlXDjzbQCCBOsCc0bxwm75ETe+pte5ckSjtPOoAQ4aoyy
oe4A2pbFkC+EqabS6jsg+CRWjyTLb3+mIoa7mM/NtXwAsSudKCcDIFkP5xuZunhd
6qTK+cXZN1cg00joClWExctxROaol+btfdlVYW58wxyKtHdlryA4An+QdXzN+YzJ
J8Z2jbpdWUdkII9v2Nc6KeWNkFwn45rqQQ3VqX+Id/599ch8KRDIRJwCdkB+7vJq
vsQkmXF1YTjU7GpZDV3LsHiTedfenEbneWj1w2UTWUqJo9hGNW9G2uL2EtOJyM8e
Ze+kynWOHRIv7US+VCqBX2MzwVIny+SzEVB+hbMcH/ObKlnEAV8baCWdkunYpEUX
hrWxOoJdqVEKuN9Cc4e3FJtEmbbALUPP8LEswQ4Qs6gqPS+PZxn6h464fyA4PbBW
R9/PyW9jUF7kkBJhhHFVQl6kvduqmTora7ek31Lqa1yHXe57PxsA8BPpVp37D3/e
bw4osT8smD7MqOoWYcVaRzY8GdYjjNsImt8tpai1SMagDqZn12Z2/mQibDRIoG08
10dgQglTA5aC0j2/5lYB3IorRLVbmTv7+KvGbgMFfp+F5OV4bZdu9zk6XIJeuGMl
iRbkPnhzIwekICIcZAOOuJTdqz+iFNrIHfZrzYzuYsFZ/CDNgVeYNS7FA9tmlhBc
5uKYz5sKhNnop3OvAouLCXGbk91VeZ8+M+tXWTwLa9GK3z4/Q3aRLwz+P5689J+U
txdujZzod6+mWZl27v3kfkxJ8G0g/wqucm0m82K1eoDUhFTGqLTm+DftJvvBWzYt
KJpoQ52yRqB7QddnY24PrM3BH2J16pvskLlAbY1JiY5OWWlAFVZGxQp8PdctsHkU
QX9zIUhdCXfobx2hOz0PFKQfSGZLbq+HouNqelSVRwv2mqup6iaBb24DFoMWAFWl
e3d+0ppkQ7belYw8EvO2elU/X6y6jyuf9z19uAJSFR/GAS64//NyWHae3QkRvmOR
1SjGaNX2wxuahN0sUg3yCnBm14TGjemOpFkT27znGbzuV4sifSqlkqkNT2RGKnU+
CMix4ND1n3qcoombDUaoPV7BG0z+MspaKvcBZLARh2Tj7muniG6JZSRPRwlL8YSi
L6fH4ahkEg5IkIEth8XsoC6qVce70djy3DAEOuZd8rvRafxaeHNYYTbmh9qmxbv3
ZGtg6OdPmUze015oo67TzQq7bil59RTKeHX6kJ7B627TwcF1MRCu8xRVEC6T4Qrn
Trn/KKLp0tW3YpQHNsDnhjNKd7bT2t2e23jYxrYU/aSE6RACurMJnkDaf/K9aMf6
8lfySRDoPECT/lfG6SLzUIfdWeX/fKPRJmroWtQylvexjmCJL8e2TrWbX/BBU2u8
ExR9ZLhJ03tBXy6IkpKb8EeV8MlYdqw6HtysMJ/en+T6N+U/UgIa8YtNhhN7AQoZ
gWcn7rOsHT80VGLwFviRQL8yQMLH+OZL5BiROzAWGy5y+Tu/1QipsInpQCTCyxBE
pU4rntH4gk6lIF4gcfzhvb56cyVu/7+e7OzL5kivpasl3427RTdexdM1NrX69D9C
amcmRnv7uDIEi01Ct2lCD4lmxk2Q1FyUmIKVFoh6mjPfEJlAJ2SmJ6Q20b345wpF
TDP5GqxqrMCKB1pM8XUoA+OdYI9r2+Ts889NuryI7T85lwX+2F71JgN+reeuM9kB
GSrOoEb88yJnRjaGYGywbPZX4wEMftECRRlwDxJ0c2dj0me1p2OC8uZckuqA7U0+
1Z98E/NoUHisEGtUJysWr18PdzFP2rzfcwGeynphsm1DKI6cPGo6JAUYjjBRion1
bNMiuQpguBtSuzOlJseMhRNqqCIoo3AGZTrxb1dhlrUhVhhx9r4JjaFYcmMdkbXB
6vm20GvtYg7cci5O+aF6KFNx+aVHpNIEMcdQ8OmuFXkd597vJa+1BXfZCXhszBGt
8vEAoK4CveLbrKwBJ5CnqWpuTycaWkS24tNQxpdq9TM4nYyT8stoJcLdFXE66rRQ
1rLyGIStwV/3BrhqOevyOhhXK9dcyg+Qf5nId5QOVhQJOaS2nk5E4Tq8xDpIsTmz
8Zu0KjkWFyT6cUFHw2xjTTqr4HR0O38NrRn2IimK4TFRzPjh26hkUJ0Y1S/IDU2R
yXsjFXgiZn3/fIEnHBR65qDWFlWuha+L/GN0LgnZ/unBdKlUP9GymOglmhOIH02L
SlUt0izNrioES/KS4ebcmdBE04FBVIxKPQ3hJJyAEL0VVHoPGWbaTr1U85efhXEP
vYl5I/8hIC2rjlamRRfR7bi2q+IdPKcInYYASjFoP4K0twMdCvA7GbHk2z8Pwi9k
3867uGMmEowJ/Cc2GEOnCbXk4prMgQBHeCfgpv4jGjyn4vtfJV1oWhBLkSXB8ncH
IqxJx0wmKQ667Fj/3XwAsc8m+Jn2MhBNnW+9t5y8nA1+YxHudHWOO7vsth2qiwly
5oR9rGw9+/Q5n8Ho1iCjlDVZSu/XBYb34RF6c32aEJCl9VegsuW/eUnc3n5qmkLZ
ESw2hf0AC8u8V8uNkQNd6ONDxVdTNtVYE8lry+Db6/tzU43KbClm132e4rz4xlRh
GpOE9yoHygw59CMI7v0jzUOwNCLvg2bmvv6VkCfx6jmrVqXHLEBzYv7j1uQ8+2wb
sjdI/N7xnx41Zh4B9kWGr9JMsZnTuiu/mVmFeXP/io0cBuWdbElmiot8BKjtBUxC
7OOJnisr56grAs4rJprbFIiSdV4yuBWatMwRLU64xSx2bOgVm/Vzhxvu08XWr/R/
5Lxel6RBlV1qXOXbVddGooQQbHD0PIC3uLwvQR9ABEt0flRbjCvroiyQBFaBaQ38
ZqeC6U/5rqi89eHK0/Ingz7BstUsy8RbISdGAPJB3aAO1NvfOIMCFEh4YFGDi6V8
YkQhYCAHKo4jGe5WOn1TpDuffUillJ8GVpn/DozbFY6/02HU1pPR5glThuaKfUlG
3zabVuyqhPdwehHUnkuoZuSiWpuaAsLEpK8Ehflm/8eRdSP4+1NSUz49N4HfZsKq
HZl/cF8FHrO/mDRvjNqkkm7COLwb/wwYYcgLZy6xcUodCqbRCaHBOdo2TX0p8izb
cfFfCwktm3HGul10K577kYXlXKyY4YWboIaB4QknthP0HyX5oUon1U1VtYgXTyZI
Ey4MUXfeQMjUbKhu/ILszmjV6dgLpYq4GJLsFFnqoNC9qW3lobZ5haI7yJ9uDTnS
Jse6u1NrnPK7H4UCy5WsZ41UVTNUij+z/79UcZi6JX/6TWzLnKa3De7vzlgAvICh
wyRXsai6D+3LxgWdwjKTGjT8LSVMov0OIRgzseCuSIiFdt5T/vL5EQiqeFR1JYc4
VxJBl96oX+TjWb5/MlRYFCntSQcMfg6uHnN002zGmYvsNQ0pK58u37kW3V3sq93e
vcxzbgE6PChZrfWJ4fuW03Vawiww96W5kmEpB4oi2zou8ROnykm9DLvrsKAiApSm
q2/O2UonSZM1r1KKrW+DJ4c3iTYhVDIAp4R80BmmXycTS81f1s76IkUC7iaFcd7J
sHiQxWgDzghmPWLyjEofGhsrh5ApOsFrwNLLvN4+jm4PQUsyB5G3HihKJrvE3pow
GgTIH6nPlwoO0VK6t9tYCoINsmzYcndD5kWnnD7zLxBmcovRZiVjxxBPrnX2TZ3b
+Qw5LObhM6otiGHJ1iFlKmTar1VEAI8ZqZenZ7HCchY5/7PbcX3Y7v8LfkRhTWtM
7m1JbY5fU9WqImOyA2rwEcoTRGj9q0jRAOVl3wM+53jAuEReFY3jReeZRLnEdxpy
sMPmL6+JNoGoQf8aGTCSi18LKJ8HY/m4qGXaw9uZC61Q22z3YlS0Osb0WjbQs51d
iN3SK5+j/Mddw8q+9NWd0/qCKfduqHCTLOePU9lYGHtngRaiSks419va1idAL9to
pVOFh9/XN3iooaKkirqyOfgtfLCHY9QqRhwX6UxE+TrxBvebn7osmR76lWR4lPnJ
O6tyL1MT0tNfTBx0PvMval7j3AJQmUXe0JTjA4mybzDiUra8uYwAEmCaGmoPD/EA
AN7KIU9JdoDzAHhNGRwT6kTVo32zwJosjqj+HGfI2SdKPuHdarLKHdE1F1r6GXNa
0FUTkkNGmtni/Hs1G3+dPMfXddiLRF1lOHIQbCYyETwo6pgED20hMR8t42uoIks9
CZhzt/1792e0e01koUksSER6hSazkIGzjsSbitIpsuDxnqLzfOPAgLt6y8Mgxc8R
Hf6J+p1EYA725HUQ5XuQZxppm4xfSf0Dkd5N25zFBZA277uFKlpjHnTsMlJl2xhq
V673hhh9z0y3ACU+F3A/SVt2wRyRXQIIbJBHHaMklAlQmPyC0VvfFtTLUFKxzPPv
XmXcOH6+gJSWBXc7wKtKWxwhfga48NKLnK3uffD8Gw210BrrecG9sxexim7g44UZ
7lMuMZoXRaqd37YuYf1Cpwr00xeV9sQFkgAdNW40RMvN58vvmoAg1YWn7AoGPRJs
GemK/JhFTAkaTSVelhjG5I7F6MLakjMyzH+RlGVAoTHeeHmQkxvcfGX/ckbnPQ29
OSo33rUPF8L62jV9hiPC7HWqBfVunvyXFFAX5wMsE/oRgC/zGWaWmqfs8UCvuLdc
EFN6mDeB/a30DrPP6vLB9zkpvZ0iN+m3Z0pllB9wUagxFPPmUQr6AghLYhW982Ia
puTvDiQP/QrHHySzxq5BLqCQ2520Rx2kg5Oxfeh7iecvDl9holsInm7Ec8/SJVtv
32Qd5d6thA0+Ib1VETKRgV6xxxDN+ggyLEGKTDVA2u19euQoSTcFLgQzg4ByRQNW
J/S24pQmpGrSXoCfa2W2ADGM2hl3hNF8XxTQduSrtRRunI70vyY8EFm3M90uQ5FK
BXM5nocKyWbSZzEDoYt7nMsrix4Marjm2nX6NqvOpdEywLKa56JdJas+VvbvvtXZ
DQSPJ9/5S+y8+d31ke1eazP8TqeafTfoj8TldYuEvJdoeyCtHlzmAOH0Z43Uwvak
/7nBeHaH5Nk+8cRh6fiefvfDlDCciC4q0tS2oNdd/p36hIfHAbSUp20c717k7hmr
Llwyp010lZZ8sKDcSv4qxp4j4xV8Jx5ZuUeA/l+DzXMgOddaPTt/LZdL171c49X7
sp4Xk4cK0KwipWtfH7ruaPWXbL7+S/ho1Seak0P+L7fmG9AlPRb7sSZuGjI2ADWP
RP9eLiptgcNZF/1/H9J3HXPF7HMshd5mAnHvF1WRT+4kzjf+5PneXm8+v5MpEwM/
7iEqq4AHePS1hlFO6LAm4tVw6MB0nCoEKzKOXPFG38GvOFu56xjz0eIP4Toi6yr/
ZruV8jwEfdnUaFf/vTkKab5TBVatmJhe5+QhwYjxNgQ20r/dokJ/zjT5daS/tiO0
J0zvf8+oo73H9wHDFrPM+1FMRLFv0S1lCBEgDG31Rx2V/QK6AKxr5OHcwsAp2nYx
ODTyWCqD0duewPkghPPD8RsN3iduDYxg6OMIrqDtQ9aaSKNRTTO7SdgYbVXFwG/O
jss0bXQDrlyu0nODEJAmAQH4vrjsSGfNypQY/cqsz9BlSUvJyXml6hBPdFrO5f0B
24hUeat2ywF5MNwR8PnKcq/KNg5+u5x06ILCs7YkMGchPJUUpVlaPnvXayvtmGcq
EafqiTMYYNIVhqrAfTtLAVBsBQSVurSbRwhw+jCcFpYjrYUVhJjOz2xHAmOCZDrJ
Dyi8T7qi6uSTEagzAFmdu7gXFS+rG266tTvz2o1MRE4qPQV1Qkae2YVolnB2QQl4
jzbDcf/5CLGFCNPXbRkuz2BCe7sEXxXvL81MDm2k/E2YkjKVmx5Kz8S18HKR3TAZ
yIaQYMTMEdxqH+shT3LUdgXvHnDd9ua8qRkfyQ68gaOPx2lOEN/038l8uANyNAnw
adWae48WYagnqb6npq2GKOjl69Ke6GTGSkS+TXTxAQ6Ff/Xps0MyKhTPSrnKwpV6
+W4AESRxNt6z/ETbrXbVdM/oUSmGJsoy/aUY4qlB3XHQsDqCLww+x9747Mmet5ck
9SUTqhUsDfOslSZd+DhJYIiepB1As1t6Xc8FZvzal1ynkns9FKy75Xg5DmMkhOUs
DWHCwOGviPywWPIAZOYXYNb1u4duGwq9mxmaSb6hyEVWFvo6WZLorWqBWOxY5UUe
nOmldj8TcK2kEGA5qP5AbkbBLr/pQkmLxUBJV9nIHT2a8n+v/EXTiaDsyYcQMrMF
nsCHms7w/oE6kYuz1fGWFYxZXS8Lq8Z14KeS2r62rVQipcCrgopAH3MqLPfIeYn5
fvNXI7bdalWLkxkBQM5t3dr+NcIGeaND8oNEpF1APUteUQMi6xPXs21djWqa3G2y
r5zSx8+J0TxSzHdTQq0WAxhHGysE0UwCkd5SdKMPLWZcHhMJRLWhKrdhBs4p8u3u
bnBMlKb39yelZyER8E2OOkDiQlEIHlLcskf3fM31B0gO/cVPU7TS6U0qOMz4tMMs
BOyhHZ1JGjfyf/5nZs0M2Idd1lygK2juFKJzHAl+IlQHobxJiGW7Dzry/ByhK4yA
e9oxmFrA89DH59enjyvhnCnLO43RzY/6W49dFh9+mC8Bwx65VpKO7SULISKZTvpi
NGfWwB35fziLqgw3lmLVPX9/QfmMyndaz8+/AzBUgsRxxJiVdu3ShvPxYya+O2om
qlGuLwbCxc3+Ti0G966P4wPn3julVHaYLH2hHyjBYl3aEOpJKC+wXYmoYMrKQRa2
uk2tICXzWe95MNoBj2LOF3MW75B6mt/UMNlgP06wuw41hDW/KYW4si9MfHllstF+
jtax4rKwe0lNKgUA+XAXMyFgpyOGSfVHBvBcOX9U7M2c9Dj3Z/JOe4TWDLOos/J/
wsyZlWao9Etf9tuTN27e3pm+4lUUejTyjab7hIXYSO1zbY0+9oPzEtLqUUWmdyYT
S0YJabCzQHL2dhsFrfa0KruoXV9caCe8R3gB3PNIVZOZOAmXD7vKpQvbAYWgduEw
yJN7ngx90NmqcxYaM8VBvlYyRt1lRs39AVoPTA2gwr9YSTVVQLm9D8bk1fP8Zxe3
lQhteObnUcWfeESyZkkCKb0zLbYHdTH2g1EKfEUYSwKd2o7LdSaJXNlQfmI/MLkr
XAbqkXekfHdL/PZ8pvPxfs3lT7BOPmHOMmIeQrTU3BmyGD8LWmEoz6jVGtnJzGOD
FmMmqzgY+vSLFcBq9gw/JAm+06oveiw6P0cOVcsSvUJ1ZIjMRfFe5ZuOkVVm+SJ0
0vqbaw9VBqeKGBAl86KKbMwBFL8nMspej1mGmsXQquCZpaFFor5PGHMnWAVxaTPu
evSY1L2FiSImSvwUNVi4c7yuKUyQnEpRvbkdZ6+lpoBjr/FeYOuSZyoKHJ69+5Zn
u4lJB/bbSdhH5JFxnT+KpZbkDfdv5Ie3b3pTOjGndeA1zhie0j7j+eZ5fIWBG3fo
y8SpikP9/5TAnNvG77M/7YeZuYqNni55R5FPBbvOnWvlvM8UijpxZrD0ytpSMf1g
7UEe8oyNAJL37Q2gERMMWyRVKwtXu/d30/iuLcOcPweulvDBNCDTL3jnajHIc3iO
yrLbjOFLOxP59K4V5Mu2/aQTkBzdze8s95d0XuhO5lBoF8p9MsSwfoxYMSJOYqBl
+mkWQi4/1ElkhAkZd8gJqRvmVQteMoMq37KLKofiCBNeaeKQhVJTQcC6R17+aIBD
OgeTv4FBHOYQDwkNTReuBvMV/2uxqSB/JUC9OawA21AFsWFGys39mWO9qMOCB4P3
+RbzC+B2eC1j1aGRDyTkATKqUcfwphonAa0YW1wHuNZtwjBqZHllwpSZwryewfjh
e+XaQ8qX7bFPzN9oZii8S3QJnB6jYUwuh23hlhDZPGqhr7fUqtBUHarAS7YHCf+I
mPnn/qAxa9uPLhTHt2EgbQv/82fxEsIsZZrQ3AeTQgac4TlMA71BAigtGPsjop/l
c6V/mZprBHmzcXLtJgUH8Zp0fmRoOHUxAz2jjo0PfgRcZ23/N3N6/GSGzsxymRHD
8Twt982itrNf6rPlEbyKgjlGwbS2VQqW4rjm9aMiwmt2NxulXZxSzoOQK0cqVcj5
UBKVjRsNakMKL1TQKGjzZCgv/sEKZkL+VZbdkUpnuC2mNwfS4aOvYR9oWMT2B/80
nJjrNTp08zAa04yqB5m2H8t7zaxXrCuMMORAqTKDD662vY/CYfYKtVJXsUwBU4uU
w+jMLXimQ74hoPgm3DDzh2YkXcK+S0KbY+WQcJPGb1Yc9jQ//Va6BHqUli+PpBts
/CHksnoFlE06CXCVEK3TSo66+x3uDsh4lg5mh5JSFYmIRPBjTbQMzT8fH+DflvG7
sKFc55tBRZUKXtGgyzoizzVxTdvO7oQZj+1ZI0h1kbFI+9P9DNKq+jfcgNBC/yBE
ewLeMGZQp+L1V24thBRkdZjIZF2CEDp8XRftI9U7xShsBOEfv4SzlpmlCLOuFYxd
aCGl6uiceHzNv5EbmWZrE/eMFnVBL3jZPZVg2PLZW7W/kHzQdqWs5nzIjPwaSVVm
lcAKikhUiNBYWp/R6KZ4i8pqclyedbFgDBhx04TTP5h8AqwnHElqA1s6rgHGryjm
HB3LfhAnUI104oubEGcDlcu75qsb15dIOiwUbWenob24YDseIitPzfCqbfiV7Pz4
2x7jyj57j6hiLRUJ+09I7cpilfQUaTLg1mz4wHbJ01ACH/wxf+woaHa0TBX5Mwd1
+/5FW3ZCAoiRRO3plUnTvicGfr5yAChrmNWagyBBkxpPBFcYAwrzEerAczPVwSAd
NJwUMED3EOUBplj+VBg2JqU+F+4d9FbN25BqoAGlQABPMhUzGTqqZbQI+uka/h1r
omOBF9SoN7kN2oUelF/B+RLGtsA+YAIsZeG2aoknSF6rqHwP7YTNGkUMYPLUhoeQ
8Cf9vZSuG7QCpx3f3Ia8Ck4d1U934ldRFN5KtDNwLjBMbI27ZLyrtMH/pfVinMvi
/1+M6P4G41nm1bNTHmAUPUK20zhiXGLeeTxwFphcEJsH+Wd9ZBQ/IgTl7hQ2FD9I
fZuZdwLWi2cMCs0BgoKqm24u27eK8YIvTQ9aFKqvdoRuH9lgMtRlj4EafkNNYAy+
d8duz/A33CU3ntyFjxYH0DejtDviCY4WsGDRHzzCNXuTiBlTaOm2Clt7Ge9yxzmR
LTaXLveqFotV0iBPkF2VjUjt0aot54m3DIK1vIW2y6sA/4nc8JyK/hsU8F8UBopg
mvrXnJE3lF68OnI2a7SBQekeJblKe1W8tgrkfbJWR8oQBqi148LVH+UB23g+6yUd
cVDBRIfiF148c4p2wz9v1SCd4jUjTxZ/a/LOYb4gxBmx6CI/oVyXu50wOX3Elt9V
TtZIagmLmvfIKFPbj2sxE+nMSKpZgoqxOgFCzzThY+JhDZcqVzFtugnaGu0zGLuc
Xnn2xU+p56Zp1f+sPKSC6p/CbN9zC0LHKCl94F2MuxNIaA0sG51JqH3iABP0PWB/
RoRCNrS8UUCA1ObKOeXLVR92QBF+rwICJgp8oiVB9qtYS2YF55tb1La73X1aGBw9
vXMitsqB03OJiVfnj9L8uvmp8PDh3Jqn37Bb/JhnhAuRI2P5OOTz9siBvu54+L/F
fPLFESFUL2WUfO7c+hVoSww8BttFee9SoOiqXA+M85ij/a2vv8PtXHHgQnEU8yls
lbphix0hZv5nuPfEKVBWvmBrGys0mWj9GyVxMaXZrXzkTlawrTpL8ri9y5djWl9f
flNrs8KhJI7cT314vv4IZdWkEFwF3YlT+f4eCg5rXe3dYyiiyup/ByVGgtcpZMed
ddXMAyWS2l3OJdvEymJtKGSFrjGxkqkl9v44w72R4Uko+WIkmWXA8GvoLy81B7vE
rbdZWPcOS7ImWOufbHHIiRg+qiEwQWfrhI43aG4zq/aiSrnIoxkR/EHVpLpvcG2r
a/TvQ0VbkqbLVVaBvSHFbL98+Q3gZM1Q2v5n6g2RXREVAYoG2BdU6JftU0aeB7C8
GTnJW8m6oNqVRWYWJorKLJ/iTu6KxcUEGMiYq0squ4RL7YnKjQ8kzBrQaIYNkw5l
eTn5rCQdWNJfO0FxjOHrGEvrVTuYJooGlOAvXxeZ2+QsSRrib/6bRmTQB53hi9Ho
Y9o3AFkE1r4tMkJmD0TCCClk6aI0n3JiVN3Cl1EeAAlxmCe7GDcMgEaJNjW4EYA5
ctHPrhk2EqM/Zue9wXBmErWLxWJskpWQav9JwMCM3LQPjhSpq59TH1WQeERqW20E
nAIcufbPeC67ghmh/rKuorsmRJGK5aacn3xX+kDvU7OUMvd3i1eORaOR8y0X5XBj
7AG89EDjygI7Mwd0WfIv49YZTIC+qa/qROup/ojOfjYGmsJmioSWWcWGiLpG3yc9
QDfhqxrrimfiK3K9l53XAyyEeaWtSCggoFG6m6ytx3ZcpOMavXFR3/tRK3RkCqwE
4M5Q4Yu2SF+Xu4JE5Bd4lLpZPW0UXbjtWhcCV81U3O0jZ1NUtBHpz96V1ogJoZ4N
AIVoF+w19rCtJc3STfI70h3ilS1PSd+TWUiuICwhK8R0SmNXDCrzkyaHHsJ4B/px
fz4Yr25OLsVOMQ9MQKwFIpRj74YFuStZQGc1B4P580KcuaviBrfcb3rEjxQTZTAd
nL9ojL9N0XmbH0iJPV2t+hfoMtS0Y+FQ+I5yCgZ4AP4UpH99qk/I1NrC0aOGASAH
3hw8LSoBG27mnyxZKkbEDqqHvtuiGI3ruRbYb3+L//Ag+GUW27wX6r+4WANUpA7i
mBE7gHHOaF1dZG0E9fbzl0eSEaTSChg4ni2jO0BeHXG4VLDla6ze7wDCEM2EBtAZ
ETGBf/CnDl6miOTY9BrJgujxj3srkLZgr4KIA6rrDdwsF9ENvhr+y1kkpx5P7VP+
uI7ujMm4vd9UPIXXafpQmD2va5jmxl3ltlEUxrmGM2Bak5lLPNJGja4M1cA/Rdkb
uaa/udf96fn/bBrljy0HDutijU0GWPMMO526QyXFDrTwe2NghtzX3XTpPV2xRbSB
s5uwgfAMnCmow6BesnzKcpEdfHhHf8oOxeYIXzkSlU2RvBaHkjy6k5vcfw/0y/Tr
DVgZ12nuXBwEziKGY6vHT8d+W+rFaPwe3f3TyJTUGjB0teA2z5Wv2WtAPOZgh21W
TAZMoL3tZ+qTjCzXO13ZcxmSG0f9yB90Yt2q8VqGj+FLTGhV+Htjfikn6QgQ52Dm
qkJUqW0RJW7zzQXBpm+qd4ogyVj7s5HByzP8vuBv8yH411yjLQkk5y2HeEnggYtt
3aUOSdBnIJTLF2mXak/1njxTjiDcgqf2TJRYqW3eAlmjBaR5b5WgeAj7Ub6lu33K
nveQ/KSwKCntNaZ/Td0Mi7tH+EfrfUr+MxjfQ9OpQHg/PjgMatVBMOj1ja9uX5dV
zSMkWP8PmdVoTJOcK3rnyLQlrbqvw5TICxTQifZ3PC7DdXsT9SJXEQHvsjkIbv2A
bapoduu5s34bSfb4MBbH4mdQMGN3OWoSa5dpYeJzqy06bFUyn7MU2JxKQhIo9lyS
VvZ4S6YrnzscoXFYVtwpKS1kBXcNGozHzOTkfAd30qn+/Uh7twKjhphZv+rKLF7K
Za9ajsVl7RatfpsFXUAvzMCOVQWwVW7w1QOdWe0odxqe5QPQEoEdL2V3E/NFgaZD
XKz66Dfi8bAIQO5qM0X3LfCX1hDTLzEZCx1ebWyAfjZdESoH8+MrdmdlLkylBEh+
pdEROczvCPmOFV5fBtrBkHfhNqX+ZQH9xiCwglvz1v9Nc4E47EjBcELglaajG4fZ
MgBIovEBIOnWcXslH3mRelK/TtFnCg4gNVUHmc2fC1wQKx5b+N4/8Rr9D1P45+6v
JTwpqoSOY82781lZRMYQHyqP9tbsO13KrgWJMrrB7j4mISd2EpaUE6Huv9/i4OCM
iz87pJu7LdrVR+rN9mqEPRdRGz9/9HZ2xEBOR3ERWgrCibJPCV4qpu7w38YN/shi
yvKZufePeuZhGQOq1fml3uFyCMsaVaAW3/G5iBNbJD0+cXOe9J+9UVf/8MszU1C8
S2ai+o+Sp43AoXhF6yodI9zgzESfGD3fpVKzRGM11M7fPGs2R9n7CvzCnppv5S4I
cYfZGKVsM+zfPZ3NFvGGsgbf3OCL0nwN0sm/1Ur2JCMF4z7/4iW9iN9fyT5LUke8
NSYfEw6Fky1+nA06XeI5ab5rV8E90xUIkx9GrebBfbjtq0NNBo8keKXy8rbWOviM
DZhPL7p0u8v3z0kf9zwjrdwr1oRyW/fIxzBCLfwWPbd+bAEnBwTyNeJ0CerKIFGR
n5pO6UuEUamsEUPrF1YYM58TEJlz7v8uVrqC3y6C3jNnRSKRzd3peKgsqJk7YKL8
e25qIrZ0nqprArZYu7NFTyasI98+fW0GXCjGx3jCtLK+kFIO9M6lH5GDAe1kOkUg
qWHJ5osBzi7wT7EqFoFOAKM2yvzzgoMkFLvaIW0M0f9qrdxlnkVUQnYANHcasR4W
Gh+JgHB2znpwMlxc44zIru+2JUpdwE2bD4B1cZBZrQRtI4owonFOzyjM76YqEx4f
ZT0tGWgqNmSMeNu//+3UEoTOSwmdUDQ2/7UBJqmI1zagoTRru6sf1tx7hVJswGbd
Yj0ffE1I4xGxCbjtfElkuUJMbZVWHPTU68F/sdexBE0gvf/zK2hcFA5yQEXygp0E
pTAI8eds00Us+/jmsZtj/cEJeCXJj2VEdTYJz908lEUkDDafES9HG8s4R6Hq/NCF
V1gQ9qPMq/gkqb3EFUbUTVSPa0QHi5nAN2mjP9e8SzcMrLKJKfjg1QJTrEwaZ7wa
igUPsGQwbACt3o7Jv+qkyT8iOAu/gZ45R09EcUQIXafw/OcadpNli7Ata+F2m4b5
lMpv6rARZ6ZXuFu9d5hPgfvF6/Rhjdk0nxY9MJJcmsKAPNzG8CD8ekb7b2lOSxof
tjEhSmqfKArf3YMBEqJ/wIe5epBEPcGblPbDGCfZY5MHNoOAYpJrWDhl0Re/Upv6
/t6aj3R+LBF3XrhCqhuuQRaXOtGgtk9iB1vnNiYFh8NKKyQ9aLu+/IBJpcHed67P
n8egJXJ4QJ8bJV0s7kSNvFQFeBlxtOZyrSHbR/YRjiacKJ2Xx4dbHYVcHlv6LYkc
fRuwJE5vQG9KVTBLXupdi7cGUI5y0inuk2yxDzIa3Tm00MpDrPI930N6HcNYLbdh
OVjnln+P7jWWttMTmV8x4auZV5mToQcHQ1xmKzJM17JAFGsP/SFXr/7R1HO5piyO
uOVemcqvX3HMa7TBcy6A2b7C63/oL4oVbokgLkiM/hEUaHrfmHZhnUJEiGYBIXVH
0Kkg1vHmLvFhI9zn6iV1KTxRFTNdclw4RjwaqhYSU+YZXR0jLqDLi0MucIVYoxIU
K6upQxE7wj0EwRGlbCst1Y5+cUEUO+s3IcYIsmMD1rC8v9wslHIsc2Q/ab13DsVp
Ds4BBEjKsxNrFo8Mozirc/omRjuDGEqWelXGac4qVRzTbXdXZJChwYNW9D6HYklp
UxqCHk5fk8C3KARbYtZljKIwY8GujMhTX/sHuep4fAqj6gvZdYZVuTh+m7QsRYeM
3D8BbmrBn6jn21NWTNxZOi4yAVOWafkuRdVfO8GFahJzWs+h3SVqMYm4qArqCayd
l+ZNCrgPnNtrlVRkVp3lYUn36ZXxy6Sw1aK0I1xqiInAj6HfHWQXQvLqWy950K7Y
UHYc7hl+67+8yq6R5Yn4NOiCtTn42A9OhCOwerruV/mpVGq1Q2FXlLdS28eXxmpW
/YYuIm6Ls4iZ9K6l2iHytgJL7uMqAdVGz+/jawRiQN8V0L92/ktycE0srHrC3aJM
Gr/RNGrclQ+7pQ3ddS+neDno8wcjkJmnmUbckgLo7ymkDQGjZO+hmpLpONtYIrHg
/qcjtB09SQvpmEoHWwBkSKB67mX8TLGGEuyUVvZXRgd7PC+VrbVvJnd/tT0Osolr
XjxxLlzMbDn0pJmvTX8aBF3v7c5AIDqTGrHNtsangxa9mDylPd1crs7sxNPbnytL
vUpDUpt7/K7+9w6z9Or0MPSEwf9sY9nZ7k+XnDqpETuFA4d8oJW/st/BGWJr2qM7
+xaPX41nvmUldRlEvalX3l4ARUHaKAxtKdT5FzVkj+R1F+7y8PlpxJPbW0vUdfc4
KrvPnX/zLQ5wsQqEd5PKVd4K92ecpSR1cuxPE63D+yj+WnOW0GQOT5PccbevQKSE
RQPmcPEDFfkLenBXQYB3kyfUPz/btXQpxbUz8p5aYCQIfgItywWaPcjVFM21YR9e
+KDK5bIXf6HVUMcNXFFnIoupfctR0Otibazd1N0hjtDgxFOBlFEAmNKk+sSbBh8+
lGz9bUz5o4VPLmCtGCyDHxyhcwFW0PPVYnP47vZs/oLgpZFfE99HpYb7ln4I55oA
rgbIVmZNlHZB6HLRIPGUMD66uCB6zX5nu4VIMLddW/7yimiy17HRc+rSBqJknVRZ
XHDMWal9vAO20LRhLXHJLAc32zhM1eTSjdA3NcHg4+8/sbpdn80/2x7BvLxVUB/Q
qhnfaxE6ScJomm6/e5ksHG1fOBMTPDUQhsQN47Sp49fSoTCsJkBFgxbLBDK6xZHq
mux4DLQKmPXHJv0dNLH8ObCtKIp+acszRpVe1NmDCQc6yRw8yZzd4sOQzvEkuUim
mMd2OS1D2xeaVezya8r/wS5W67TLxF0dlZCznPfUmrQVYtvLhy4wr/ZfxFMpFiEJ
3suFrJ7YvXnKp1A3qJVMuEIQvKCMSqtVdZBF6Fxq4SWIdv9vgeDQAL/ypTNQPsWr
A+oXtl1AyroJ6WJg2I8yy3z5a04uZKB+BBEGS/vAahPlCC1uhvc7S7GbXEeQsSZ1
Go7HDwV/5cRvY853VzuIABarvvyOMVtgLnnQjKdDU3M4wHOAvF4IER+4NQmhWgPo
PW3zVNyFOUTd6TyGXngD4+RY8iRu3QEYy/AUmFcstR8BXae9Ef8PdXC0g3Uz6A22
3rjUiC42GeanLtkR/b8aTTfyF6GirVY24SYro2RR/EkQU97ZyRqoNYJuoZ2Vs/ht
wNx9xVdR0ohzOmCRD6lOfuaUsrngo59rVnUW4j6zSFltJ9V+VAa21mtuHESKLPfo
coRUXb87LWopsbf49Wp6PrCAnBJY9jjS1z7F4jWyXye2pswpU2RcCbnnt7aRUnuf
6dAb6kdRK6BKl28qNEpN9mNg2rub5avgLCKHcTFo/A01vtpPsxjLH8qXBOo0e1tY
GtK7Q4iVO4ZqxKUX0oIoghBZxjW7NbCBirk/XfGg2HWXd/04QLVQ71F5CNMXaEvD
E9HdCOEaYvko3CwpIIkFOXYiBXvbX0KtfrUpXgJUmA+daIychB4xlIWDHXvPqzp/
BVSqEvMbjc4x9rGEU+vbzeXo6YVPrAvZsqo2Rd7Ne2HtUyeQ9OSeoRA3rqMbj405
mmQ+6ZniZ+UC9v+kWfYE/i02YoKxnQl1FxWhFo0t6vjjog1cMyW7RBfssTV0UtIS
8bwasDFyvA6dkfS5zag/P5g9ryEJbhQmA8xd5972GD5XRsv+I++2CH64u5Rg4doF
Y+Be91FL5v4D2GIwH2jRgU+6o5w7VAsuXxNNJJc1d/CqWnvllWdJ7kcVlEivQY6/
D14nB54V1utfa94k1SCXvotKHpD9PYZZ06N3QX2K+qRfM1E+JL3CztW9DyUuYusy
tW1MXi6akoUMDrgVclAzrZehxF7+dC0LKVHkBexG8KHGcjJ07djO+25TXpJos2dS
/9eZpNDLKwQ5PEdGwD+HghUvLyzIti6NjAMpC6Q1yazsAMtOCQJ3a0da61tbCqAN
0TgZLdoID/qSACyTPLbKJLOB0X1UXM/XyDAHiD2YFMQg3e0/otkvO1hGf8O7/aVs
3X/wTL7NP8/k59BJcX9V5UQXq+HfJJg/43Y5oYAQHRwuuuy0YB5tfxJqtt/qj9wm
AVkr4FfdxaExaJgo5fIDar8JtFu0jian4hsn3XC52jQh/koGSjYz1/fsnh0mi1F+
sKOkF2buU1hKABb94wS+KWolibFBh4o37qqpoIf6unaZzwfkZ5PM7ADpYIoOWW/p
W1CJp/W4fgdnGqL/QYdZUuypoZGb/JWDmAX1E3CDFgmf1WRjzCVCDOveyRW5UTzG
kmF+limi3fUQ9JfPpruSS6PlnVcQgTI4fSmsxrgYwIiKYFLrG4LUn8EV8TsROrZg
Pp92RZsHMDSwDTJsKeLQA71yFb1ehVbWtGmdcXZAk5ps734sluHeRLKVrCQAU6f2
DV7o4Vz7YQqllMPVaDh5u+D4ur2D7FbyaYsiiPNrJn1RfZmX1Tc38EEqVZ2euHjF
ieZrFOh4KgnF4MQdLqVeq3P/rWWcLmiE8/7B7MpTe9mw5d7LzFiv5DfJZnY+zmUY
JFVj1x8V6sYvK+7pBjtlC19CjQQm6vOpaUtksYZdjUt/+2iDkctaNWnPyUJaxdjf
PoyUOa8Pf73LOWQMHAaWA1q8fVnuNYlwD/BWqOseQ4EYmrGNWxAy4tAmhwDEZaaM
BSNi5xd2dHe1WzvL3nlC/BCpYWH2/2HHdFUejpqSBYRo4/Ljwdr2Iibs5YTZcsB7
xwgVJyQ4Efc5J4GicZTZCo/6LpMcWuKkQSLruhq3Oojrak6TfGK5YCkp/87+VAWW
ssDTJrHzUN4uOFQfNvA4de6VATQMNLWLk33ZUY/yMfXIfcvdZuYVtoTMqV53rflA
XO08hV+I27U8xJiQ5Zx6nXUWwAXRYdIunoh9JuR6lHKX8ZJi3gpK2fRbTmthJYLk
r8IjO8+EGK8DarBf9trNFp8QzI6kE+VZXq1XBDrf2Eb7kM4xHlpd2U1IUGCwz1rg
`pragma protect end_protected
