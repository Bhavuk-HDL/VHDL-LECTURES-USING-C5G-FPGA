// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:38:59 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
GC72GqNyXlpA4X/DAisGqNUMoG6oMFZ9RtHPtfIw5ic44nuS8aPwtzzkRs96VBhC
qdBl3JmLhgCHUDkKrCOyRw4Z9ZdwP8+KzQhH73TxWPRoJePfK/8xrTNY3NQpyiHy
Pr4qY/yTBpqyAO57QFeEKd8o8gayXcWLpKVFAojm3uU=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7312)
N+9CuUsvUYCyJUKLvtGXSNDzCvwTz9450kA25SZbnnIb97cDyWOh3O9BFkCqyQK9
3NaWGqqj3GtfyWzYA+1RRPIWiwhyW+WrgWgiQOBy9vMpvODYBmpINZCUD/4sY/Ib
N/dvYVw4vkTZci8Sjzb+ugYNOKIZ1wA5WAjId6INb0ftpS8q1yPx1lbegepfm9l2
gi2QO6RFxwFBLm5rNTMK6CVpidJ0eZGt4xA0s24k/H0xbpNhTsUBVCQbr/zpKIlq
6rUdukx07PovwhukH65T+JkAAjOHgTToiwZFT5QnSWEYRWQUzl5Pa+yQcc3dV030
JCNoxhCnrUVbAoGTmsLR+jGOImqB72Jt8ZcSRcrJaKzqFbc5dTUAap4nFvxunqlF
JDa/+bymY2uRV8dca6rOPdOVVEm6CAfR8URu9RXwMz1h3uMgp6T3FrF3p/UVKMRD
2OpYBGnMLU5qHMu6Xc7TQok/0zMUO/MnYx3ah/XqOzZkpmj/dOoZWFtABwwN2L35
n4uE0TOXrsCL1JO9foikmoeyd9Ds4wM3UciKemkW7UcW9/TRd1fYM2866GUPtM6Y
glU29TP8GYG++qOgmluPOgQh1uNtDc5bm609vjV72RELCOKkdUMgdeVJQIy9uI25
ILTK+gIWZ5/XgfJHvEMhWsgnxF/ud4jJWCLk4xi6gi5HDHiCwUrkpM7Hz4CpQIAf
IAngJwx97VVuWw/g/T6DFkszpCBuK3G721AC/YWstgAwP4wf3QZhhLgv8fC70/vV
pvMlszyQ2KQ8YHWYAXHJgldh2jvtgOCTcH5JcCQnBohpKb2JF/GAXsvrvx5BoLmn
6dzYQbI7DQd3/9/segPWsHAyG9H4EixtMOwlO0CpU1bqvXaootGuLsawhdz1ABL7
2VF5MjmuW2GpvZNbS/I330wpsUOa/GVv8dCHyk9kNZScXp07RoaiDiJLT1iXrjYn
i0xgp2OlYbTjAra/4GidfaAVnHZNsnEfftUQLg+GBZak5J8eFHf4S38LavPUSjs7
4yL1czzOWClPRfNceyXpR19/0zyLVPWvCrMKL4jwoGwHXSx+Yxmh254gqsNWtktQ
dsddjE93F/qYGuDzMgoJM3OGmQPvxaGlb31oprBb2EqCAmLuMLoWakEpc6zdQ/9w
KZ1aA25VoyasrUbT8wr6Qagvl15ihXlQXvjR3pV1dM7w/hAt8v8+em6jTGPveRH1
BRD1ArTT20u/yH1YV0ucpCxQ1yMZMXpdolFOSqG4krAY3eA3DeF5WoSI89dK5+CE
a7e3l9wJYIV5b2hH5qySggbCnPki1EDNNUP3ts4mcH5VQ1f08riAZ64jhspuPeDz
ucglp8iM3couMDRQQF2QOypAytytquiXjMQKsNOzOSwtRkyDL0p8ejJgW/5AwcfY
s0MzAONrI2+WA6hdvw3/I0JcdpxauKdn+XR9UwDF2IntkJnfjsLpY4Z+f4/jGkel
8K39RY+BJJXplDFR2WfS2Tf+h9t1ExAje2Hp2XtSxC1yIH04dxpa9FyQy/2F1iyg
LBkxyp4s51dsxpvTIvV04VVMl/lq2ORrfv/Q0wmS9UHuyGuxsEF7FBsFEdOJ3rec
FrN5Sf+ZI+dpgxBXNTp7/eCWAYpcB+K1m/PVhikLEZvF4c/k0NMS0tKtYdcYIQxf
oBTT0pe0u0k79l/fdSZVBBqLWaKcsfZKI3lTGV0RxyarUQSzoQhG97uCg0LX/i7b
P4fr/nlUMyvkOzfZh2NEcmv0V0BW7vZcwb02OEhB01ZrJGdqGv0VkXRZLXeIgogS
G8cT1Sgf+bSMezQvtKhS6YDX4WbtFxPbRCIUK1s4l8TH6y9iS2M1qewynbjbyjp4
05sBCGnMgZL6P4wl4uC2bRrYweZCR7COh/u6hcgFRcM7C+/9t7B35/4MBylWi2i3
wPJjlpH+eAW6a8WWPa8D/x7RX3tKtQttd7ViExZNwhfpuq/0pmAMC6hXxMysNzXd
Q8wr4+z0WeprdajXVXdacbwqU9Rjb7tCXVkyAx6sohi5MFnh9lN25u34XlpQoCwV
N4Ny4PWQMcQNWudsM14Pm3qboKjuRKKJtBpB3v25JKrE+PtQkd/jJI+P+GOeyiOt
0pOnYrpsl+TTwrcl7N/D+GCcSCcvc4RqfYJMjWgRDsVRr9B8RYZMaSFwj30iT+1A
pPFcBJwmjqEaAgKbEfxfHAUoRHBG0d4G8dLhA3Xrwo4+V5F5YFDAAJHO1xADMS2G
kmRbM4JrKChQHnCk+KIoI1HJmxhpaUNfAcewHH40jafddPGO+5FR976cme1XR90l
DPSPqVmq0O5O7KqckgO1nkhGt9j7F6/dnaWPA50uYAU4Mho02Yyr0sgZ6uynt5fY
/BJXGDCCeMcKwql0LYgGgtQMUjNmXQhKMXnFkjTQ8JmXUWanUEjPf+au2KiTs5F4
qr/k1TKfZrLjhmRfRbe/lh86U72SbRx9q7YVnWG4gYqwPUBYZIf2zIeZEfFUAuvv
YEBjHVxH04A4qQTbWBUlETapXJ0xsD+CmWpw8HHFyJrnOztAa5dgbPkd1+U0uwpi
UK4ManOfJy2oviZFthZaKOPh6Z14DpcS2e0za027ecVPy7eGbglMzygMSqqS/Rpv
5Zr80K0d09uoeOaxOgbRVQcWZXqUzHLw23cnfaIUYvugp1oyEqBq8xNZN5lR+MlK
jU0MT/A9WtuUjF1x5czcQmXq0kcbGWQuFOY2eDWGwGVMKQ8NjpZ7Sk3A5yMekQif
lQ4lSSDYfxzNlxUQO9M0mPMOOH6fqgLmioEsxpR62SpQ5nlvNHltQ7WoaQbhS1D/
/XL3nNKeR7+fr/ydZhQANf/eZUxwOktTR2mxMS2WyTssHTOIZXiXMcTWKYYlOcQ/
cbkBHafgKAWLm6jOgs8YtNWqS1OWYae/7MXKamYx9lmDRXnsTieZrFW6lO8ADorx
8Jn1969JoPxNfGqpXZ8LU1PhOPGfx0n/f8UCvbQeNUIG1y7qi1fTRwXcWidNtHry
UAxN6yySWGShq9EpQcB3G2iElT+MZrF6KNjH4IFPs0Fj55gClJs2pQ192jp6SM5g
feekKzC9gtTTQ7DJMI+1okRgYU+DwPHK58exqxmA+kOcDZcBVJNViFrpyIoGG+eb
xw7ttNpzY33u/Bx4v01k0M+UWWXwGJdCb6xI+mn6Vzabj+29M/NEXtnuDCscti6v
uiVeuWZuUYv8fvuXx048z/TYPp1ECMFRXFkqsSnC8bY+UIwx+7/zdYA/vT8UJXBm
2mhxEtTYBTRXo1YJCO9S0M8LNrJS3qId+wpPVDr8ggGFV28n7O7cKcL4ZguRKc2C
3hZadhX7RgyEghfaqf7Pj2qb60+9aDKoCsshnZnkCBJQq+CNfJc1JwXpbHl2phVF
6z4jA8IwL1iMUlIccrRkwoILXZjK5JD5pnrba6ZQ0Z+ecTUseT2MBVpX/BIB0oAh
vRRfJoObcTjuxCru6Mz6WXz16CCSwzeDrlkttpyTQi46Xv6IbqlVH4kaYqPylMgN
/TQEORNSVY6P07JupD0duJjh+05t4EPYFzJ9r1DOVgAWlcbtNX+kc/SofiQGKNcB
5pG/TpxCDXBdIxcgRBwxXat9NFpWrm7z/xg5e+SJiwYt9+uLQRhemKOqpb0DYDpl
bc1m/2TPH/NyQsZXvEMQ0qNhurK9wQxH+SvmthW3eBG5ZtVJkDFDVe09gKWvM82P
17zBxqw7oJ8Uo3n6fGDqHqQs9AR2xdEmRRcSas73lp3lj/LeTckdI7wlAX58thJd
rHQe1nLTxu313R6ljuf2F6idf0uTYxzz11OhxKty1YmUmbTLTHdWYvwESBeDFZ5l
fsOXdaRSTo4ho87O/XuxZ5W1IZ6VICZtXVzTFI91QqRhdioRa9peKqZZEQVmSS4O
YC0IJxCQ/VLPry2W3TMTRWYZaGZDhvmP7Emk6A7ESeZxuSWDOtzG91We+eS1Ejq0
RKn/K0I9iWnyyFz4PSgRI/kRz609IMsI4+eg8Qc4iTFz8ujcbqc2QvztYOzZvPzo
mK33ldnOrAJ6oE/VKNRQf/2PiU2Hrv4+w+CiPf8mBQREtNSTivwlL4NZb7vGK/5r
3aYSQgLeqbgJcya8OvrBgkcdJ45x1WZ9t0UwnEO94PICJSEGgXJBCORaFVa4tkQf
WkTANRU+1BDVaZB/5ejdmbu+1G2qJi1WmV1mKXkG/twKx36uR/tRaaNwnsR0Oxfw
iGS9aknoYYssL+cezFeTA7r3D1t0ROgJWGlMt1wQhsTMkATBT7yG4s+ky2NOUdcs
X/1mTJSLCGt4bKPFWMJxYxR287omq8A9kWxZYC1pXGQSvc3ZfpIksgy8VDFF/wuJ
dT9ASLqVdYwB/kTHlTlWJxS10anPmF2KP2oryzYIakifsIZzkjt2tpdXDlqqrM/M
HehSXJg73zkHtXvBtpO3lDpAPttxMrVfvkDodnk/Cl7NDSwv7I/0iRqtfYANAGuh
QCl4IB6AKG8PQoUq2/ikDnUXjZ9khiA1gnXCYcUIK0TBnMDTon4OSo+BiCYO4cWK
fSdCa6W1IIapefz1Sd6uoQb3wEe7NTvPR/moDYxarCHaOxaRS51L04j1DJqrB+eL
uGTvrhxxk+nbBwJS1mu3YpevvAxHZSwUXEgIzKbAiKYK49FmP3Peb7zkkbZSxGM1
PlmTeUV+pbaC4zBvbRromD7VR30CJfByIsmCsBrcm0wsHJqD2bwMiXmvQw0GFFoB
atZIWw5HeSnkMd+4/BVFc4XxkTxARt4dkgShDfmAeciPnKxBiWG02N24sudKYVof
RMoTNBkPc1xYt0WZaFEmRj00mGaxQmV7pn3MGneQ28jlu4J63JaaiMay5lIfM832
Aa+d1usxuFnc4nP3gADfOyDk7kizjVflZGnNnbEHtqnBKmhbicFdnl2aeK/ScxWv
RdHvOzAJml3jIhVkGtTk3lY1AMciF9Hoa+jzXxctgay39n34WSLdA5qqRH6zZzOP
4BaOE5SMZOkVnOUb9gaCtcWzR4Kc1U5cIy/GsbSlK1MfYWcwGJOtUmR4l61AJStR
qZ1oTUfb+W4KKWdpc27TQ6vx12HklgxKBykg4Gp1rhrC4Hi4JhfeJ0I3NsqxUzc0
inroCM1UihvUQzFxvrfmdqbDmv1G9jGQMexelBVtH7t9OfdQf/kuk4B+Jt9QNFLm
75GCALoP4uYZTxJVRTItS5UZp7BdJjZOGebVYkvzBVdZnX2c6eDdEEmfvoQFrx1L
nD64J6TQ7AXTDgVMNC1J3AZpQiV28X16Bp7vh2z1MHQ3f7dh17H/Chwy1EMZnJGX
vp529jZIYFhSrWK6aksiG+GtsMrBvEq1lnvQWM8ycr0YvzRHTDhHb9yMwAvpyRzX
RTofM71KtbJ1yVdbCL+CkU2kJKu/v2lMDju+CsXV3GFBG0+5X9XbWDebyPTdlKXu
eZLVHj70kIu+PtwjxF5Rzqsq3cvgX/eABdjDFVRF0j9kBMbRR/RTPzFyJf2pI6uV
9ewy3cO1FEb/zKRkZgfBWEdLPch73gHL61CCTpfx+VPAse/N5XdMrwVv0l9m7gEz
YHqdp6EeVAwjNdADz1Iagd3xR4nMwIOeRjxaTzYJ8dgZuUpOehP3DoMcc1YuPF4y
dM8FoFbHreGaJdV/ktHxj7bI14biS3cEu9UwdyYhAol1xR0vvDHHBp6FAL3KPIc2
XCF3idGj6E1R6SuMYf2vSp4ebD7BnnTnutmjPPqiZix5EyuidnXdwV3mZLSayYNz
Z7xWieDXUyV6e92hlsMgl8bVCWrpDH0XrzVpvpcgbdwY8TlCRMNvTuvVkVjv1kbJ
eijVz3Epe8TH0sQ4nGwMnNbLKudMVbSyPijPKS3ACRb1At75XfdfoPNLiTjfVi7D
fshlM3Mx/OYIzACDwBnt34eMv7s2rbkMTef1ZKXJxCFRw1iBdjCJ3pWZHmwdq6eY
eWr0Bd4T0UgbWuCGzNZpveaDvo/edzRWW6bZZYILxQbqqgbTpM3Em2X9J9ymJq16
pD4fyXlbSyiYmE39uyjQG4IDo/L8iYYQYJ+TPmtFW2cXhtuRQB4jGYNZXYpMsAQ1
4XKwtSV9hNJ7p7sPH0p4fxzjUMRvDDkyzfJYR4rJX5/pEYhdLe37aD0KnDGjfnvQ
j5aFbU/cQZxgzB4Hsyw1tflzqlH1MaAy28+eCQtvemu2u9Gds8Xuaxcef2jx1fXX
+89Sd8jNzl++1tY29AZUwBDv65FWABox0qH7l1OaUZtXi2rKKTQQlaaASS28Du3D
/PBHfg/74NC8CEiW6A2h13ewHLNxVe6OeujOMb9FvUnAd4N/rBLL0UITIJrf7oQz
o8t/iaUZburxVW1kZ2n+ZNSoPvu97wV509tqE+29l7BwDydZLEK6wn195+Na5ZZs
mFFypuh9dqyp/ybsQUEgeZhtjUfI572fKezENwFiJ3tCxiJAPJuP9MqErJX/H8YB
TIaLjvgqpn9mdCEP3VtxnQZr/pQERU40YuSr8C3jQmOicARYw7FRW1s0SgEsJxLP
Osw5b08bJ0merpHejtw6JCEwSr/FrTjfkkGgdN5z2M92Vuida4B7bIvImycD7mc3
JaxgyRt9kPS3NFS9IyRMPWFCzqx/z6zU0aKRMALnX/uOda2ftTWxmHX/HmpqdBfi
OYdyIqkTB2pG+NQgswGv4GhGWx0p7+syknwy4zpzUJ+OvHHfPcvg8J42pd/y67F6
gfNoXjNbohIMv0VrC/xOZH9tHqa28IBAb03rjUWtXo3O6/8tRsxxTxfI386aE9TL
plnnxFMDCMqfEWE828RAk7diUzB0nGJJHBgy8XYEIu++MdfxFJiIFMgNZfbJ/h4q
qAqGsph2HCvDMp8X2VQPig4LzJjz9lQ8W8bHuvcQ5TH/OBiOHpETuBmvC1FrkBso
rHHUoaqm1LdocFOxvQ4bEdcbuPRwpxG2gwq5kI+4Nva943ZKW2tutMsuaArBBi6r
H9XsDWJP4cV1J0T2MFNuAkMjLc6LOw59yvqSZjANlW+pSoVwvrsfsTIrVbXeYbJu
lSuwhMy6BMv3DUFUnpKHvSZd7J5nU/inp6TATPTtlRKnF70GI4CkjDYoBCS1OEbt
EK410w/e39VmpSoJmJEBY9dydXebRnjtKE2whkcjqz024uIxVrYVquDe380Hxf8d
lpdNt0A514gft8QG/BremTPcos0GEWYJHu9uiiOF8HviziGpbVc849epSZuHCcj8
DqTSVjgKlgdf/HvEC8WE4NemS5g3+tCv1m0XNCcfiyPMOLaNrm0EI+wfufGolJ0r
dMRQa2+DjBOS987dnUOFq88gweYsqvt3OEsTAdnUAgXMYRcdNHyCPvVyzkp2q39Y
vgvSmrBc2dXLGpw2Eu69zWKAf6nSyPYJrAB4aJNeWMAhRUOAqowl/ng0tl3dR0+J
g0x3/I21EVdp2dZN5obPTyfJCwgYvqI16ctTcrDB2WwbCiNFZKKoCnNVt0pKHo5X
7228hyB2JYp4Ow/tmHq3ogBQnYkn32TRjRrnczT9ZAXRkTO4euiL4N7lhVIwuKV0
xhtEOFrbz/znQ03MoDIEPFCvF8sjdOAHmJD1TnoW6BqR/tBQT4hxrEvDUI3M25RH
v8AseFnbhTjOSWxVT2Ue8gHFI/4Kbw3j8LHIVlI6gEGcwywBXF87PYKlqKDawd1m
VMxTij97PWy46qYyDx/TIPjR++rPkxmMKDMoc5yE9nd7d9/AZl7X13wAhgomlFDd
AV+uMpNyo5tZaaPkfHWsTOSXx212GR/C2jy91FSihiTBMIcwqfCDjxe1UjoceW9v
mPkXGWTBaTRcaeoSPw+ZoyEF5mwsbIF1JTFiFP9+YdUlzR0aDEBff9BurrzGkc93
3WMnMpjjgmzobJj/PZkZSQjDbvcOmKQQA7cLPyc14XkRDTUsvAL5PU0l0bfMuXUy
YyM6yV75KOH2M5Jd2EDQZqHPKY5izGncSHGEcHgpKvvnRgOrz2anYDi7eklnH5yd
+42SjnLWbUHT79TWWy7LbuKlO7GolwVpNb76TtDFajKr23s9i7t8MxpfuyasflhD
NbPr+Y/lHPekjY59mvvIx2nCbEyeRkZtU7VsqW2MP18OF0yfc2tI9kUt3of0t8fc
SNIVFDTubMPbgka3GyUuws1t/Q6cyv7XaZed1VDHoIvI/EUFwr4bDKGpnG18Dk6H
nOl6D0jbjX1CeHFM5qzCpWvZUaC0GbSo717QuseZ8Qn/JNCRDszaKYWO6UZ4n3/e
PsbhM9qWcUwRrDSHRRK7CK1zLOEy956+BURqVbkvf+c9dOUgM5ZKD28f2aoD6LdF
nQIqsue9uk+/0HWQDqhdQUGIl43Ay3r2zoM4eJ1a+6BAVyOQA3ioPhRmM9pI50tS
vefbv4zuvqO6Hubno4bN8A+Hk7DZW9RcPxx1DlIuyCaGysBI7SA5IGuEV5AUBtZu
e4WaizPalrWD1SQCy9jCTRWkj7fUluGf2lHSY0F0Cjd5jgW3fH2gKvaoOSo156vh
3MTxixKURn8qwgxppMe2kSAu8aFNDqRt85weQPC83Tq2nKlNBzg2E3b0Wq2GmQN3
qitOPKDlPfS0awJ02PGJmG2pMTQyfeLe8cOYOPV2njK4Z/NQn6Xd3QtrdRiESoXF
FjvDP2cPrYwVb7TkrhlUS4Bamr+X4wLGxngaQP2iKOqDQgjVcnWu9YzVzXw1ocwR
Og3/NruyoSNvFeYqtwnk34CV1VX04QsJyMPZoR0zdJjHr4YQ3mil7h64o3WjFyak
+JOB02KWxw2R7nemMGgZGvmai6rjIL1tYOzvLLbKXO7++DWjYn4t8X7dQckblD2N
aleMzezW/3lCPP1ptdcI5WclCRS4RjMTtCuITJK2n4Dpv8t9UQTksGIySqL+dA+H
8uEd8IzoXRQrYIAqORJqXxmmZpP2xO+/IIxU3B8/7KCjBgSK8gRnPmQn68ooD/e/
AmSREJgPaTT/7HfOn5yaBf7NWgR0HFNnEdrO8S6foWv/1AMtD5rdTTVAVuI+lgm+
zaiuvUCKrcSxcbEw9zGn8+IYoF27psrBLIX5TiOeCTH/3x67LaZwSF+HOdUYQiZI
ubJ0CERCsTi2a0rjr6MmTRKWjtIOLLQ6+W0XWKFkgpBjloQSuOfOibrWlR2ZEXwb
jaUxbNOwiJ+3uaPMyhjfNM/XsIa62zDiDrjo2A4TGRQOgwEsxR/VTz0ntmIbMPoG
RTpCmF6WVtVaYK2tdzfdPREy0NkSLyK6WC5mmCZKaDSMzKVDki1+Dxuiiw+7d+5b
sruwjDm/bOyPef+jboyb7OKQyDQrWVGFNzWNeOGypMrIMMW7rBbi4Fodi7uceIoE
kHQKFV3vJWx7B6YJAbp7x842OFUf8n+CAxw9oCNK8Q21s9Xv/IdyWef4clHspoWX
ExPoOeaclwoX8fmDXQeDdl9pSxA7NeJ5oOpGQXLsnBi8woBVUKeB8/sL3LCZvkQk
gDl4VMSoKVWKlZJprbvRwS805dedsfKlxLvp+EuGMrYLdSVnWbn7bdEsGmzLXTdi
FBdwv00LnUZ0eYbqcLfC6lvxSnojdsfPJyEHO8eBXwL4pbUUKCvWWVMNcC57NSv1
4YTWJK/GS2GiBKgitiQocD0vkBqcy+3UEUCD5DpU94dveXryv4Ce82P0EqLdGjTA
/Dj2sB6KPzSWQg/t5kR5vkjDyd1nLqS2JWMlOg+moxIOCfZZkTqLEFiHDzfh/Ut5
d4DBfkvVNjdOCYNl3WOw7g==
`pragma protect end_protected
