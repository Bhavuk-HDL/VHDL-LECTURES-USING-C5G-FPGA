// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:39:03 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
kBSdhthCydHuAF/1NEkXEIoQ6SGcmU530qxfM0ekiD+yurivHVwdI3Kq4FVa/mIr
JyKsjwMXaVD/mqFFEw6ZQcXspL40+2BohBnpCi1MfssUItuO2QRLajjfD7zd9wm2
HeoR5a4rRoEF/lC7Y95ZXcS5X1HWKB8+FtRx0SMbmi4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7424)
BLKEvkPEOiN5LEvqrjiRLJn7vXViPoBBoMEQ/tXVe+vwKgQNApTXLbOvwwANf9zx
MstlLBd1YeV14ZdiWe/Qbo6Yffm/OunBpMBfsFmocnUP+zgk4xic4wHlI1KdcmcA
4yjDd3z5wJb4sp1yVabGN+PW+pvKXZHvUJVNPd97TFf4qkXBtwza+tEMd6/WQVnC
p5AaU/LrdOCtNuc07F9qq8m/+iC+baF2mCBmK4jCtXtoPLTkwAk++BspGz7E3iuY
dz7VuDwCZ1HJFKVtFuEgEUFyWpmihYrW8Rdx5rDxNlrXA6HlUAkQK2qmzXVYKrTF
lf8Cl5GUsPb+P6E0ceiCuxz0XIxqpkJThApQltoD64RYVXxUVoyYEhUBOqpg5jwy
UGAB/YrnyQ8Q5tHrtebaKUA5mTZ3FT+PRpl2zZPut0fRu1vXsJkgsg6c9uIzs8Vf
2ejHgSi+Ig2vBFB+hDYy8FNk1OHELqMIEbvdrAnSifD/PMqDfqb8s603Lq7BGrYV
bVqztPM4fAWvZd9R1iePd9GB+Th1uh2wzfWwEcePLPL2qqtATk55C2lMB0ocK6Vy
xD4Wy/hT/q2e+1gE/t1ea5Q3sBozCScjmjZmPp7AraY+WpIldeF7HV1xmtx0I9nD
keFVRVs5u3s8xfWOgIzOgFi7QAQVo4Eq1BHNwgAPYPZ7Ozx4+WzWmjcK+RfGSHgp
8raz+0SguW2sbgln8Jv/7f3x8smO5lIc0TRc/5CANNsjGsj9DbHWDpdBmkEyrKDc
SwK9iiU/pQLacciYsfk1C9X/CrLO1LvoO4ykIJGI757n8cZnmlxZNV0FUJgHZOzh
Cf4rVVT2Z7mS4NKRaAycyEywBObGq8T7ed6XKHM1s20HS/Hp8WRff4F0YRtJoBXh
iscJdgcUie7CoLcY3/72B7944D3O+LXlT2IUmmOGqQj8yk/yy105Q3NWal+n99Oe
LuIwpuHe5/4/BrSeP5HmRCXge7NQ4LJsMbr8Ehtuluru2N9nKrPjBNHk3CYH3Wns
VP5t6USeJFYksNnDSHAyvuyhv/9I71mrVjC+icG6PYWCkMdxgjQLj1UfdzoF21RC
JcpEm1RLhtc3HLEfZheaLU0sZ888ulUhZB5rIsH92Ar6E1Ptnb3dhuYpg9Gbbpb6
J+hqoyxeRjbiKYDvnV1+tt+0Ta9rwJQbKF2UT+gBdopayRWHLVXdwT6NYKkpxNCJ
7RB8aznENn8+M4WcdfNG66JKXtlxGjMMCSGxC9NBprvqNCEVWQtcSW02MU7o0vFi
ZmujpYFWHJJJquU/7xW08ObKt6Userba4QVmDZcUGQww2WlTLhOtDDHK1RPP0Voo
FkxFhwnehhkg6/uz/6IFiLXPktEwP65TWHKGFkdBMCWraCygrznOaCNy4LZ8sFtN
rwvh5TyIZgVbozjuIkgMqEoAJtFOAqoziKsrqbaigouNkT8mA80gsR1Buo3HKgps
aGjFLhCr/yVx2D8tmrqtoUJEw2GmIe8OtfWnWy389NSqzpCOJRogSGcESKgNbBv0
GoIKVSIP4z+6T62iCb9ArSfGJHufSNC8DhaYT76sTJ6c553PLCbFuiWBvQScXwgS
pBKqRDOEjfVPj7wq6TyKdDZlRgKwIqDL0aFhvo3QHoxzSc41qG/lGiMGSjozy6G/
uOkkbpDrLDY5SHZdPcNA9sf6SyVZMyYFWwser/x/CoNaMFgGbwgjPGtCsv2ic7MG
exMZLS+eVmYc0UwIHPYO1cgFCy2oZDKH5cNQT4LP5LVaWuZJ+r3hogMZjLF/yt2U
eJ2fu+mMMk5Emm4jv14PLUjAtq5Mfcmi0AHU3Q5loJctmIvv02zLV2kJHxzVwatD
PG3DwqgoNvEnx3XoFgoSD8tXSXnm1WRV9YkIeiw+MUZ5/HfMe0wVHt9CXuhPvbgU
qDg9NI2b8PGaT/JUxo/RXH35ohtqA/+AM7BMhmu0zBITA39qPnhLxSAb+UO4VAPg
sGvtBMe26OSSu6k1FNWr2dspAIZRkeK5gjQjSDdnEFn69n0z54RfihxBAV7K175v
7VZRNfbZ8uL1OIkedblI+kZTApCx/yx6Hk+EI+nXmLImz58pYcb7pNTVx3hublnH
R2BfM2Hg2eL+Cqd3HLaFqvRnFt7qd5eQKD2MEsdkurwv5yk/0NpYglRT28WN1qOK
6kdvevCr6wYA4hzxyVjiRH/RhaywI3gh6t4FXIO7khMoZdQE6ltHTKXjVye+G0B/
DuC2jZY700OZvuCgfIvn7ezvFm1fE7b/o383utC20SFIiI8+UyuaWSt90IIk3zIg
lBn2n4XTeubSS+sY5n8KD9HhT+k+kBmX18MOJrOW2LAmLssegclupj9oaYk01fcY
lGT0BRPkWYyswczpXEzBhgeXb7MV+wrYOtQhhtPe5LKZ1q0TESISEHdohX0RMrbb
6Xbhg6FkOPUv+OxTU8fSC7aWN30YZibbvg3PRjLxuDvkqmJ9tZM84horbSK50A7g
rTbaVvqVkdaPNgl5gtK8sZhJjVO7Ih068/e0rCXnjZ4d3oN8MSQaflDNKz7NaZCf
Zny8J+tbzPrEHi5pOHRrXEoHGWKdWX6dz+Mb4fHzL5RgLuz5/BaUtuNtAb85FvIX
08+IajwUyzdgthZZ04qiMDZbuDZvggcd4HrD4viTSlSqCSMCGKn5bxRMl/L9gH2k
51OF3fprNB4mv2k99j7OLt8+qftNlar/iM7P3Iu6kbdWMP8SAQgAGVbKsP5P4VIb
I6XSHjoI8KB5bzSqz74ZVGH8TKaR2Dh15W8VIVjW7PA0h+OacjiZZuGVj0zzR3jt
UPjcE1y+9uE+jcBR3xy+lTuU9idrCwn8EVIDhX2xUj7sToGdzT1hDXAsaps3ihj5
CDzcpMYS91zqg9uypkNRGnqhfuMxjzsJDLvv9lbh5ythKMhf5cno5RQtIP5PJeh5
/lSs1Xd8MaUKKKY9jYYN7dqgxtXwnXXLKAYNEktO4C5SKCpQU5RUP4665q4ibIbH
mBpHaypUOaTIigc9ABwH2K/foWWbhnfJ2XNK5T7SZWEH5eWs1bEcSGnKO1JCtVGk
T05Qiy6nb/VHpV3TWWFXrCsWTp7XGRqMKDXDBA6k3dMJPZ2jmuRfRxNA1Dmkt9jC
2yWl8HWmzrjkpaW8+/NMjnGSgJDudWy59aWmdaopBB18Ba9B3gMgHHzuWbcOZmw+
klzzd75R1Wcx730LU9C4DoFOlIy654VDXf8bwF9KYKKXpFluxwmvdkXa0wQJI0l5
4GLGcUVwpFJOJnJf2SbTD+smbDV+azt6INniFiBpCW747ZagA9IxtZjGa08fiB8c
G0+I5Pat9mhRiOh+A/pN0ZMdVSTtGODIGec4+6REdMpNi5e/Oy65ymYuMNJufAT6
NZ0M/Gn/Np6f/Jj7aon2gnT8HeH2dLduEK/gvKTqErNwD7m/pRuwVTdiyLCTfWoM
0PcCSibQJQTA+LUMHHYxRktvB6Rz+jIUfKZ5CyzqeekHLTr1hIDKsTKL70QniMGJ
WaYe/rVl2kNGGrCxcHvKBHhrbYnV5knSPI9wmWaMg6w3WlJRDbwrB45hH+qhW4aA
C4gQAG9Iw672cSp4OMX7wK0qRNF56wr6nPU7OBsF786ngEybVhHk9F773E6UYafO
CDmf54fDlvwRXH3QJ5GfpVQ1Vv2lnMgrepR62tCDaX/yJzGNyGPnNdOGVtNDlaoJ
vbBHt42BiDH6fVBfRtyAoVaHnnwgJdXZCmOUkuGnS8XEm203eEmJX+PgekcLG5fn
xSu1RThzDg4yWUgLfiMtXSBDoMdMbRjxxzyZA883BjMVrKEeOQJDq44zk60EdHYC
7yLIIpMlDjYof/77Ah8mopjDRRhxORCu+MyaQHMJxE5n0HT/TIXMajSK/a1B7w6S
WRlPOxH+Qwd7RNqy3LiBbwX5UNHiduSLrN72oaeGnAQ9DacNyv7f3IcybivVj4PE
EeSdinXyc74aRkpH3r1TyZrI253nNrwCv8Y97Uiu7Km3HAZsybYUtaSzcvx6t/pS
+HfutbNMfSta5NRWScJ435Uu/NYF+pUebbfHtoWOV7z875QTWOFhVYEnrwqc0gXj
BfSVZQM5kcBXJSDheOVwI5grsIVsDeGlJtwn4QAbM+fEpoUnv2GExz0/rwjHgr6W
iIyolAVgfCuRnq75fV6bkG/r988HQJ02YWT4CkJ0W58rcbTd1Dt5+xWlSgeAMmua
zTmz1UZPvo2hge4Nh/CtRBmNbeljLIdTugSHWdXXx4kad4EVHlJd6/j+ZPwI6Pjw
A7rOCNFFoCQwu3Ec9ImVWkAGQixIVv2AJgp5p5TSEXTuyMsNQcOdMj0om2Pbn107
nZbZdbFbcoDUF6h0bGTqFAX+wb7Sez6rNnxFIbY1xUr41TBC/LHH7lMsGAmyV4DV
0Rah/1dh1wgwvGjH9sfv/hhabSYYvufAWgPazN4ZRB9G068nn5RKLw+JNxQMc5pR
d76l8kcut7AtD8ovXIo20LcbeXB/+vv6eeLr1CBWurDhv57b5urIVKK/aq3SEc9u
9a0NMYQrV4bx1PzeUI1HA+cnB0Q8m1zw3alztZR+iHlU9HdwGO2kOhhajOPIohUp
1YQeekXlqHyZy1e9WUzx3uqtfTt0izRq3xcxTNpFuwC84jm+WoZt5iwJeNwwbzXI
K2P+mZdwa2kXJXCGNPuVWsY+Q6kJo2MCT7pSQ5yBAvtfGMNKKLfl30Bj2/Ir2Hxd
I7AG55ld2WsTJgsPQYPbwXGVV81KfQiuvqSh0e4rj2Yj3eFTIPA8uxfOfLgELy8L
4fyHijRmggk2ppiQSMHCLgsMYLELfALSNXV6LWfYSh9hoRDoWUpRM7E00DtPKFSu
BqeB2PNCGp3Zvx1WjMQMhOajhP93wD5DdTwHPvHGuEgdm5CCUD3+dLyO0Z2OOJvz
hXYE0nnriglQ2z88IZiBZ6zZqbMvqWzIxRv7brLJWTr6Sp2MXQ1GqVigjgWSsa3M
MIjWd9NAm+KR2v9kBsoHX5EO/oRv0CDRYvMfNv2LuTbJtVoT4eM0P7nJAwfRvfcr
t2zrI7dM0WTvWjaUEhlD1B6bCMWxoGX+hu3pVO0MIjIYOY4ZKbubGHO+oo9P/zob
pX9uKsz4Fv/hrUmnz5YdCIA+kUC5p4ubFzEWKJripEJEY8V1h+qrT8cqbgzKMBbh
ss0M9xWTOQuCzcAjhlI/QUvHyNnFcEHPqClv6QKdOBXlfS5nBQaOaHw15dm0SqyK
gpoml4lzPyPvII7XO9ylcO4S46Ms0N96RE7DYKuQg9J6vOS+Xx0/PebfRtnBB2uJ
f0g2l5iT8EPr7CsIzK2Nn7ccxyZ/KW2TAv97hFtNF5eQSAK5HAPTghTtDw59lK3D
fOtZHvbBXn1Ol1JSDyYG9EepWGhFNl/wRZOiN2srLQlFg5CUf8kRWvV0uhlqsORM
Ttw59AW1Il2HNT8Hd6PfNpSZWYjfybgefgqZOgmDIDnFy6cMdNxo4re5T2uar1h9
l6p0T2xy/tKXRUa1VCKYe1UpYJxsEV1nZsgiv9G79GsF+enN/Oe+DfhvZkVDXNFT
TUUSIgdbkchJxgqws7K0iJWCzeD5wNfA/RtmHDNhEQ5ZUWkL8Vm1elWcRa9qOelh
VBKTTIM2kN+6R1KTvWL7Ck7JzouKDbcVn22/RNecYQYFtJbmG4fV8NU4e68PepKQ
xTlDHZnW0ITqYRGA3ujQjHG8PnmHpf5NSTL8yGLQqBYrHG0ILaONRiDzfxO+XBt3
gfeaoRNZAzffkVb38wwGv5+A/vPWhwtT2kZUn3X59p99ZaHnsH0fn2Djft6pGqog
V++nGNAfGWnNKkCQCMVktFI2xYCO8N9mt/znu4uis6cC6gWh1ep119UDxFaSPdXZ
VB/09xvoQUWaStt90j4RcslMloCx/hI34l4GnzIb5D4qus6W9sp5mXSrdKW2GtxD
IaX+pF57f/I3nZUqoCxaaXrlQ3FvpqHzQqZANcFB9SQwR6Pw0s4WMrAGI1tKiqIi
jf47DHXU041PIZtewQrSvQU3atHgNgKPIKeRbEJxGKK2dblTjie42yTTwIdqOfi2
TW5VqykUE5JDz/XZtYM2idzO46ekMFM/AbtOuopqs+fLbNJDLVd/1p6q1fWa+Y+I
WnSeSiJiNKJ8Yqb/+36YYJovW7Swmx+XtnLf+TsXqXlBnL8X8n3ssZH+JjK+6fFc
ZYWd7HVSSLqwW+X/7TeqngbCL6ns6R++l5MKT5C8qqdgU/SiHS4I+4QtCVydTxD2
Yp4o5pkDFImuy9kKezy3aAKW7bWH5kw4xLftXxZv1mHhbJHdmAnjwJYKjYXYRb1z
vJ+X66vg+jNDuvmpRUnkKNplichRaz5c3k/KZa7O4Bnj1ZkTUSEx2fG1Jqxpmksw
bqPAWBg7CpNk61hxdJz0FeQ/0+e3yt+ZrTGnB9yC12eLTtEcuVfAis8jugUfqqPC
JcTnO7XyTze01kbNjHTp5AlkysUvKQlfL1kZPpMVx2FzKoXffVAkmiq1A/NQF9hY
xTxGX0yoSmFcsF7V3Dgdcre5XUDUevKLfiZ57yyXQkHgmoCudcAIqx1ftC7KTYne
ieBr0nV5cm/4mUvhp6LOMk9X1a7LFaZQqChrY6WB/4iNiNaWd/TnDuA57bpM7B3g
TYMTTxw995tTi7006cDvfKErufjfOes6vFJ5hy3BAs3YNC+wMrKpzEt7fbAGutE+
c3i0sgbRtN4SSDe3/Tl2VSi3R6agx23krAnFixmiCHcSBj5ub5JUyGUB3AIfFZqY
0bWTktz8G0xKO5cUl0tM/0lmmMT7c45bC7V3vpo+J7ITXjTFDAblZKO/eBOqjbZP
wyDcBcdAndQ0jBCHrTaWspbZSGPBml6DgX8Gpxvms5pvv4vbI+/SR1tyNue/lyP7
pIfUyrCKd5xeB4XkqmJmcM41m7NHtw9WkWpJLxzrPisF+UpJZ+q2N8zMRkR7kKcO
abrIOioIPKpt0+AOXlDbAurvDF12v36KJH20SKBYqI7gfRvxq4wEX1qtIdkP2aCb
NLprqpqxHt3b2LkswyMZI0W1ZC9vH0HovQVQc4ogOflar4k4sfy8Va+AaaCEFeh6
iwfkagMRgwnjHjeAqSCB0uE8BebToneqwuqqHXD7g/szzwftN1OltuF7+ezmRYJN
ei15Q14IVphQq1bba5iZhozupZmo/wv/GzSLkYBP19Mq0iLYUN5XBTYdBg8wXxfO
FvFuafHVHpmNvy4am0sboHYJ94RZxJvIxDTeMAlqziWT5fv15bxJiu7e4U6fKSB6
0k0ang5rfNgYYhywoZ8YbqW90WmpEl+MoGYjRgYmndUouZRSxrKRTJcxSCu1wDYQ
7gSG6C+wM9AusG/AL3G1Clk6nPoF/Ap5hTYwaSLIoqNfRRyZ5qG+oOMGehdmIk0u
oMGQI/koKwZpgpi2wD2A4WXoRoUNPj4wPTWHlbvHbSwYqviJa+u/0Abv6RTC6rm9
2UHHNNjTOLZvB9M93YXwwmfhQQDHVcqedSroXMWT7bP/oDUzLjRLObrhl6NnFvTr
lm8FPZTaizJtm0EOylN67dAcSTu/udAqEy5kQzRmjxnSMgK/3PFIrSCb9MUOF+up
aKMl2wpzW1Ab3Z8TdXPyhK4TU/04vAlRva3LU7avbZCC9cYWHwD+yZp4QN2I04hx
SVX3pBE/jV3xvFm5cV8rXjiLlYgO8ErOlUhKExMm4mpKm9sQOujECAEunn9iDOl6
5PGckJucjruFLy0eJ3vWsO/gX24+k0l4Wa8LDkSAQcdode7GbCcr7d27e8mYhAzd
vTfkxm64tv0BfVlE1ZRCiLaV71GVQzsKH2XuShM1YIrxzRBDXroKdWJhZQCAP7Bz
4B6aO/T/i+6yV0BIpO2I4v/NH4kxWpLudfhBwL/dkQcwUD50DGAoPizqKHrpLIKM
HVS/uQ+eeUx3fi1WI4pWsiErr9SEzxewhIhQttHNx07mgejx6CPdybE9lRph8vhX
xMDYCi7E2ZotNdTxqtVT0f3JcrW+sQiipaA+hq0kxrZltVx77qic1YFgEuKEjd2f
vFA2S3NAxtaEDZQghM2814uCi+1Ud948X6DVY1FljNnw3+aY7/AWmnzYIaKs3m0a
x507Yk++FfGJTWrNIJ25wYNSyKUyUo/3ahBhLC5oYOqyHJ7CQp4Ykv5iq7r/vkEY
DV2V6TbRcm0TJo7GxlQyE4+rsYVJyGA1JOhO9gponuxz87XKp+and6Q1JxZ3ZLib
i1Lwzu9GsSJKuj6Iu45oVfjqjre2LJ66M5sL2AQ6CFKCb6gkO8sDsF8qWj4E13XY
iG8pAHuOjI5+MTdvqf0ONb8YnYi2tjSolyeYopaqZ4TCQs1a+W45+eAKVnrlmUbj
lkHyiJUEC+YMm3kqyRIknwWM513i+MhHE/vt1Y9LZupFKGk9Vr+LkpJFDPZNIIao
cf143Wa2BYGOkRpbhW2hvZccsgbEKDV531JcR5oQjOpoQNGzKklv5GpJxKenIIrv
qz/a0KwM/klVw51KI/E+dJYsJFHXskGaG2iIw6RcfAnu4wB+nK1KHxpUUCIMuZUF
KKXgfIUruBV/o5NJNUvZNRz7MGI4dadv5S34nAC+TIIK9FjPoksBRi7Xw5fUIj4Z
ukrZe+M4ns+r90bamBJ8BMbESR/awy5SPhOgokbx5NcfpHPSQWpHMiTJ6cg58BjH
4aV4PmKi34YXlZ0ThIFygc0/+0psQQa2fktGnSz9Q6u/Y1rlCxJbeS5xNrINRWM0
L9IngM+88FRkfGKF25ZN0l/PgktNFLK19jmPlzXofZW4hq0h8yHAlPrQl5ZKABMX
xNV/QOq6oZ8qfzl73i7pxddXWH2dyj7k2JkEqXhwONgqpglsmG8jv74Ouhsiai0Y
815OkG0T88B7eyNbkhwn9Q8klynYiu/RfZ3gJ5RDuomuneEbuN9QE8ZOFCzErgg+
Oa+KTCy9wlR8mQFTq2H0BCftUWnR0ofDgYbgAIpeBIxnb+8+ULeOTPAqByao9h3c
zy7KtavpeZweCwIJsxov5baNhHjt6cQP3jFrpaNkGj0FjfczDtsGadrdao7h9ooK
VFBLQ0Q1OBa3RIsLCXYIVBgV0GlIOT58kaFc0CHCbb5lvtr4cpaFub0IESFUQgkN
D8vbSwJnvku/+IIj7Vo8Ed9eUeoz8KLC2teDuSKpSm/piJEKu6/7ZyV0ApX8J/PA
8cKDBSPqFlAl1SMqfK+un6pGlc5WREeNs8GKGlYYzJ3Kl9cNDJn8j/wYYMqKLYIi
PCGi2hdy7UOkjCSB7G/pemQ78Hc20utVgmvHuVquEdPe6K+5dXZ+2ACJY07EC5sh
cijyZlDdBvaIgrnXdE/XaKxTLt5o8V3QCPlx/JnAku4JZTnzQorjG685qlTH4opT
N5ioadoG4yZwOU9Iz+7uaGw7uI22CzlKA5TdOoSWuWYLxDyCbXU867GzTkRKFQxV
mPfg8YsE8jn+PjKDhyYMFAMmivOhg4L+Uz90wa6cjOXG4LZ5IVePqypEGPDVB1XC
X5f3EYVZ6Y1Ju5gbkB6ek2RwSfEoP3xNcGT4KotzKr5SpZuoKgSYEWtEZ4fJ55+b
c72gZMNhGUlamaMCxwx3hxC5DYb61NHX1Sf9aQm0rNAKIkwXs5LHiOifptFGBoyO
+cqcmgTdjmUxx0PQMdt5uXaW+CXKXrYOz5BUGKTaIHmT8oxHqp2dcKosza0h7kdR
PhccimTTJZcPo23IdQnvqw9e/nhOu51eJstk8xiPv4FmSZaN713Cx208o1jiLlva
Q/39nhXWWouS2kVgVcNz3h9IbeXXoyzj1sYrGMAewijL/rz6ylt75JgOx/1q12Fr
8dqa6ptRP8Ki+ZiSDvr+IXUw0LvOZM0QIihXV8HIF3c=
`pragma protect end_protected
