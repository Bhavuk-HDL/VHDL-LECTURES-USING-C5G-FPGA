// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
T7SnnWP5pdMLkI0ozJxB3PVixWwP44hKL/iGMa7R7QnD7H+HTQQ3U11C1Q9ILD6p8lqIA5AQ2945
4+iLVpsMmB3DfmjOwYABbZUsF8FJGOQAB7ZoZ5EWuO/MRXx8xaM6Uyz5oDAHlucUOO+KUYRWAg4s
UjL1qusipJoMsiEJDKsjAV1DzHLcenjmxQX0vikFPB66dNFBChZ+1oEChtnc1hEetpQATktlo9GG
w0hJhO/0kV0pNi3QwvNnB9aHubNYwqo/MJP5e3omnDqDlgQH7vLy43y7x/yKjtlWYAzNT98EtBZN
PjXB9vSV8pLF8S9jjHYK8OAVeqtc5Ut4FtUxdw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 30032)
mre/g3QeFMqPLIkPFU5RNRZHNA+4KptYeXq1LZxrDvHMSeES4bGd9rtpCJa87M4YBIJ1tsDswdme
xud+vLpPP7HvaY9BwMu398vq90a52kphXt8rGnp3Um9vnEgXmG2ohgBzod7RikC8L8jNMcsNDtA8
d/XmnS/bW8FO7zjxKMB5SOXYwsLnCpgNvuH2WCv951Rp0pEGikixMqXCYEQKqOPpfPrKWEBU+G6S
o/KESPsRkNcb6+tWEnb+gwG+imRGbbaielsTwmhPWevy+ePrrDbTTTl7H0JnjB1DLHPLSUgyWwTJ
r1yGW5RBLXzUvfP4xyB16L7kXk0VCO2qB1XTpgOL+63EfXqPy9Cl4rkDBWGBl/w9OW0tvZPa80XC
zVLiMZp+blV5KRTOwNh4g1MC8g0L4B+ptWenLEpmanaGtH3Q39SfVhzKdfy9eQ/h1xukHYuDAtpm
xgadHT03jQogxI1VgeWWkHb8sd/SNthhvsmHJVOr1p4mK8uzXFgM95z7V/nq8/NuLQWhD41Qcrti
PAZ+Gg+VUg7AQZvQ+ZKZ6PacvixCqX8KVv/bbl94zfF1P3YUMuTLd34MxLq/qFZ+G5N5v/5HmmT2
FMMET1zoIvod2kuM9JXMYRnms9sj4uqzEVgqldDPYVoeVDlK6K3sIVRuvUAycmNTybzIFKQ1CuSo
HmrBuONDymesJ6YXQfPB2/FHRFbFGglKnMQqRvB06++cCa36gce1eBS5m0gwROSb3cRd/f6HMVds
7HZeFro8PoRpYXU6/YLut0iFAfBCtmjYtWLepGL2JLE8jX6VDKqJyKk9zP+QgBGSrzRIVO+BOjFN
LFo06WXaykHJQh0KrvkJ8DyNwEcyQKGddYd774FyQFC+3ZbPlYPbZ6RpQsHVjATYQowKa/gM264W
mqEsW1WjWpjAIZQVZ4RF5WOR9RhRMwNWsSQOxyD8zRAEgY+YdXkP3Q/duC3XvMw07emZ0xR5G2lJ
Po2ZZ42sb467VeU7W/eVi2B5Y2SPEt+d6uT0ItS47zbSykcRZe1e2UNxK+kLMdVDICcpTfiSP3nj
KJeTju+rbZrZeApOv2ROnvg3PRDiw00VE6kW33++Cd84ANMDowW7ieg5bgT/dn/yIR85qEXb6hnn
mszWgTob73EzzncZcF5eOMkXwfB86x807quAByi25oMKeRWyEFTfAXKSeVaUha3vlo0T/cd4Lhaa
OVfd7S4HMdasLk4BXnU6U3Rhok3T7y1BpkbaI3h3DQ5+25Wd40/7oa6zV9MVPopQvIqGOScsFj12
Ao1sSKeJgLC8evAh7UrZnbdjb4wXltsSOj+JZFIP/62xJ4TeXBF9QB4UoqV+a35VL0dVkmmyIGQN
2WW0qpbqjoP2TN/rWLwKUYXCKBYO9ukfGv9lHFm5SEfJHEwgbP/Y9bDL3/W85jAgtl9zHRrvUTQW
n62hGmjV00tKE69j3y3TRM2rPW7gJ+Ytq/V4my0cI80SI8zG9Slm8llUohfLli7LULy5nWMXCGUZ
fLx3sBBSfBUzZQ2AxTw1nnPQSOsxFs+kJUmUUAPvUICG+L4CTlmboa11XQGYbOvtClUHZ4i9fNv8
YA9wk72lkc9AuI9ph41LmluOLdl3+pvbTb26ulMk92vucEsMhi3hmApcD1OpYe8oMG/pBGGCSp2z
6ypWJw9uS/YtGlzczCLaa/sNYIN2JbLDNgKDVDedD2tG6ZFiJUht5QPze8j8xXna3WEDAjDIfeL1
Eaw4e04wsmhwhE2xpqbKubjOaLhqH966Yn34IghSjXmDAqhCRKLviUchSEaZ2XBQSKM2cDKpkevl
1hFJSVeENDCaRSUSAbG6WF5XaNETosBPRf1E7k+YJjzwB+wvqSDsKMJN/Bqc07XUQFZB41XM687D
mw8+ZsMUe+t1sgJHDFKs/M1RT6Oncb+ICHFUthPoYw07ALM8FgPUk0vSqHxjJYAdcjb0paT8qGyA
hxGnh/7sFN9oOqELv1UZRtyyxv3BoMicCKaR2XdCwSgMKpwd9Mk3ghCZ9kwf7jPoGRfoRUQpdyPL
OAhpjLbjmT1k5JGlwmxPYq2zSvTpNYtog3pv+Agv7irCXR60PCDQ74pdQdA6DZZ0kC73eVN2mXN2
0AWIQ8XjX5fYE0evNTI34TfzpwKFzpKvM89nmI79aGA3DAS0A9gB2pAC1Iglgttqwx+78F2hNLD4
qQKheAB7Qzwg+gggsLMD3srNPZfmjgTJLomtPer4Lv4RTPukGBDeSwoom//AzFMIgHqTrQeZpAwB
Skw+sG3L3mM5Yfkw9bMMstEd7LE9CPVWOsfCuuOg5SdYPH7qipCBQbJXX63P+quj/Fa+Nm5riWol
XLzpDE01D90lSczoSexfcJKFvAmYdVpX+kvubc2v2JrH0VAIDSA5GMXaHx8JDVO/COt4/ET1nO8+
hlZGuxuZ3v0HEXcyFXmQYhiKEbLDFWCGFPvGN6yql7npCTYxv2QhpyQYhQqM43aMgWOBUhvWKpAN
ykb3yIS5RFgmfNjbzVDtOuZneYUohKsG9hFTq684v2y5P4FLt2yfdRDsq+LmZYbp5Z1CHsHvjlgL
+4okT5/Wuz+elYKf/9EsPHHL6VczBvvwVqX4cqXIQdlhVt1OZ4rqUnwnw6KFt0NSULJgR4cY+r4a
wJCuWmW3yOQIIseahLfh+AG+fiYculrPnygPSIAetXSZEIhLVzdsLQvVM2yElsu/zk81ldbBjG2X
hiP7oGlEdPW+nVMlD5F1EWtE3wqvscFRwSJoCoTwmNWrfgr43XcFjPTLEnl5cQLPcZu/g6UrlrcJ
J5ozcRUH//q5CxTXc+JOXsiCHYD7gH2azudnCkXGpF3ks87Vn76OdinD4/oVp00LJ0RdgDkl2nzc
TDQgdNCx3xAAaC3upiVSfgt4XZFY66XOMiG6RzqHn7N4nNkkybaVgeo4WdwKX96zjH3/Q2bBGATU
gXz+MTO6fT8+PG/Q9S2hj1n9RlYskKAdPK4yCrRlOeUCJe8dHn+AHMSOIQGmMc34ijh3cW3yF9Uq
aG2+OszYQUjg7aPysCczv+l16Cp5EycdwTObW9HaAcQzej4yGXBvZo2MVvheQL1KHOEDFMg0KnSs
rQT4qitKI8gOCUtciGLBntctLlm5roB8EVeB4r9NOHS4+KypvKX/2dxTUmYLv32TJZru+MEKe3Yv
240O0/MrHfflMpmgNDQrTYuYsEjho5X9aF1WjsvR9rc2zKn/01eh1+RPk9/PjiSRchioy0KXS21N
6Wn+zQNAtz5VjApX7Wp0nld7NwBVznt8fhsv5mLdxNcFj7cCURCvx1Q0EP/LktzDDmYSZcNi1sCy
THVtjgtQ+U7L7YE1PgUV7LIHYwoebzjBtxWL2oWXzaIN3biWxNbvhdG5VmcLzyIe9Zmrc+nfCUmq
dLZqzRADiSJS3w+P7AsW06bqgBIJInlMuQ/WClYu7UJ9ZTog04nhfaJMlneHxe3i18o7waTPN+oY
WsVXHZ2lNq5PWOUhG7qRLUIv0D4E91P8g5tuYAgQlql4esyA0xxbO05FyS8UqMDlHAxXE0r/C4O+
60cdiNF3/TUsuIxqPm3tNs3ZuygHGeLTNsPk3pHzZ7fUM2GkIhVuRsuHDOf5aHcIIO20ByxN5jxq
GgWefWENuRN6KOt7HsUd573wEDrq3lMVggzxBkKwoDk2+5MM1ApYflW2VZpj+Olpm3sAdcRrrxGL
ZvZcF6XHCVPkgD4sWq/3eB/O3D8Ni5CglgGlNNnxbXSheoOqVwau0GrOOY/HOB3fyc9FiYZSophJ
BjAv8MWxs0Ift3zs+cxqHrl47oOzCph4t30R0ZXM7PUfSrc/wh5Xm7LDouigRT42qXoJGzsPU1db
0cgQVthNohjcelD8QURijmm5Zdz/2Ae9d84haqZejZFf65M8xgLAr9vRCYk8Qfc4MlGclbXSGEOF
s2xVi+P8bnc9VZ7nJ0IL1hWsSOsjD9qpTNcxtM6t1+8Qm5JfI7DjpcBmxcbKR2IaXDv2gUU1ugAi
ZTy/4+nJ29Oiw8HRhVgNrqHth5vd4S4qTJV+AH/Pc4BVQgJtokUz+7y+qKssiBjFFCB30a7kZzBk
0Yp8f9rv668ZpoWUtEa/jYtUpnvYJJt33iE2TVoTuQnC6ky0WAO0Tz74WOYv9aItBEZl57QXkQN9
T0QKi5x3MkH9WlK5R2FyrYzcB1FpD02Fh/acOFCXaRxLg0M2B8rlL66+sZvkpzeH2Z2ybkWnNHz6
Oytp0BxFodXbP9aBvJ0cQmAY3iHVWCCIMG2ZpoaI8waacUeJoJkC90+Pf7eGKiNhIPmitbN/Jiag
t40zHtus2vTmiBSRPNa70jETpM7rdbX+OtTaIdE3exwLfX4dg7AlXLWU9CBe7yxtLHIWe2Xpe/uG
6PglAAIAgH/5FnNbwnuolWn86nUaB6SFwW22SAS7/xAkOAgDVeUWionrC/LDFTDCmdqip8UpglmX
nCSY+WSj7NI8IZyucZlkDCI9nYPloJkB6K0hdVrMQi3G+kipUqefYSRdGjtpOzSzxlyudiFYY3yq
aXgeGSrwdYMDvYtit7vA5WTTYJBY3VFffmaoILZrHT4RZfX7fMLhoi3CUoKrWaXq1y0T1cKCMpYF
c6KZCZ78kpgJCWZmCg7+x7VGhzAITLWXDTcnLrHxloFqUUvJglecjdSiEIOIKByWpMa9XU9IjqSe
GxlYQ0sV66Ehx0IF/0I2Vxu4+mY1lnyA8fB976CT2Ftge1ip6JPYP9mKvl+W7XdddoSlX15Xy0RH
BHRbGT2kuj9BLBd+o922wpeTrCsdVd84DPRfZwy/fE7EI2ucCMjfxRymg9y6WuhH3keIUXyJFhsR
atRfxSHgMY1/hro4yfMYsNa+LUHWZ3rh+YhgBa0Ahxt+xfgmI9nYCdQjSXviIAL9mBNaiGRU6PdW
m0o+k04KA6hQL2CwA1OUvAVBMMhIZUwVkSG0sArn032nKe2QtwKHefN5TqqJ3MVp9Xf8cnO8LMMH
QRHPygiP/pL1CdDqUGu4U2H/K8v9mKZlRIcgM/YVqcIYJWJOVhS8Lsx/PdOLFotV9rfCaRRmje8Z
DbW6jYPFfeftLCZi9GPYoPugTJAWJGq0vy+/xrGdLt4oDnKZ8Z+8kBJrhOuIahDPqbXfSC8ay6Pg
Xya3aMr2lPzj99DFKS0vwrd+VAk3mDM+zffcdMGmukiNiIuWD5vMOEi3wozMV0/+oy7YeBqrLmKZ
fx3Bb5NnRac7j1Foa81QiX9+NbpbsTZv4fkvdnVuEO3Ck4NK+3tnmybHOfKKL6cPUf59RVSTy7Q/
1KXkd8gBMubtXfdmQ8YW5S5tagrexbCjV8qcRpoy4stOi7RQ+42pGFmw5IFt0Xgymj+6uWakD9IU
TNdHzqML4iDjRK+A/3oY4SGy87kZTNb8gYj2GRP7aw1uXJUJrvOWnrVhvvWAc0JCCVv9x1llB5NM
jfMoLn/wcyr2dFyDLAzzcRdJT4+Eypl4qWCtyLibZggfbeobb66wGOflAvyXzmN38R+iSX4GrDmK
Or5aMJWZZwYkrAfP5Gmp6wdUO9yFWKn8xgkRpIvug4BW3W9AZVWSuZLLprfQLozdDOUF6w2xMV8h
nw9RK6Rb5aAXGjtCtmg0RZAr2Ul7stSAiPqGhzCbTTTD7RweOTWBQx+JGxwAvSR+ytin2PT7gNO8
hNHEehU24KUikFcAAOuUuJh0pQUyvzQOU4LkTBz7OOizHkAMZiS5uuEKk/QO2TU9CFcQ8OPe0Oje
9rd+MqrwTYLdy+yza46AWVQvi+WXukGFwUQU6f74WBrqC9Quo+nDz16vIHfUXh0AGDA+1p15dzZN
4cLeD3y5SOKdohmDMKQLXmo20A7MiPR9AEyNdNsipaMYv6KrQoPC0b/9vuxucHqz/jd56a5hFf+j
5Xgt3QDUAYMubg7/WKWyUofuQsGMKyJxGHxXFGhxyugVqF4hAWhztWZZF6iuJhsi2Iws7Ge+ea83
F5gvXLTa2Ft3zJY7k58OFv0q5OW8Ls0g8lIzU9u85QxROpBGdJJupjMxNrb8sDg2fMVCiQudcxdM
C0eDeXRSfUU/HckSYQ4vqwB1jl3XqorIidC72Hf/08PvQQ2dbyfFwGHTJ55yn++zUx3AgZ48dqZW
eXkaGpQfBKHWuY4gB25ycYSMfREF4Bf9bePUs1kCnUhjfmHYE7DvjXKiv2N63iX1rNu8xGo8tNDw
8aIyjk9KrLN0U4eAFzZ/Rq8QIe9Z1k2iFnE7orFXppev9gkqbTnJDdGYD3ds6TpAuiYmGlShLpmw
T65lVUTz72AnR1/rlaCbgiKjJgFI5fXsty1dpO12KDmKvBBmolbwKFDGnXoPSv8+QDXnlDCS68z2
odRzbRIeoql5Bu05IovhuIGjBCZRwXTpRXC6S4hs18xYlRCb4/f2vgS4DGMUgJm3A5a3bedhMXy/
6Zp9dlCTw4HesHPvCWH4LpegJC+5Y59soIvClTM+vl05hH1fvYFt94CBeIxrZyyJ9AwJinOpznKP
KBMqWl7juoSPhKr/VY1CUyLfW4w41uAicSOHQGtgZ4MhvdWIPy7iPEEwXrowuIM9hpQipyMDjhIb
Tbp3nTQOOfDsQiUxcO7JVVnyNNY4Zc63fUlAZx3DJcMAbHudwKLJqQREpXt0DuP1JGqLXayy0+cT
v57M+tbFnTR8A5DLb/HgqAmQeQ8GeZaPgKK7S9Un+PyMY5JC35Dq5GoXbngVnLsHtPCDnduE33xs
Rk1QKQ1DIP0Rszz2WYHIxF210hk57wUg1ui4USpWLQJkvVat83dAKgPNVNwe5wdJ71K39hGdXWn0
3sfPwcFM1alos6tTuAEpB9fnWNpWUDWNFn4JGbeAzuL5fwE/OJVmtJg+XBWPbbaIyASpaTsS/2QD
0ZW8wTYilZWv12O2lt/Gi4ZK37KFJl34Vsub0htKYyHB+3H0czjs7yxB+82sIUxaWleuDW0+2c7Z
DIkmptlseuuRvJ3L/iMi7xu3gRJ8S46U8dIigMa2P9qaLJR+zQ+H/6nCisv5C/6/lPPdQ3AYFjxD
nI+92shS84eJbaXKkMT5yazdWNMiQ2QbARxR7CnozP5JZ+ILFD0ovH1eQRMYDbfvLwTNpk3Mqt8o
0bQcwFNsfEU++cxhpQW9KmNwY9Cbv9Dwz1UJnZY/dNKostJmT0tQ8n64irxcwVjNOMSuLHr1F05S
pqyfUco9KOS9uIehYq25dck11WF77ZLpCT/9VFw9K2ofg/nyHguvgadPABzjPT6d0JcztjaI9sjh
7/Q+por5z9zffkL1R37zGD2rBuMQOqldcOjc9++CAOEXMGbWXgjoJTQtLg9Uis+WusUFJCWTxjPz
pUqXfwcnX/X9Fku1ro9APjM/Mnsut5vNkjlfK6p9Wf8TxB7Z7WfCFXo81ogBeyzRo5KiLPngSJIT
skfbA9/6dwL7FK7REM45TQxQf8CXzpJ67yfUGvYvD6tvXXqNoy8xifFowAfZ86J3yNRHcf60IZFq
sg9VNDy888UA09JmYI2HDKh54GzvTZKu+xV02Slzum90QIBdZSzJQoTig2H7E7VahmoWiWUfNO+J
bvawH+XbrE7lwjlmsQ2go/LaC1y8eg8cGiMPmRnRrA+rn3cU9iihMUPH8i5MteFGrgaRE7sGSYof
rz2OmxrzeSHOlXiOtv9frmPlXDF9podUO9J/Mz1596xTQieY4gvHF6LmK7YaSNo3KD3xFafVUa93
VE0aEKL2BGfbZBYZ2DhS/EVQ6nelgQ4k2rkZvEVz3XcFMIDFn3GaajUp9f3oOFv9NCJMU2QqyD19
dhZZoQWBHCWQeMEG6XtascGvQPCH8erBBgIuPlvibRd9X1YkwIuKiVplTusUStvkqGZF2DKi4SvY
OnUu8hSeeaHjB6hPSAjYT5kuyJGca41f6DRoDjyXbHWMxWspP7x0wsYY94DhMBtjty+a8BAdUxlW
nPpSpqeppNYo+8GRLbsTm3phPZ05MHL5A35YqRIrljCtFU8SmjoVIMEhkUekj6OpUEtlhEPLsZrs
qAgARkotFwu/3hA4l/EFPBXY9EyJN+vAfKxOk/DALERwSFod7Mo7hfoFhUMuI4ToeKZvX3ntjwHK
MFcSWF7/dA0XWqnXqtzwaD7BKbZW7JpX7K6UhpZpLX3E5tsofqbrfDOs11Cpt1jUBsQWAm+1s9z5
v/vCdkGh5MOzcVhg1sjb40XROhYRtv4LfYZUtvTYKBUoyw3+2Ib8kTdh9UwRWMEPHs4yaOJ6G/CU
q4K8dBvqSOLns0sRv37d+5cHcRipup0UJifhip28TCXKVBELUzKeoanAqHO9Bsrw3cfmeczTdgr5
WrnvDrxNHSW96brScJfvWc+pWgdLnou8TXEszxGOaLZoLgW/qwNtWKq9I9sycZG2b/tRtThK4Eh8
K30I25/lLd46swkxcMXpC5CDxk3apyioTBK4I3cAcchdCDizaNbqbfWjoDFV7VrbVyTLjD5ru0hS
6YlLrtKY3ckkbMnO+wYFL8jY8WkNbuOYUFUZB7txRrAo4Z76F1fjih4ul0fIVscKJLn4ZLa3YtaQ
PfDoow0lqrJJXH2/gcz2xNcfGBltNT9mcZvAwPmA+t6LBmpxzVsS33YDkXfOFmjDiWDIHwo4eFMD
z4vLfP+fKVAWOlzbqh8uW1QGMPUppW/Yvj+56TusdXozBdWjH8I3yAcdmCEyvmFW6iU9Yze1eQEP
n5Iw/EQU2cxHgsc7XCPmSGqByz1slpnFvT1ZFiMuOJClgkcnA+IdOKW1kqCXSjBgvtRetulg461j
2FHfd0BpQekqIwvqR6XX4wXuKLcYvNkSxL9HPk8Vq/vCDGTLIFFGrUOrDRBPKFRaNKdK3ujuI73i
wcD+oEclNl8w3Hs7NODgm8hkRS7wNLsKHo9yyoCMg8cpDOKhDu+RhjywnuSnFxn2W4TE4OwqU6M+
sqW4nPIS0w2GtdPZNEGtWhlL1YJ3z0MohB4naKcHb8GPfJE4T1kCSScwJgXBHe9uezn5wOyUMHTp
IPwakdO4Bhbnk1vPDqnn9ucq2hYE6pDeb0raDH8zB+9Jq03VYDshD6ftMEGEqXQxaTKJs9KT2KZJ
j8NhDqIYmOdvH3LCUhuI2NuZhV0bGvIBrW2j/DPnLJIac2yKg7LdwY5MznnszT+6myrSOhp4l7vj
i/cD/pQQMQbZhNY2nFxj0E2kuf9PXW3ZK4APoUPzaSdpr6c3sPKeUzWwq84Uo/4V9ZsVO7fZ5qJE
dauF+9+mCIEHhwdnuPubTL2PJJJR86oweiZqQFUD6F/sXvO+iYenu9bsHQzphUG2dwK5RlKr6G26
7QnFDAgN3+zdoFQv1G9Uc7ztFgThnJzUKk1scMjDZBcPF6wu7CJ96ES8T9cNSYoRP9JIpdZPL0a0
2eoSibNpy6d64/9+4lu8DT8y/yA80q0Xs023sEbPKaUQWkRdd57Ns21dRr6VXyvXlykbZNJ3Uels
j0IXEp+9wULmp6rlAh2YzJduHcUB0vNCVbb0PyQemD2SZZEhKD/N4wdhPUf7WBupKeSJg+NoQxE0
7jYvg80LayM9R4LGYMUFSAiDNStlUQGvh3bXms91foI2m2LS2zjLQy6YG90fvpNyR862inobojJV
unSJqUaW0ALR5i1NX+J82mIKJvW67QsR9wpeP+whoD71UFTyxT2LZKV/CeEVq+LMzu6XtejKSAs2
8GNEe+ZgDcA5wsFwYb4Cs7UQIdBBAFxV9EJQdOvYWSulCuzwuuWm9Z8WhM1sRGTke148V+DU4W7o
T54BwiajcEif8lxJx25Fnd3MLveZuyJfiENE03kG3Y++UWyAyyYBpvLkvut7JHElkBQehuoQ+3LM
CAX8dcv+oE7dftM8DN+ajd4+KNwY0y2WPXZAKwGhksD3vUrc7jeasUyizjtihUKrM6Dujjacxh9t
L09Uo/q0qs527PMQEIwkNebJ4WY8+khQlc7Hk+xr56JOJumU0+sIGclFfL9bKfnppLUytAIvNSeJ
AcTkPY6Wm4mimaTSq2j5YJfa5rXPlc72pulFGvByxE9wRW2doYIuTABQVW8n0Vbq1xW58ZoX6yjw
Gg4DXNxtlDhtPIYsSFnSKYf4BhKn/UpaPQ3r15saBV7z6LyBLolrhjoVvfoTshOOLO+Mp+OeGFJp
ITry4VJ7q8pCF07eWHTA2MND/gOMq1QRW9WhcKE8lkevTOacs1r/uajVPMfx0xHmG9OBCiQtHLgi
YhMTU39cGQVuYtcnA/FGpZIAfeTn8vY5tOsH3bGwTvJHa+zKx9SasPVTC1Y80dKuFBlDFTzO7v/X
4Kx2O2oVGdFbdJDxTvJO5Ea2T9Clj6Vg2OtQ4Olssw2bTXwEKGlPU2As1kKVh8GF0cT1HidwqBlk
iRuwmfgNsgkCQECptb6tQh452LRh3YKq7sXVWRcXkIF5GcK7BaFFqx4TxEQoy7vBGNv+5le4HoVq
QHS6TRtbgRQ3NrMV7ShUco3HOhRqEuwWPcDyJW7zUAUyR1ojRuN1t3UFeeD+eIq3nAriiVC/3gxq
OAwEUqLC/qlcdw5htQBYGtT+eBBfJDQka6toOrSYwCkiVO32iu6d+XnVELjrnWPIuQkFzYSgj/iS
XPYl4zF86WqQ35NKKOzMgzqK1rJcjpKmazqNX6KGaFZkqSSioc3aO7kYXjokMlrnSt9v6knoGGVz
4/jPUF0swJpNnOr7p7FYe7vS25ejKPKCD8BoY/wNm4WmSNQWvkfW7HGFb1LFzAMNY/S6xx2hC2Ed
YtzcJQKcEUEh2cXVj4eiDNn0tO1Tfc7TpBFxXhitMxFmhYwCemlOldCGRPNxVx6EZoDW1FzlnR8d
U5QepyR4I0OX9iDmgUjzu4AIyoBZCI8lVrFkL339fhZ0t/KEFXYC+R1IcnszfEP97rHf3mk97XUW
0Kdp0dJ/oA3frsSzHPJ+j/J6B7BbpvGiI1mk6AQA5M0NYpnwk5syZnn48AJU5KWeqieUehwzUXq4
mxNjiBogQQWp39BgMytd0yYbCqyj2tQ4Lry00yJEo/lLmYVl3376BpuriZ/dr6wYeyKgVeNOwKo/
3K/UzFmfdiBt+eDRNdeIrRR7IMt39zy86P2ERbV22DY201otww9NAO+M+7cSilLOr7uYoBdjqcGY
36PmoYygePKYmUhUg+EZ0S5tjV2FKqaUps1NFskSEtMqS4GJquLbYSV1Ig98j0B8JKCdIZ0a0G8r
5NL8hf5YGmwjraahVM/r6ssOHRN2uuMFVDs3GRXbjPFw7R1gLtPu9r9bn2ha+mx1Uh7SX/cvF95O
LOaQuRnCsBRqI8CNJ6qsScdGmDgEo6FLOf/pmyiVz8BkrSN1hc1jh3Epw3EthOHah1QvJtxmG92Q
HqLbxfvFrsC8/aYgL/uXU8Nw4jyBe9lylVvjKf8AURE6YEH/R3rd9bPilb0xVCfe4SL9bxbIlIdG
WZoajbu4JkjTMLgtkZST5L0qEuE+pNl//JegCm55zmhLYqVtxtwxDezC9qyKOrMwF6z52DOngsR6
ZBofwhiPoEDPz2w1z9Ka7c3D0nGECTrDA0NwlVbEF4LtX86NuWfEJ/OUz0BFNR4Rg2Wwnz1TMY2L
xuRzyT6BlH3pAasjgaQbQlGEJbFBfOktsEMyUp11doPqpQMSJGlo3cWvootF3fjETj5Qf6ly2YQG
d8UQpcCm+NbtDDwgA8yWnSMiMeGlmtTJy8HkZgd5dy5lSayJClPreAuUmXvRzRTA2VVB2fbZTdiy
C4EPX9Qj+jckjg/k6y1frrFCQwZVGW1ff34ZpZf1TG9LPbM/zWM8Rh5gBhERzhw5eydYwIbUYt4g
n0CsGLrZtsH2YPsj8XEOZ/N39PZwnreEy7lk5dl95njHzhzlZRwwrkNZTENiDmVPULXpInFc7Ku7
1zqiZqrbpNND8gFyd8OQMlevqhbjji6fwGB6GJAENbv7vm7UBYHknFyC0W9xEU6lE/rO2jr7DwJ0
dUek49nIWW3fh4Aw4EtPg7c7kU2se5pHSYtL3kCQeYT099zvtcakWoUOGg/AQuQZtoM7/CSXAdgq
qZK5n54ZdNvheAjOr3tqAOQv9idmTi3sMQ4VQ/ENbl0I1vU7UX8OY7wEOyUOTZvufN+iZz57rX6Z
QZIlsHd1UTW9gGWsDcSZeiUi3PFMd4Lz7XMBCXqMDAkRx+pHF4vhFXlPYOF+jgqhnXuz+Hf1ej2m
CWHfTLNQZMyF5Q4aVpGGtNabsV9momn9sQ0Fa4u6IcwWmOKb3l+S4ekKGaBxnfAmI5QQ967F/1kX
vv2DrwPPfGVxe9Jo0Wb0UpzUyof2ltXCxc6CYXyzWUFGzGvqIEQPRbprLpxwX0lkMWgPBWdUIqTm
cOXM+68onCFfsnCSCyZUS8GE8uYR6ipSXVsQHE/Hg4w961dXpTjH3Pdr/DvhPa//KGQOsIr1PVTA
gNb+5WgthRTFn/fZ5SrG8X+Hn+Cb9MNJPlDN9RagFCQlTazh5sRwvLMby17NuU/8K+IneM67FPvE
q0Wlt0YkZaKjHWSr94SIgs3WcVxiCIzHv8XRDxzq1qvu5XA/rTnvWVDaXrMJnGYCU0eTkKjiitfU
XRKdk/quYsKpUt3LOLxaPilfc9OQu4GGy8lx1GDw976bOwgtYVutip84W1fLPoCtF/wr1stirI/o
RZqtjkK2R0ahjjKuCTxAgRTow4sOiIAi2gXT5NEvVvkk6IF7pYMdtaMBVxKC+emJmUg8B/j2resP
H5yW4gu9jpNZh9oFMuEnhL2fnTfAKrMsvu1OcF5YcdltFCWH7GO/4klnVvu3s7M0VAhypK9+oL4i
CVtKmEG+zzLhXQVpFYR6WC7k8sYZuv4aG26uylMcMVBbYwoqx72IfG5u8W0SgxGNJI1ccQgMozfT
LA2fFwHjzNKM1UV0e4kQaasspbXZNY+ipmQqaM818b2ZnK/ouSFsfT/o/KApVypLJFyilJ4ltNSR
LTXxgfeAF2o2hkSWLpoyqm8+ChbafjnprbessdbARvShDoYbwVBvLhceIyyCSfD4rDKJaeZmED34
c/gk8Yli3pLLk9h8GxXUWCBq8xWEQWAr1ssZJbpUZt0OfG17pTA+pVdnKS1yV7Ulnm9reJvEiLBn
cwpeOIagykVuVEBK1zqqbgozpuKltWEFsojXbhmGEja7XhPrygM9j46DH7guVXaMnYU6xIo+i43K
CMqtsmhP8geZWh66FZRPZWsokpq+8wWaKnOcaRMGWVlRPdvJBE0MsmymwdFjgU3OJJUyYgkBmEwE
6Ox6uXamg9cEJxXv4DiIEBmAajckM1P/5ScS3DnH4KDWQATycdYLi4so/5/n/3k25Hf+lPYXZ29e
PCfGxqPJOQfKCIFaLpI+YOZn4Wh5nMolHP4wfr81Zh9XbZX97ElStsM18zHtqWP3zGGHgiEm8MKm
ithcE6/umvY/jgsg3OC+uD/VB+L/cYBXHsMukjGtLvxK7m8f+aRlHE3PbCt+Wz1tpIolV2EUrOLJ
HnnLAxbUwh0Ydmk+wjwY5UHQZWOH41E0lMsz3ECYMup1KzaMp9UfXSpCZdBJY3+wjYXgJKJCcnF2
j0FBdQT/GFejA7K2A8IbtCqfyhkCOp3y2rWLH/yqPKWPARXnEA/eoGaGVWefmuucNjwNgLF9rfGB
rks6NaoeotPJ3tAi4CBeRBegNmecsgbtl7egLiQOdkkOH5zjeJW+imRT9Kk2mBt5IL4CCyMvemX4
jfPBthdiVQOKuRlCyCK4SQikXhu/dCTHyp3KMTm4h2vdBJafDltpyPEGxStdstcEJwgOF0/oU7cN
sTM/xkIRVuZRVna3Sn6r3KqnU4qf9DHMQlj+m3zST+oXddsDi2bc2sHka8yKyLar4zzl0yTn2wzb
GGiUDWeF6CPTprRj3HKMnBtEm3lCWM9nVaebXNbvLESMfUryzwFqLDfBbKX9V/QKJbeyaaqNc4In
qC8u/KH1F4rncHWk+5qtlQFxSDb1juixGdrZshlxeqf5NKQ0/nr3p7BFEbQ76fmDJ6i0EYwauWcW
cvXUfQG+R9X9g4kgzQG+vsuaZTc7pTeYaQiO6Ht4EZD7+Ysi/QdpffuDnDgK115EoWwnd5To1eC/
TAspPxDWTruQ5gFpTlTr7eD7qLMTsnAUA439dDmw217sqxij6YlkMmwjbOrQMazTUDL3spoJFsdu
3jFyx7Ix2I6yjPoF7gacKfKoAOHWyiJQKUeYMPvXjDZe90Ob7bmX7MDsvPE1UVxzNkLp27GbmNnC
wCt59KSnfCeQAAu1NZU+EV3AlfDtRghGouAE+acll00JjYc/n9X6E+yfncpwa/kTqu6ibur1vK5W
02kANnHfUobUEyAfHJmXpp4Ct49O533IMs1zZ++ghPzX329v0uKaJVjhaviDABX+LkVDsul+2i1b
Fp8vfqWaL5Sl4NpnQHUn9E2j+zJSIeyWnmKcPXugK0Wpo30K1xivHXIK0tl4l78jUDo+LiAf/AJ8
NnaBdlDLxcR1GfaYD1d37unvGSKLA8bEdY6IXkL7V9VzGFcp8PA97SUZR4QYiiPv4mcJHUHTC7DG
ra1xS9hfpEwJxhEBfUurNFyhwzg4K0AjQbSqmHL7mKCQMMD26/chP3j+EeG/to4lVdyjI6EEAqU/
w+17AcL7Q+/FdEVsz6FtTcpvN2NT5upH+f2THvI7BnleiU2CAoFAiLr9AvTHZyZEEF3gRBro9Vk1
/LRX/qWvuUiEpfPfsLNiQnYKV0P8soV6Cil2KGrrccHflv1thhu7MArBJzz5rOk07YIsIQvpmMWe
NwD3Cdou4iAyHVgFN/oSNGELD0r7EtvxyWqH6LTlsrl+DDqzzPv4HaS6Bx2H4KNq8FKMUqYRQ9y7
MltAyZaKhJvgKbbXeu1LIFRD8IjhR1Bf8rj/sYkIRVgmRFtAShRxqaLZxLnKFj3S6/scnY3AJf8Y
nLkF1/npRsY1jQ71UpKd0dJTlkkbM1clrhOiDWTd7cVqrgpNUV/cRs3k2rjyOQPIL5jkisU5/95E
dEAdS4WiDL4pbtwkmg9lUzYGmZccJVd/LSuegTGGcA3a4S/xXbQNZ69L0VDfiQDId0pSN/OWzauL
CkcX4VsQIYa0qShY9k22MnwQJYjN/35ycv7UWJJY7ITaS/6e921tZNOsTj1t3Houd00QBtMBd1ep
PfqWzyytUBu84GGve7qOCAsTpUDNPYSE2tqzKq6h5zHvqIoHyNdXeKSCkSnQOR4ZpP2gHBU0Faju
ExNyi7h7x/ECQYMRWJGfxwcdfTyKZyFNDuRy/Y7WIh2US+aAC342WLG1Vrc/SIaNZ0qFb1ClH9CP
iEVNgyXlDwrmLW5oEJsQMmwWePixGUpmGbmhLq2m3I6tuNCPLkCkF5H4lBqwY7b9dK4M8wJ9LIC2
M+PfUlC01OwtKtQOjrQiNBJv/XpHS9dvgQwFoFUZq2BISdf7Exf8LQPf4kR9wtUNgfMKOmRKn4wc
h9jU8UUArk0PjCU3Mp06NpuhO18jh7I81cZ6RLwUbBvworQAGTGfuga+x5qp69PkcK9relDaBe8w
pGmkDzFjK82J+Z9/YjcCdamHX++RSmib8DpUJyJekchC1PljqCvLy8CfTCRIxSvyfGi2hEhxUIYV
VBC9vXsa1kTrihjjyS68AS9B0yqv8hy897B9Jms4dHyN+/GXXgYyX75+YzHHdxC75nE/InaOfJ69
7a+Z25zV3Qpc58M9RWHc/c+VEnvphy1I2F5MR1Idrej0n1xmWDdG6r9GIQ+eT2TpUpfIeHqu7xx5
6kT6brWi5fDCbHumEC8OFSJ0EtpLxosLy73GM3Yjc+IlIEJJnQ5bQul4C7RVDOq6s+KQte3MQseB
BKTDGs52whvmQ8c0woRViA6yL/3/KZ325hLBT3zBjmbw1AE9l7CM5qBRmMyBJfyMu4NsxdvtElFm
fD7p43n6QgFTr5aAj8wiV7s29TPMyIdhTPC7eRbdmplPpnWy50TySg91tjoipxbuZRPTlggvVfTu
iD5g+x2PhImYXQK7u8T9kMxt/bld90mdmGtK3ZpDuyE0dozU12UpSIcYHFXbDnpX5aUqMxa0I5vp
8AGoeatjKSK/R+29bv0ikJXknctBySzjjrO9aBFaaP1/vOcbUOthIX8xThbdzxZuvcpCEN78MrtC
iF0PYnAceyH5Z5xeFRLI8kFQsElvTrSAVUVp0k2888tYCIs38Vek2q5qmeplSBzSLB6FYl1AK27H
3ozJPcSb86zpocsagTL8Kst4bBlu2LjotbRrj+lCvqXbFezRL/P+GZmBzL6306BdcssvD0ZmfyUv
CSf0E+lUQKFJMo4uSmIDUC66X95aWQnA0j8WnpkwArydVxwaswjyHbQTmWD++H8a1qtttbBZRAID
Ce/nTwIdAaWnK+A/H2BDO743ZQ8CjryZ9XkNcBlbxp+JMmJErOv7gPDU12AQlqEj1+153+TdVtX6
60twbGbhasgvTOeRZnkU7ymhp5/mEBSd91tNaRlHuT+3ap5XVh7aSWbM8OW0DT4ntEXJzxWx/onv
gKyPA/wLt7WlPCt2XMsaQI7tyoYmiqoyT9AjjYWwSMTlhtDbM7JwTnVe8rU+401Q4+3Pxj53eu7e
du8/I6ds2CdLn7e/nOhSavGBWc5xwi7B70HUG2/nwXJtbdfwL9nVeqboWDiu9zp04eido1F9LSjz
JvgsHbrsxP12S1QLjgbII/kFAHkq3S4ILhNKWnVmWDK31IY6xI7t97K54yRIRGlQzxogGOKIqx4V
mkfU7yPuMUlZSTQZC7n3uiIwjB7d9u5Ed6JDMB9AVWJDYv2l24WeY45UrKki+iepXRo8ePp+Rryc
Xv5GjfHTVH4r85xVWk3w0K5wMlpFANq5ySyzWIZzzkBw87H/TbBDc15pPHmU3U6xFcQMOqgZvq1P
r/48J3GLNRRJh3n8oQiopUJCmMBjlXOXndrqSamXD7/mhrfW2vlReW1OP+UKS5cxsTUabOXhukkV
VQin/e5y3LtNKFc1ey/FAWCWHUqflbqxrhA834iOVNtzvy5+XVxFDUsTmpCfWHl+bSVsrZoBelTo
zYqxDPuvukOA26SnEYDQJkdwrLvs8XVFzcrYmcYbl+jnq0OHd/3369avwqjcAQAiRZrKZvoYJ93W
+oq7SYHytEumZuHB+DvGhwScw3//ygN989g26cgVOm03rjgw4QV4lfn1yzyWPbwPRZ7/w1aQwkFW
2XD5w+XaKloXj3qe4XfbWQqJjETOqjP17cEgksBjy8CxgJqUlADjfX0qYzUlIGQp14pXfzZUbgLH
F29F2n82dbWUjl+o9W7uW5DwomOjlJLxJ2DbrTuKBJ12AUA05d7JFmwAEdUr+FP5IIONMrOT1kMY
UQha37McynX2SH/CMY3rEvSibEt2R8fpiZOumGlYcs9ciCU6vzBcNJRXGh13dgK4x0IeIvBmLIFJ
Mm8Yjog0GjKdZCIH9TqxGf5WuTRKWskE2ieFf/G+7LoKMomr5wgrITmECWbY+867pJhURmCtU7Pi
SxQG/aN+NjxakLPVuxRSD6tBuoJok7wxR4t1EJ0TaWRfSBOfVha0R3dwuqXA538+/RPX4sDYaBkw
S9myyNDoqZOBZXRwOhpOsmCQw6rgIrXJyO7XZ7n+2OwqP+IbIDEBkNxQabIqleLty/j/uV245lUi
h2HlYGzcw3G8nCus/I88sWp4dMogd3Fhuihl9+5hRn9LSmPVYZxefHqaAg/E++18k77+xjLHanN0
rW5ig0ulo/TC+Yp/GdE9ZkzqSowW1DraOPgdHrgOJlVzMCVPEQuq8hAlvjKXPVThp06ekH3DXJzb
8PoKtH6PYVAgC467K6PwN34C/ie6U4QtwHboyD9FzG9cIt6aTVHCBkk0ZczE9luLGJ1MYFr10gnT
U6DkKvVZV6gWciEtAQp6hp92UJ+lCpe3hhWNT2+hPAYQQKJh9uZNoQcRCLScBGzNPuIsIVrZ1lUq
vCRHz22O6FR/pJUJQlL312upBu99Jw//YAzbhXYM1aNrMPk/CUY9jWIpA3XdY+WOmJaw5oW0zJxp
BNPn8rt2jxDeQhDDi6Y5fkfdRxx+jDmfbwnFSuzZnvrOyYyS2s7zUtXdA8Yko+WhQDY7bcMWGzN4
Hbxbcc9d+TOhEiUGOvsfuTr6v4TpCsD71XvkXrs496xdXR7ZFh77j3jqYH2dzkM2wcefhSF5JG7k
JzMK2hgd0tNFEZIfeK03ksISHA1B8CT9wWUGvAX3JBE4urgi1r7xrL3bR/VsHD6HY6OWmOkO8wvo
yD/TCBv0CzWpd/8MfML2ERrVG+AGZRvIX73d46jYg1tk7QuODGHXMJsuooiT/q6PROkPuQmeS6NK
K4sMSCzkNs3uX7pe8z4EsgnAklUjvhSFaI+sfIprM50LwA0mQETL8y4hF3a7+ncaXvt7c3RclxAm
soPM2UTGG+YIXjCRNNSQ8h+Sgq8umNCL4abJ9a0AKjWiZTrJyZEvhwUVrx7L9CXx6PCMFMtfc1F9
dKmkn3zp5YmInIL2fQyudykm1HNzlgitFeWt8Q0OoWp4n+yTk4XpG95D2lIH6aGz3zMTL+Pchfjv
g82fBoIHN+ST4f3PYQcgKT599p+hu9NAkZhAUJNDvtEy81cwUojfHKqjSFsc/d+FAlC87+aa/VHR
d2YSjXfdYo8mSMPDX6A6spfkBCAH1F9C+rrvCLpOlLLis3LkotpbCEY/IVrXnv0fo4yMeAZxlmrT
d1S8LumZp4a/H+734/BqbfDgExEfwxGJxc9GF85vtS6jod0DOEekG33knboq7llj1L9oTA9NA1O9
eldd/tPPxkqweefcnt0t3bJihLvOevKIi/IuKit1tbrsxMy14v2fkQ7gA80OAyfIQ1UsfR7suz0f
uC2HgD37yDWZlGD52IZR97aaGuXlXw1ofzU0GbXy4RJxtkgKYESVIaRAN5heN5wf22z2fNDaL3RJ
GqJEaFvgMK1j1ncFntyc0JzmIFBHvxLPRvpWKzmywuJmfnmQThRP6HRVna9iopRTb+uTdMTU+xuO
+8lCknv1iszhcRe8TC3pbeYrsGee/jeWQebUyWkxHNTIoYNYHiXYUkd95lEczgtQc1cubG1aOea8
DhSgIwwQwZoDeIMwqBFr9uSA7OurNob6f/7gzSi0H+8LzT8Uz6SUcmU0/2dOVuNld6TamBFKQPfB
x/wg7nvb6rkFPKxPhJAMRqmj7ycAR12/viTSukIEA1Hy7ov9mlxT3ge7r+aZ4wd+PVYCet5Mt/bP
+ec3Oh6hw/WW+r2DH0KSzLWDTqyq82KHFOXSP+laAwNHZec5G6BVKhxUjydIdp74cDLeDdN4LaXI
RaPhhOJxKHaLcaZhHc12X3/IRhldvuqNNFFkHvLCsyg9sYHZlUAyPc5HwY+fet9f0HKKWscKZi7X
D5iorEKl+b37C2TFxIvIYf0BDR99OkQfLy6xeolVPEnypKWWlggap7lrQqDYjq6L5wmNFkCMAvo7
+kcTpHOdFV5qTT0pE2o1lEKnM8Nb66cccycRLNqWuEq6HM5pZSvaZN4S8e9T3lHuMH+hv1eyiNjm
BzmRbyssEUD0J+O32HRfxrxJ0dnAZBEHaOzzwTw8fC0vPAGcoy3Gb40s3slqJlRyTLfCVZnu4E+q
QdUMWcg95JV9QLTmueH+i17n3fJGKBCzdNVdYoRttJcRX8rT8kEb36emA+XTqJxZvcytpf6HAyN5
9opXlUseq9U40nVKr7Y2VzwmJad5A+n4afLPKycpf6adt8ypDR4jcJ45yYlJlt1MqfrhK3WYUaVw
Onj+VOwrcagU+wKY5Oq01GRb1N01htyY1CHklTI0id1kqrgBU8aYkuspe6mn5oOV7Rk0IhMIiZJk
rxsMlb3lylUjOI4zD8dedPZe0GaLENVjCkYwtZj1u6jxTnbl5ZtYD/cZZFVwry2du9QBkRQe6qLX
vPu3G/t65Br0+Av1LsiKfE8gTDBputnwdqJiCOLgsgi79HOT+1/qcNvP+65FCDaPtni4IptY4+zz
52J/07rNMe8t8BHChl72cgzv57XKJMkz639082RT8+P45JZPytbwpWd40AsebyocG/JEdukdbodQ
jB2r5xnq/KGX9GO/OcGCVEvJAzdp2OydK2kumZGKJu85ckCsj0PH5NBbsQnWp8ByXRg50YpcTe1h
7uKgAedR7bOECyK0S1V4e/sgqU54t9AsP2ytLMDCCh67ZgJHKkljYSwbpMXxilaY9JuL4DtwcIh5
oDGyrdouzvQUlXWy8qBkDbTUxSuLE3r3MMkXVKNmCUzw4Pc4Pd/TDvOZ9YFau6zvVj+Cq80V/x1/
8NrY7Sj/MwNbLfZIGxsLrWjDTMPNoea/XeCewxuQlob4eJa4b0SmP6CEf7tn9A7f+IlPOwQIkTbp
x9tD/SjsUrEWYgn/K9xBUW2EPrCxdeEaB/DWMwprHuUo2JEKjRaBDvCO/+CXuBJ2Nkdasat6RSYL
0zocHhoEmXKidWJJyZfOiPYtlmiuIXa9ycxaW5hJt604acPx3zaH5quqoVebwJYMhhiP16i/+Y94
ooqWuI0AMJu6cI6oe93q0rkzUMX2+SCh/RlJXJO9gulasMnfffFvIjtWOF4Q++TwGO4CvuLai+bD
j5BwH9fImBShXBb4NwNqLA50P2WYXHRiOogHhvHUbuFKc7azvZPvHzvUuyULfpjSEZKx65TgvMcq
qiDHLBdfkVUHtkREevJl1wcsHj71MVCov1SZwiS8p+c+LGW0kKGWWvSLmcbjj4KQi+otyy5BfAod
adDnhL4nvl56gOhY6zK1baaKN0qqwHmY3v8FujZfzaqylmmAs54kkOwHqAGexj1fnNn1cjOY2eFu
ryc/spGnhmf/Q8i370GcJB3Ah6doLWzSqHAQTQSRoFlz5+Vz06iY3METSndAMhBH9wgpAsddu/m1
LMMCPwmTjNcQCnORolMiRNSIIJWd3AastnTBss66FpWy/bIitk5+2UIs5+lPQL5jUtuw9yTrvYKA
Q8ob2cMmB2HhcIapDB2cf5KoF/d0fEKDEElhWGuJadsqLCBkZDXa+7akxGP9OfO429yXgTD+yy4F
FadL8B/nHIbKnCMXkhgET6s00p5YnpldX+opzIWmj01iKj+W0OLHZUd0eqhNAi4542j7Ysn6J/Ti
UQKUbsj13B+ilce8K735gwSR4zi0j+q1Yq5CVBcbmDR8MU5FV1HsgDTqDO/nKrW7p7rE7mIZuddW
suFsNdfF5UcfbotvPAtJNereMXFq08aJn5sH4dxhKSQw+XqLpzK5Rl5QwnYLjCMt9HMb+Akz9V9V
KhXKSd5ZaNX9yTBremrnktyBXyD2n2/BAz5D7EpWgr4nm2lOsJSxZf/44rdpwDhe4Y42a48cKkKh
ZlwZInEpkqdrwp31K5m2DTIiH9qLkwvJSusM8tz//2JUIqhnfQ3O3360UFUSgZ4ng3fNr8zl8D0M
QZUTDCAd6aaG++bA0C2QRGoEm9gxIfjCcj4TB6RmuCfaofu5j04Xgz6SRkuvrn+7wKSDuasFUXIg
+nu93Dko0N0oGN7xf32RmvowKY6/wx/eGk7+p+uct/pKumYsReDMm49wCuifbIVFkK9DfEUxX34x
/j3mT5i1h9hEs07D7FGXoKuCZW7/FDBl+23HtpucjxUfrzwnnhzpUnoe+EYoZpHpdNmEjWLB3f4k
7gIzQMbItjZHNrxqLCDkpWpFKf0LqaiRkQ9aRaw7yAmf5PeCd9Gc5cPWUIHZXUCXJAaMjpwf86Fo
CWIvrGIjtYBxLmQc0pZd+7EGFUK8MYXjrMEYmPX51HVxZXbKo8qHb2iLo0438m/RoixoW97aj0PN
SN2bDA0HMHSkHu6dVbSsCLmaP5O77AkzRyM5+RUFYzB1kD1Z63uSo+D3ymL4NqS3k+spt9oQVkJn
O87a0HTJjS09M9rcHK3G5OeqbMefjxnmfLWXTQk6g5FstJeosYFEXiR8V5tHBBRiMyaCknlTD4Om
rN8lIgkRoZEGoKa7bLAq51hEk7I5bcboL/YzkljNfgh5ktqqpRsEBIJPSK63YemrNX7435PnF9G3
aSmDJxkhE5PEWg7Kb0nTXdk/JoNBrYCyJyaiwk52oyf5JArxYEq60c5/cHwgM7hrlTiZ4b7W+WBS
drfnQomWckNfFNSoudmO6Mm1wqO+KqYwhRW27Yu7d68tJvLbtCsnEwE/clVmNgLOdP9wEVOJRiGA
Ae6g0V2eqeVxkhKfWSEhRlwolh8rpgWsTArop7LiUXIEdBsWuFR2lReMhAb0wZEduZoK51p6OjWK
j5CWlAcLEgS1JurAck2s23g/ui3zoRqNXyVg5TSfzHAswTdMLI8ulVLq86Wu2HePXBP6BbJZYnj9
Kst4368jX/X5+d4BIK1lLxOmyCkvdMmdWI3K2gGrbu5LYytXJmj5ZKwJcbPCefoz8S0x8knzHcx0
/0Dpq2GxSNBn0fAiebXrmYtkK40UGVHe4HS3JR82h7bb5AI6zGv2+3u0dv8ltBxL5zhimmrEbGyu
BW6i0yYvWxcW6sp/KnYkghDo5qtjLu/uAetQY9MWe2+S3b0AYF+FfjAKVtgZw5Ev7ygW+sgNZy3B
+B23eRIx9VSw+rGfVJWvZ4yVSx7eEW2TAvZlEsYdjSrqq1r1zoFB1HOs0h0tCwvSqT4aVTlZIocd
Hj9Kfnaj+muaWeMqdLEyrjWlFJYsRjtefYVDXPV1MTvHHx7uR2WOqgGpwv0edN9wIuQUPYvZWJc2
kIx6qnSqeqRXmNr1G/T7uYQ8lGnkh6BiC1bQX9xEArQouWlW3NvfPS2wUqJLotasYPqrYEAyb3nW
/ro2eqvrtEUhkcOGhiCorW+iq1+c7r9lym0GoTdYGwhu3qmrFsNpX8y8bpwOonWZzu6Ggjhq+Sxj
sNHK8hPnMnjWkjH+FBQeFC5MCJHkBxcUT7Er34yonz+L864S2XADz1ZXMppZmL4OjAWuTWp8XJKz
RHzkAywWcqrjObslS+YmzNUeTuRHeUmG/gD5wy7buQ4DaCgOr8WBa+CI1Sz0sDuD19g2cW3Q0Awl
Pe5XACt9BQ5nTHmH0ASlsPTObrCCDBYFC6Kk/9iNuhLsr1T0lk0v97lu9fLTW+gtTYvC3zoON3u6
1p8Z05DAFxNxccDS3GqVgBnP6fGwPiqzUW0pJ9rZboYCSzd9iPgoOAEf3yk1+eRYjxdye6j6Su8n
KzSgyOZt8iyUp74r7/3fKpumOdVMpHzMf0CX04K7W5egtHZAALofdZb3YlVmwwAes3g49jGIjUfO
Bgs9/b5aA/pA36Thcut+zYM4VM3svNy5rQeXGFA7C0K2zbEOACkPHHb5ae2YsvUZ1ItNC9dGs/T8
HEQr5jYfK1r0eSoHOBoIjOQ9RVB5LgbQTUHa7geCqBlgdx73GY+8XL0kBqHeqNzzaf/IpB/9+4Sh
zZphRkUBWY8vrgPXyyDFrvcEfXNkvWhg2jVaX+vYzO5YENCpiz0L8MCsjCN6mCn+G1DWOs7dMktZ
0D3vFfaJxmKshMrMXlPqoYHX5zr8MpZC56FjI2zg884ZPzx0FXw2MgTNCFg1zx+60mZoRS2LthlW
S3kRBl0STtYr+bmZl7BHoLn0lQ/8Emuq0vAOmKmpQYIpF87Br0Ggd/9SG13r0b1802Pzq9L26hg8
1JCAKsEKzF3S3V1LuCYKlcVGkuqZ2ZXZps+sf7f5DGSx5Ggs8cCM8OH2vqG5wx4HRxJggBjVNetL
wVjhrgOBKN2QVWbbQ16HMFk1nKzok0rbEqhGdoxzBbTYC1+gptFW1N37jagNq9lzyucdvmJovZ7z
TqILmtKQ0Yz6T+oU0IiazSE45//J4vIshtnucqL9Ts2VPNwVZWTMFGVnpvHNxLV9BL1nU7b+pULr
e68TXeogGiV6ZDO5IMbaf4cZkMys14uHrwobNwN5o7i5n1uG1zmjlFdkX8QIoWIXSPdo2RrxMQD+
R03XepdIsuuHuFaXfxKWf9XzH+juq7mBKrhAAIB5JgIpnaFcJbCHiqAYsDMyNUQ1fa2QliK7fu1o
667jcGvhHpW4vrj/L1ghVipfTN6yiuUQmACkmW3plFySYM1hgsJ3Uhqnr5O/eWkTvD/sKN4tMES7
IRMoEb57k3UcxIX0OkNKLAuj8w0z91rjriIBizibchP2k6bGCf8zQpSJ+iCqA1nY3TgYBaDoMzOs
K7ov+cxoQ+TvCSwX71/cx2DN4Y+f4bdcQlFqO36Loz2LVMxveaEaVvYMtjFPgEu0WgvymvoixWTG
Qd/SdbF6M8hb5k/zq09IPYHZXnIQRW4aYLFlH0AI9C3Ipgigl9m86FTea3FpJ/pDKABjj3rFb1aF
hKsWTbJZvgunsuEae72XQ9lszUeGUzHh5Me+fczvo2ZI9WyXgf0hrT1tAu49ouJHkyp3Q6VdS0Kg
PmsP2+wclcMgFy8L0v6iXXLYPr3azvrlSWznKUyP4QcREevSZDG62tUtA7MECv+he/KRLljFLqcA
Ttq/LWoFlt8VT2/4tUqF+9Ab0okFBQWB5JAI2R44wNn9TEnxjd2Cjw+gCAp7UAU4usoNGtqrRk0v
ykt3UrabTTccn8+lEhnOEKfo1L+Ck6NVYxcL7s/uGT13MIuPs1o9ydxBahoB0UHifRYTBdQvA0/e
sBmtX0GOuTLMKnqXwzgEtT2Fue3H4msobhisUAhQdAQ5/XX3Ctc+rPMc3zjn3n9R/O034eOBuqPe
VWv/oYnT/riCVCqPXG3NhvSjUFmi6VUPbsXTQSrjOjRS0KN7FCbV4u57miv5xgB58SvDzjRbtG0/
eXVwKr2ajBKo6Ib3JGzZV4ZdMnYy14W+XsZ8/ZP9rAslL7MTlNKiMFTbuIhiSLQrRZx3V0nl/owg
URxELi2EWYTLrArgJtb/9mHsbyFpIia2EI/dugrze+yU76Kc1WSaaxwomBezAzyhd1xGkI3SsV0V
W7jA4UrGC/owUH69heZAW+KKzaPMc9LPw5dFvJ4AdzMeae9dy+loBtrWtD9zB7mtnSnHT7s3fkao
YNk0JuOofTs/1UE/l4qNAWGUcd3Js2dRBeDma/ivmLykCdQOsnhc2ljWKMGIxwQkVxGk9J153BVw
Hi7KKw6oBoTOpOIUQSvxr8aKURFnIwXazxzBWhq+H4eZhb79FK3iuGe8reMuR1F+2/p1hZ++wwum
QhQlGIcLHQeR/qTGSqNUtr6QrnJV8ZyBb7CpNce0wk72acY+ZDccYnw5zstayaZRKer5r7vyewIr
lv1WmEUr+HZLP3UAGh6H1luO4IKKE2+qzK4p9Hh1KB0Cw41Yb+uRezPeIAfw5uXYCLGy9fP03zwv
SYJkErBvs3V+O4iMSaXGUQpRpyI9XLEolrBAHp6t8g0nQMfDmYbTU2c0QqUcXlgaG0G1P4yyo9fY
axNPvHFXBTdoEUrVmINOAPdcekASDAgd9i4F9HbvTi+HLTG2P/AYahB8k+n1okaLQfqjSHzq3wxw
l9LpS9jUvVol9ECVIUXf1UcMwp5cItntYXHWdm5XxCnehJHSs4kkuYPSDM4oHZukm3QWNXtScTMg
5Nb0hlspYQX7kN3gdkGkCboiIEIwphzSqygJeyDDb41rmOn3EqwFyp+a1X93i1QAJAfrpKpBEYzb
9CgnEeEzdUdMgW4oavdqgo1Cuie0X1gU8wUuNXZpAQ0CBeaptDc6oBvccKsXbM6zQMe0LgtBuMFh
iwpfItw99g96kSA4lWSMx18luMhrD9Wuvk5VNXmsm23Fd77KRfgXfSJ0zVENN4/IOf3aCVZsiJbt
tAZtuLWAjcyOl6/9HuG79wpcWv9ONcQo2EcWbktydRXsUlwQfYugQ4YTytXvTOO3yh2DWXpvPRwc
ZGyuvrwG4v69OQOcx0vtCl9os8NTRLQ59o7nWk20O/FMYYJRQO9SMZOK05pi/MP2KapB9LuCZ5qc
mpX/8wTcnh0KNY65BohPPdNrodBqdeM23jJ0tDe5kRf9IcHTLCu+KBTYjZbt4h71+jyW1RQqsjZn
NSGrqXyzS3mT+Itszp2KEMxBQ1aZJ3JsctosBk3t0gwPa/HNbBBHmADwZCdelIKEdSpTOFulcw1b
uHoOSf1HtsQcC8BYJ8QD8AREO5Mc1trbiTO7hhiu6P6WWY7SFaqdYXv7SDehehr0ZNIZXcTfc+Dn
QO875HaEAfqpsRqjA+CsfvAzR3nOWh8o2eiB6vW7q0XR+dJaTPAsRQ+mLCd0R7Tzzleb+UjWxobl
BdRNvwPGki8wQ2CjRjNZGj6qviADuqbYTcpxBo0ZpxWh7DrpTG8GZzdyowxoT9WujcnRvi2nfGqw
fRQlZN8I6oW5yPSAh3KNIsl03cbGijyQCxoRvPaOCcBDALm7/k57IVsR6xWRdiJZZARX1Qva3CxG
tlrbDZjy2qVVN08O4CVYt1CTLTxq5GdaQK7//nnG/O/TRx83EG3e7ne2XvUQn402rDOsp8Any2vi
ikMpqfiYe3wmGaSIDKgxZxNiyRoRkEUPXm0ALoQRYHC0bU6vOxG4GVcujRK8cMRpSDpBCxFEk+yI
hYd2XuKtWZBoM9vo03PuMtwPEod1l3njuseEayx1ziagE0+Zf4mbw4lOqUwvR4/dIQUs2THMRBeU
wiQwriA/kpJd/n5AR9gpI7put00NvjXEPgWh1/in0GTCMd+aoU1cHdzKVjy24H4LmXKRhoGMJxdo
SxXmaZBirajRI8UOY+tit4L6D5lzCBYpC71J2zWjlwQepEV8lbmSh3Pibm2Ag4NMgNBpPxrKdpmo
wmFD0L3LKAT23GTilZbuvC4VnofVOr49fCtht+CDyPTcUQFTf0De0Xnw6xoct3HyePmTBYhbkc0V
+rnmRNdE4UPnUToy2v221+6ScZui/oav7QPp4tDxi5oB1mEKWLXLidycU+QptklpzfbE7KunIN5q
ET82veQOqhwtuHBTYyw+PlZfWUGx4plUHJDYP/96kSjh1RBHMqJl7runHK3z3JeAPxsWgIqGfRFo
BIvTgWUmojJp94J+daLPcvvMSRs2UbE52wehw2evQpg3ayp1Y8lvlAlQRhjWBYWWFvlPNamjwBAf
JcPQXvYvHEvoGdNM7/KyEYPgB4OjG1G9FDCoufFupzhCxfxrvfmhjmiArsPVA45Y7qOa1ZKzmaC1
t4bhRLXqrxG/eE0fkkmiJQPnpeQOKzf0yXErFJmWWYOtlR/8SP4Rqcu035K9OUueoeW2MeV5QJEc
jU30yOtqUIbbxImsKf2BQ5+8Drws4WpHVnWfW0TFgdUId84cI6XvfoHoiWsEvCLIW6IG510nizwY
Arzp02BIDsHLuItRfF+WlIFuYhruy3nF7BhkQpw/29vsYDCgaqbpCT/2Edp/rqfdiena7w0Ge1/N
ZcW180MsdfihFNLvXrZd1O/Vt1dmlp49W9Rhl0ql9XKLJyhXfEWBsoWa/RJRHipbYQ+kJqN6Qyze
xdL77BILBoXFxGUxe2ZLk/C2XZFORzp8sBm4ISX/t4zQl4p8pvm9fz+ypHhwXz4o7h4Gf1pfhSkb
SDEM1kxOpih7P3PaIs4hVUAm6NBtYI9iexgnUs1SAvuF8mX74AKhQnax1tWC04KYuIuJXHh8OfSy
vJsICU5vZQz9Dki5sty9ipVH9z0K94KNX+5hiZ21Vk65Gjs7WRwkxLFUbXUSV4rO+hYJgW6aB6Kh
N7GrjtLmALaif5mzcvfLf/cB+DMM1S37/aaNYwSHZ4FfJp1aXIWLuRhcXx7KFIk3npSHB+fzi9Lw
9SvBq9Jkujw3Bp+uKJw4iUqTeLQZd8Nu2nz+hDx6vL+9PvojdiZOU5fY8s5sKWAnrOmd+0sRpFC+
z9H426huYVb9bTdCJXOjlp84LTVKjv5heVJkzLln6GlKKzcnd/hyC0vGzNwsGmmlkmGtirLozJ0+
/zN8j62/5JEQ+rEiL/ftpz98gIsmUnD/YN07v/KfWvmUyYkdGOcYYKkmyciczvAEZ3gvQWUyuAVa
t7lMr5FiU5fm+aeAWX8//6l0ocptBwVawEyC5rfz58w7u3Eo6rf+5wtJnuW3GEu8sxIDuEYSXJxq
ySMVb4t1lpj21vI2jWDoKp9ET17qjAUPgJ7HJgYvDr1Z5WT+cpHhKR86iNjTkxrSFUgqkCxkvTjD
kXKNvBpODtv0v3DNSolwKBE3MUOybXEl1z/RnPR8CoJ7TZS3N/8SXYq6hN/ZyrjpkzGQq86UKBr+
uB220QPo10LKB9yMkDlpyQZuIN0u/TElLVRupK9Y7+ssSpIVCnLLxeM2okyOmxtSdcw21hrhP7Wy
noy5KjLWeqRrWIGQbqYiE8TLFGRK4dltHXXkQidrXpNMLz1Ny0RWM6S1LGK7m8fR05fo3LmCv8dI
uVhAkf/jeEDJN4jSdSI0eo6346rG5J8aLZpPYMCT1yqVs0qn6eo29ZMjCXyp/KENqm0MpCPEj3iM
K9UbV/t9BAxgQ2at+C6XuOnHGaPSApHLXvfoyKhia8PVV0WtcGJfKb8zwFo4eyiCwhSXD9ySNF6+
3gSt6CWJRlAvEX9B0eYchx5QBRYn/vkVPe1w3wOFneMVt8EJdxf2/Nf0ANRG5qmavZLABbGeRB8R
KvfGpdJbX9ijujQHLGhthRS6Pchh6s4r6/Cq3Hqg5I/Lhtfnh7+a/QSL0+Gr1a5iS0rUPaSRgIRj
DQEv3sLk4piX1u2Tz2vxnKQdr22wCCEYxNbgBPPoraONhKgiFDt0CRptLFakGbcgnuMVdln89+32
SImuufeoUflXK5Lft/A3PK8cMjOVKYcwPJL5KcOUo4/rf8THuIP+s2d2T5gIgjoBWZiYrgoqY35A
FjDprBr5ChZ/mXHayfGYx8JuWZrBvK7O19a/oXKb0xrtZVJ7cLKv4i3sEAqlVWAESIMvq0dZQDst
mbSmSx45s8va39xW/K6MoQ+f2v0Djfn9ATJWUxC8i/OVYMrbYCIWOtWmagkX3Qjshgv335Asoiku
jwoByNgkpN8zlrb+reW0NO/IbpSuEzk7gT0CyxL3wW6vIvJ0gK+shjzl+qoMWylJqWLU7mLaQITx
HEpjttRKL1ZXxzbCtAZHShzGnoC6EyQFAQzGXY8CrGUDP4ByB+3VASS1Ul0xOk1J688xFefFz7ZB
Y7g/a5KZFVCQFoJfbzNpDamv+GCnj6dU+Z3ho7MhR74MDMQ2W0ebW2u68szE/HvHCcCFy+jMIxWu
mJbdyhlaAyewhq5JyuzRoUSB2nxkNSRGXkLtqL6eZg2ZzDgQkx2c4cUpTry9J5ADPaVI647ruirj
iTUn8y2zYWKAV7S23aRWo9hTsSZW9Ia5jrcvA1Ym6iPwjnuzZOnXebF4nbbf4f47Nj+XhGHHKMgA
Yz+I2gbFUfaA5GXCgVa7NiNrUav5EYyeGklne++BVz1MOBPX8xrZEWovKlEAmP4NPvCY9FNiBSLy
TW9Z8NbgHPgCOtWLmgjVypBQWQIt946F+n3N3vMBJnAukrzcuhSjKn1g8oqjXwHC5l7oSC4+O5fw
e2axrkXRIcS9I3z0acZ3+frHo23QAKNBlv/0LjAvEUePS2S0GGPyYAh/t+3+Pyplfoh4/VyC0Qie
BMnji0EHfT+BUE1jIILufcz2EZdeW1xISnKtwfPsa6w/aSDcLSMcUj3vguMUPDS0GMYS2oTKFe2h
n9liPUOkbcE61gN5EJ+Hecz1jEyV1Fj41IUoavVod1J5Ay/gJuSONNX2IExpkgwa+6VMHF36C/xs
vXivVLLprJsvtozBrd6/xMuF7YyPZC8hWAU1ctVLckWhUS/Vc80ZUFqSiFvmr9xJ+lbyufqgKiJU
NAwrJxnzurtcIhj970fbXuOrlBmcQx5MOL5MAGODhzC7I8wV3mmKjIEecriudOHy78cr88o9xq/W
OKzGngPF/IIbLgb9vAVfDw4SZmQg4B93zpzcBCTkGkIBWnzTmThvA2Na+YIuJCAqAh+g4QKHQtM1
t93XjT0hZd2aALJfFLdAAm9C88l/on0nnXhS2usqJg8E0J1pUVqj2o/ZTO6wMnSrEIpLbKHwOfqO
dAYbXGlE8901z4AFSjfW11ZxNAyZOnDiSyc5zPq0a1IYLsq+NlO1kmXz2ulSWNKYG4rHFJPKLHeU
9zZXQ+ISgavsI/sPgQkqMwqii2IsGWrS8lLmY2EcmSeQqY2CIFqC9D7u2M9F3tpHjpzW1h0uIJ/j
giwuubxHMPWhwr4pmn4kY+viaed3wTt81F4EhnwxQGEEQNvyhpcjLM6Do7pinL9udWapixjFa8ya
Z+8CwTn1c/jKYKfFeXVeDZfT9JKkVetzQWmqEdK4ScbJzjV6qwfAm2Q5K7FL3OFfxVvcFDNlr4wq
PaSHiGpcEBjWeBBwo28i/2laU4DP4REVRDWMy1nPDJeZALB9hVUjRHXBnVUb9MgvApeusXOVg+T9
cRi1npzQosRUee7AB1EoK50Fl6cbg/ZWfhi6jTxJvphoFtN78Pr3l/y6NVo0zqHSVgeAA5QRcz0t
skQO3ljy6S1iveyaQSWpQyQSsBracwJ5/4RcVMklsTmpP0KBWo87EjVOdEi8Kj01PO5+UDBSVzeJ
8h+UAgrxlBTcB/idHu2eyQD4+QE5cSd0Nf1yJolI5SNkzxtzzBMxwIIsswVlvg2A46D5N+hTs7JF
sRM0UAKrG2RcyS8SsIX5LIORUA01LrH5XvMzbAaMVv+6WURdni9CDvWPey9g+KIdYzoFRefx2rmY
D6VUk13qOomsj/xIjvVSzUfenni7kdBuRYIpsdDpaCg7QkVnEFRNhQnrzyqaCDxfOqMk4FIv0aRw
7ktvcY+hjPmI0fJlzaa1i9emenORSJbF11OrvFYu5BCphUZKk0HEAiEcDaQRDHp+H8rI71YCOaas
3DGyR1l4HzzuRpmzUBDKlrfrkg+D4EYkBgJ6nxpZN6YVXON0rSb6qBar3qwRN7ojs5V8j+LCKAtN
vqzaNfsv2ZiHC1YWn+YnuGdqoDKB2ZXHAuyA1UAJz2iXtL+aC7s1JJQ2tQHxZDvKiW/8kjnWiBBs
B3074sNf5jamv02EvTWRHrLAn0bByqdWzZ2WmjCiZTfppMnwpTvQng4aPKddZ9A/Of3pY/fANzG1
jNTonKGcjsaPnvQ2DbgaCoyJ2omtL3EIDw87zYJvZWuOGB+/KwKTF60oqPCeKBgG9v10fOX2mDq/
NJEBxAY60mKjayPkRJ5KuhOp005gYWuk4vYgrQnZe88ZvNoPejpJH+vUkVBPMigNTzt3UD1YcOrg
pYCeqlnOb3lZmTWqb9K61DQHjtJDWNpmgF42ad5NI6It122OAaj0DgoY+EhISw4wvUdgOuTJNDCH
yS8vHx+InZ3QSIzhPLYj9Z2qFsyZk3jHK0raX4yOGTRAUPz1nvg0fLGLKgl66jKQVLdhFfgpdT5b
zF+DjP4PhEtTiIxDSBzgJiNROZWCtMEQfHcLV0L0tZArHn6KDh6iMxFiyVdcWdAqM1VW4ssfj6pz
m95WDYUPoLOI8bsbAV3wNT3fZsBgeDBAMr/+QH0zmK11Rop9d13d8AHU6lg46GwWyu/IgfCKTv/c
EfWzjM2X7+lmo3jViSjRUvdo8zmzT5CAGjz1jS/rbI7NYR+qyKurBoiHrgw79M2TNmeR/PUeIml+
2K8c3j6T1YyethsGcKnKcivm7V8gNlCPWViHcjIUmEsUaopTAMuSKDQX+9W+wxewfzP719IBlUhp
X/E0esRML+Z9h6blb2FNQFJ+62SkR/eArIZa4hsWBp3Xp5BsTopFaQals9Lc0ynV/H7vxhA1x6u6
aN4fDeqMEmJrdYPjbDId3S/pxLfAjxfZSXStFSrNunXMKxnClH8ZyAzssB0xdqce/H532yNV+FZc
zWdS/MyyQeLaNbVraTvbftVRTh3gHiVnhNdtgUnS+clnEBnw8RpFew/CunYAXq7U2m4OifvXSM6D
qQeON2ETzIRrGPpWiUTi7+HagZPUSO671qhw4/kEz6XVouk9bDWG4lGNsoOGLMWxgVyCasqVD+UX
luFgWlfLwjEBW2iGxRGn54mSoP6/D5W0Y5QEgeqcMIJSIsVc4Zo9E9Kv1MLQd4IiNFveeb46oLna
Nray34ffpr3nAl8KNj1l/bSR3tDmN5I27Z8lsQ4m8QYDL+8dBWNRPSuFu9SllrimWWJN+/7E00ET
l0PSw77K/GsfrBphmX7qdWmcGK4EFy9Hn2H5dVgOjfd3aeNB5xnbcsQ9zhQUPvTKdDnkHDrkXs6z
5z1OAAduf06yhaPOM5CdT1nZ1PEQvU+J95sqFEaomyFEZqOy6CQJ9i8W3U+YA4Dv7Ci0WgRrN0VJ
ccHArz/DpPxNnomHJ0/vwubwyguxDSLayQ5zvMmjpA3mWvPBK2vP8t5ahyEFG8+6FDOGOZ2FONid
Lczgq92Iy7ko9sRB6Tbz0wPmyGCo3Iit5OBKmKpIvmg9skfvVRjeqLRzS9LjiZVnN5WplzY3dFDi
cde13KD5w6cTH4G6+Ew8y6i3aAPM+s353XY2Js94t4uprneuq4dHqA5bqdn2mPwzI8pvVmDt3W0V
l1Inxt9BXrJDx4vNB3zMtQv6NbucppT2+l0G9VvDojV9ieSeU7mPt9+Dm5JhSsLgoHJgB6Fp9F6w
EQh1kZRDJQ30pRQ49GHLHiAXePiyz9DdOPmvC6xB8GDNLNpa6OJ97PoQ7Mv0SLW0FpFBuTpXRSYI
9L+6BMPYhQtfaNm/c5cWChIToax2Lff58QJ+K2xuVm+hCmq/fGVBuV4Jwiprj0KAfrvdboljYCj8
cAdV/oNd7oDtd3gsYTSS3+K5JTqN3mVj7ycT40UvRfGqkG+ivzZr95+ER6eqU+dU74io0bmD+SOO
JDEAxdAJk5kx4uIGpP21XIsBSbofA99X3FsfJNBc/WZgpfAGAGaiDRy0dzzTK0s+nPfIa5JzyBRi
/vkXeffGL4aAq554pmPrkKVcrBVTYOq8GEj+6b93fReh2Z+j5TjpmRA1paapbqCH15D/JVvurDUe
1sZQy/c8LObOr3KAQCnaAHQSRke6e7JLo2MbH6iPawQHsfoZhyHgMRZNhtLJ96ielLFjG+QUa9Y2
u45F/QZoDZcH9HWGa1zcDqN2SL9Ed5s/ls2BbIYxRfze+oNytuIl9gYdtgdnmoFjuCuDCSDLUX2x
50eiHcl9pXS/S4cXo9DPvyb9rtOrYKubSg3llHc1xQiB+hEM6xGgP0E1vKZGlRtppbGDp7DUZi/O
q4C0sntY+iH7iTnF2LnBMQdOxgYPNXn+5n3iX1hrAMJMOSl2ttRxktS5qITajfy+AzyssFBOGZBE
CpFZHGEnHDoQhScVRhj+2VPLY8719QxI2X7yj/iQAfNrw9D6pI+t3YOb18x5aPgVXRrip42xpb92
4fXxM1PYnE8sTVssW4ugEY1GLLLyqjtclzRgP1bF8wqwFhM3YHcMLTBQoX38jSJxvl3tM25Ys58g
FartDANNuvIaUAMUc53YU08DroqdBRd2RkGx4uIcHjtmbuzk2Wgq0VBnyCalLsS9DS3w4YeVtpO6
lZIjYcl07mFncQGd/5yLKomkd/7kDWsJufxSPEmxWKmu9AdhUslF2HSX95z69t5d12AomSks2p2L
KAlxqzdl2lDnlqOaHtPsjTPaN+RH8Hs4LXigr2kr9jybqPMxaDGKAmtdEctkx5okN1AenxOgWIu2
GBms1vJ4wgtJcWIdImC/YTtUUco7Okp1iBIf5h6q9vWjcrfD2n0veTs6XeTZWbEvA65oLgd9cqE+
rfPx811LmoYRb7ZhUEDHNWhRZq0wO/W/ZiJVUsD4BUnSxSkzdn9wqZAvW/wRPb31ji7A4X7Nsyql
9TyWQtFQc283uqtMtqFjp7TNLyMbFohdlaPRDPERcwO0J5ZJjNaWZD6spRXep2Wgrsna/HjK/QPc
YFtvHFAKNuKYv1pCKxmynQGG0WKaQzPyExIh6gDDws3X+sAFogXzOFxfaz5djPz/FMog9VJ2N/kM
8vHCMuUnSNZouLFnq3relVkrbXR/VcLgjlMaB5SxwsuJ4nZdo7X/XUtqlS+/Abd4akSC1CBJx4VR
BLOMWPtgrWhIMDVHzpOgAJfr30L3aTwc+8gIaYfupNucnBdG4GVA1mMoIoGy/ukYK9/2cbhqPxgF
rkXdhZyBTgykUf2A2REl9Tc1rtSiF2Fo88kCaO9lo+vt+USXIMIJ3yLhCRm28SuB1kisFysMl2+J
z3vb6SMsIg25l+xocvpVhx2VjaLPmeE585tRunGTG9pliCa/+93t9wQzkZqwtq9pQnXx6HUb3oHm
QWIlyLVTkfj0afWnxaVLj2//MDNi2uHJQWA7pXdiFuPThtcuKXkNqlAAUQYIZJsMDY06fA2TZwps
lXdYWDDWcEQbG/Cpl2q2gZRAHllSdAGKWUnaBzXXH1zTrgVxza8pRO0GfxdNp3fKm0RX6HUqWsMZ
hlj27wU0u+OIUZzcOH5JwQksCwdCque7D1Gh5Sz5IB+rw0qIpTfxizEiEkxXB9+E6DAIZPnXHQ4j
RfsHcoDEWWG3bJZyVwbuy5CaUS3z79TwTX4p73ISp2+Qx7u8oBjrDO48Oei5QkKY0yUEAmArUN0K
koGewabHGPx2d8r0Z1QS2jSaqvwPANijwKpAbOKLlianiMPcGFSdb0ypFS5PQ9nSu5GxoYIdiisF
Fi56ICcm29Kuw9Glf2i2dAYyqbwDKYfJ0U/G026kOvBsZXiAvkoxVoojBKGtSnivN/eFM1BP62mr
yiHrTXuy+P92WzILc9JcgBSV8kT0BhWy2wIywbaN7AQ7j1M8Mv/+J2yidw7CJ5qS1cucQSAD2Gfp
8LDAc6fRr6n3HxiB40CGuURl83MXt3pb20VIQ61Lc2aHfsbdOe2BKNPG4YC0vKwDHnNVXohLCDQc
BTeyyRWdTV9BVbKwA++YHtoI+BV3r8KrQmasCbKLT4QrpE51MJHB/PB1Fpv6IzKpf7Rb5BVqlp4B
cE6LKakwLEUZuA3LaWlIJlFLcCrjDM9gGM82sEDo4G7cqZQGYDRWFAc/xDSLaef5kQdmSkMPRJHr
lQmLlRhVjTX2Lw2rC/mbT5258xsTS0FkcLU92HL8cS8jMsdQ0CPoodRdGHvog5JxGhX3fgegWEuJ
9GhyvezLYZmpCWkrSZiwP6nGV/hRNS+twA1601m3Y6jqL7RB4ww1B1TDYFBWiyFVkoJjeK1JLd7R
aaK7WtxadD+8mdzQiRQEiEog1mINVHqJDgSPZw/u9AbhKwQC6s1WXN3hxcQomN9FAhCTU9KtvIJE
sQc6dU4dGSu14LAsree5PACCvgTtRE3WnlgSvZf7EAtLKE6SbyY5kLZimNnjVyB8umz987lqaeAD
23Ttl5/CwrRIWBQuOlSHZ5uTM4eTEZLzqNYmlGECUZq3YY63O0BZhOuUbfUVyOUiblH+muiVy8qG
onviP94YS/JeR4QhMlIbeGBbQn3tv6VWOpiDfxgbXsrZd4vVxjohvTyI2NB6wCHXw+4hfshQd0Tr
i1qEdLPpf03Gw4nG5WZZGKFGQ2UZahKIT7k/BpjNJUrD41I6cM4qiRJpAREqa+TaBWGPTs+T7FVI
IPfokPPW63+T03Ae+p85g/Nu0/HA0/6Bm+r2YRawnib931lAQEyxm2LbniuCi7q1uRRcEz4gIqUA
fDL5w6dapqXYW97EVwhjQQtn/QzIJ3qXVjLo5UmcibxqQfdZwxl7K2H2xhwOQoAM7aMjysK6jO4r
QeEO3hubRDO0mUmpDtMRR3xZplzUEH/I34rC3nR4ED8IuzlhOBBbtV/8A0qPAoBpScPum6vm+lwP
LiAdy3UIvejp0Mhq9p1HLJmrxIMo28Qo33hAEca4szyxys7t4qnQdmLAudQ1j6S3eNw/t/QB7N5L
YbiLxG6TTaXGaMg2KRbilPAQbzpgIiIs4GbaQU027YP/AvoKYbefrNZ/NOnl0GhXiwlVuEVkAfAe
Unu/Yky6d0wd//aeW1oh7c25jQYcX/f35Z3Fb0tq6lKOQ+jN+Wb9i6ULkALp252t5WSqc6d0Tvg/
tR2uOBtJwUyUMzVWqESoMhEg+O+3Nr8yf+6YWKUyVOMLX4o0mVECi95lfKrdF0GKnNoOZmFXNiW2
axv0IttWotd64jdah7UGw4fURmPKm9GEeHqec1eREPGOF+IefWJj2JCvlFnjY0LiVRpJ+uGSxDf6
QYDOU43F4IJ9LjSSlUPUADagO2lWu9/rlfMXaVOi53+u/COEaBYrtBiVfcnZbPBrhBCu+ahtWtKq
Ap9Dn1PQbAowo8KxFHr79XVhrYxOnm8YFQtfMaULEszq/boJlSImwaSy2YlO6wgaZXTYjJYse2K7
Kwe+CIwqu3EgjOcUdmUK26gZT8pIZRIrxRFYQ0aBCm2aXJGrbkUTSNbTQupee9AcawSNLPkO8xIK
MKVAaEf4r3fFjkPXCGQVKRV3VdU23J1O2g46UoN0xd6zAU/Fs1aAxXlmg/MCFUjeR4qmEGXlGjFR
sw6gubYqwT7yXL3De8ZLhaCB6lTJp42l0tA7o6ZAZRoP8SYJIbFuLEHLbl5oJB7Tz7DRlsT7k/4F
AhYEkLQmjIJhzGtmW6AnlXGBT+P9MM62EOh5OIjeRTnkhqSTYWTUsYjANFSridHf5ueT51+bnT0z
ZMfdr5mWgE6TKDDWjK5P+5ARdljoS1Nvfp9LMNOkTJB5ISHEojneZ4w6qvZmhof/On03cquM+Zyc
WQhH8X1G159ftYinsmlG5Q4cm73AJH3cluFQkzXMzQjXozERbCmjDuKQaxrlrLczSrXxj/ptg3HP
UBBo39HN7LM5uzYW7mtMrUeccQXSYEm/ppoydL4vx5KemWAPFyAbPVCRw8XoiAxBgDn9WqVZcAAe
b6gvjK9qpErIuMMlyww6LlwensOadBfw7apfYXHtoCm1MLhN2wVodu9X7VisOVjFJsKDqSQOCE4W
8GBNr/h2sobm+YJ3htGpAE2CMZCrQljduYZ3U3PaJJv9918i7t8fTsN9DYsj2+raYqJC/I0LKpnU
mZYLROaI7jioFBN31hAn+HRup4WmVf3+6qwLDdaYLJteYZ5ScX1vpo4J8gHttvU9fAGmr8iVwEUI
Kl9T/tf+EO83UJhmk5L69lBXhuud9NgDGOcQ1rIrHvvL5iSOeQ81/LyXFAZ1t0g6Ano7uZOAiUup
uNEiNlwTgxvm7utI+F5Ez8RMRl8HPVKMeME/9k8K0/S4LL8tc48OiEkb7phaG7cYXaNEEQTFtbND
MMzNatHFIBLAOIdRdE07NpGdnvzqDkg9dlbHbfJc1jOEb42JXCBNP9Hi4rJ1p9eZ+Irul2X4JpJs
jO09VUdh/AQNC3d7vsBhRI0uYtc+uPC2NDRnfXSq2EMQLZ5SXekJR/DBBEZhEfizQAYUtZHJAkmh
qSOU/ufQO32pmrMtWJ99nbxODuN1f2O79ecbfP1tF25A5GZ0QBecFxoaZ/vHUOCGObx3g5KD98Wh
Trb8u/LXpZKZAd5hogorMLg4KMmpttQNVDUWOFlGeCZt6UJJc93zRIybEmBwOGCeUDS/OdukjoMw
zaOvt6QwhuDPdrfPv7xbvzDHLiZP3wkm67MY5IhmsRfpY3Uy96/cpZ9JKVtiNJqPNgaU6EHTAVpS
xbV9r5Okylfpq2IGJdBFq+72ChBhrMv74EWpApneCUKgD8/dfrl52lgeFlMZjt142lOrsUiAqrAU
FcJm9PytorObinXIczPf2piMw7pKyYdbTBwB7KCag7Sslgp16dnmGNlpmpsxPPalT+V2dIvmF1WW
2HHNnqwlBvUtlQjLqVMQA5hpBImTtzf37e70n1MrVKZ3QeIh2F3xyiCuZssCFIRRGn5UpFroRQFB
rfYi+BXpFvofBo3KgbOqG+hDsDLFy5RzeJiN35fx4vBaPNo/yBjxCD47bnQscxWLLmZ8CYM+2Q5r
ldllTM2HbWJY+PDOUxR1PRuo25JeFdmNree23vCMoqN5UZK56orxMvilUFuV2OOhO3ZYv1usIAvl
bTUBDF7GOf7pflRVB3jxkG55R/44zDz2OctYWC7LpPLWAT/VFmOsvjCkh17/9zR0jMR3bdvYJn1m
Ejkx3SPZssxOOzlvgPw5UzfCNOC7FwX1QPcguVAp6oM7TMZcgrpopjduugGPxBcuV3fjFdji/4zl
gN86JDSpmrZWvNTA6WD7uevzplRXVYr6aVTVUdqrIZm58dgrjirArgcnu/mb0ckyX9wCnz8S8JVU
xcrHdBs7/G59DgApaBEnZiZYZ3Ph00KPIQpK1tLAM947AxXZfVS5By/zY7S5Eoc3P158XrYhe5pC
49IBqkkxDVNdPkjbiyUbdOlHCEnNdiZRuI+qrcXMEJ9qaVyx3iWDY+y8LKo3NDop4q+KfszLpEMH
zxSgv3UUrCmTc6L8UfIftnKwcvDW3etz+SL5NvvsoP/P6oHx214EGtr2KvWguAp6wPU9D35OcBMk
1iEvQd7Ihj+A3Fp0PVMxFcXM7Uh9wIZu2TbUMJmEU33Ys4ZSPVYYsl3oa4prFs6/yjeQuOb3q3aV
wo11nClhYjc9XUw135AxOaX9JqLhwPYrXNqx7T56m8I2Z0twkQlx/oY5Hef5DprgLlr5bot38Dk+
Dvnn2q+RDBRmwDkND/wOoNttcN69G21d7Xldykp/ECbhSlb2Wu8Z/QlTR0q4nn8xS+NnVF6TsJbE
RH4scSG7hUdm5hLtIziIvzwZqbdd8uOqgUwMnQuues4nGvwLyqAEd9fvLUnsuZV8f7Lzgctphzie
Uu2jJHjpE45H2zBxu9ABwbAd+3OEJB98gwefORzHCDqqiDVr3atEa4lGWDglJILB6cODjdO0CciL
nu1r4vOk/SLSjwCgBMo7ZD7sf5zvzNgPLbjjT1biBrg8g9QKx4XiDTLydyoPAmIH7KoAkxE4cFMf
vbnywEC2rU+O/phuPwoLeXHPTSH4db6BiVcXsLqk6p4PZ8Z/3ZrsSHh3kUJc8ZdAlJxm3kaJsO9D
7K0TmwqMktM/C6R7luDYrr3yflD081qRCmZtfrrfM1NDV+GN0qZVZ1jackQIHWe4wJHciMpY4+Z3
sxDcXw7bUFC1ReqpRa32pqHSj2inrlNxt5OWa2LgICOVjYrWPiTYuNefUPnfNy1gOtlhiOWCm4rh
bUMa0RlEtO1lvuCT8Dbmpyi74SGGmgJ0mkiL4w7weHdihCNzO3SHw+VA0CP3SBF8Ny1nRYjyNBob
BGUDOyfB0qvqmuf5ZZRn84jQnekWyptIw5+DUmyVmn7EBdMeAGS/bnXilVnbA89csJRQTqLGipBB
ZjnqBE/xBx38+xhp7kyGlDGt9ghTGnCNuE3gc9oC868nWBX6BgK4q1maCGJrESkQebbsQv0O9tqs
Bq45dQEj5YARB9fSuatjPszTl31GNIspBD4+wQhCcy/ZD6olt61OC721wOfWzlmiwTyyEV+4hYkn
u/645j+ZwaLOGWgez7w9KzW2jsvrpR6JudLIGVqzwxszBl0U1Hs8TGvJrRiPifv0/BsBQbwipMvx
lae2v+h7n4ixuwmw42cgFCBTciWlhgKzairm97yQYkSU8pZe4t0NLU0SMNgJhkpxaV/AQWIs7tvD
mNdpij1k0HKTjjEIVfeG8V65fBKiG5fiU9F0SRCjwKX107PRsqmFO7Lkc6EUQXuw+wF2akYMy6cj
mNfojg9sFterOmC+5JuvXTXhkcrt/oUQzB60GVDTCoxQtqg4t6Tx+0VK7BCSS6LL9vfxiebOaewc
uJLDMrCc8ruAxH996hy00JQiw2UXDH/Qj13q8MyFP1Y/tajqSF7hhEzF0YjqoN/8BpsvbNF52TGb
LzaD+fxAQUQTFbXvDPMXxArm+S/9epgzjiWU56KPYsJT91xgzmd8t0F0jt5/k5Ypb57WEUBAqBNH
FxIn7G9VeHZ2kVyMBaPzYazlEnVCLq/T1vWxVLfXClnmWPh3X/okZ2zBh46d/WzelxM=
`pragma protect end_protected
