// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:43:28 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
MJSFri9twRRL6zyTHVf+FJRHgl5S91RINyvyxeYqRrTqOtX+llMmpWgekSfWfvbk
keB96AGmM8mTsikF8keeGClhz26Jz/Gecb7oGga4E6IQSODLhAlLINPS3movkjgk
dV+LmpMRnYtqoEVl+qaRzjDh2mBntFf0zGiQ9xYh6MY=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 17456)
yHJHgY6TZjqB8HCUFvlAMBgQbK1v466BpCKz9JE77Ri8KgfvW6LIp74DbJmaK/7B
bllu3ozn6X6X5Tr+qWF0V3mvf8hUQpC1DTpK29xL4Hp86r89DQJlP0TGQNgG+akv
K0huaXZbItctfa6MAQPPgQXblecBkFk5B9fgPFx84evCpwbJ8nY5UTXEX9HLnlTH
nvaxmpGod+H1jEVKlWalHT8tQFqM1upGoP9Ueh4CGHubTMTZJcaaaF5lKalZp2R4
tvqaKNeEBRrw68pUTLvffTKhVGv/azSrUy4G1TF4nGJ0giQiLaGTMUoQlKJ3TP0S
R6tuzhSPTJGULRNc1xzPW3UOFoV9kRvutzyK7fhO36AB316nipDY1WFOj8lWd2/A
4AAxzW+HGxKNOEy0hAggzMerbIvLjKyunjCaHOnHNsuuRaCZ6IJN7Aq6SEQximcA
Jq8VNAVqdd/nIvaY689sykQW8T2lOgn05/P9n9fCiMPIbUDCEy2o+O5abLFYlHS0
8xKFnSP6CtpKyF6+d30CPPvQr5a3sc2A4k85cN5iM/fhZo9jdISYQmcbpftiRdua
xGfrcMMT5FAo3x+BB1q9CoecWlV82znlaJrtX+X8uzIOtxWfQ7gLJuhp96hTg+Pl
hm0mldpZsopun6NvkFCu30NN/qFtlaozyjCzhRneYA0ySPpzjLT3yv8ozXke9syU
9fZToIOecjNRWDNMQSjH8sS6TTabaUh4ia8LpuYd/z0BdtentdjMXqvHkzpu/k/E
N0dK5fwM0LHodGEHNrfudxlAymwYW6prTpTSjZav8J9RoaqphNLwEkQJfBbA5EnS
k9MsUOki+Cr5CIOHTwohoGSUwOO/ZzDn9x7q3UOcIklzB73rcrR8db2uQ6jB5bWd
fSbcNYrzy82aAZJrpPrrBNmf5PQ+TZJLqHu63lcdNZAuJr6mw4i7NnrtSL0wiXxu
Q7EAEXlVZfJNCJILYrQTGdNjdRGePaxWHBGLY6zr+7m2uc0ICoKWWlaqgVB4jHYu
UNMOuuR4kKXQqZdo8zSdQBOkkp5qAJ+ylAdZptZOcnS5IZLsn3sagyKucHYdSIed
/EbjPrbW55aImWiQoupt6JteEcsUCBtk6jVq8padtmbYsXLDLknVFhWwRIOgQwIo
YjTRVjKr50lP562VUA2sa4HwmCECWMbtIKfp2mE5PCmC+ZHeMadRlnfmK531gvRr
PUXWcBDzQ+nL4aELsUyzLw4FUL/viuovkoRnQ4WPmtAj8S08Vaxmu9awYDvMPLxp
3MKCLXDQBt3ZN4uANtVMBxOj5ho0os9yZPEGMyJfE+TSk0tHfPclFHlUohtkAe/4
46zLHp9dcnktpLpAp54Pv3WQ0cnjrIupdTsi8y76gnpBE6MzuLVTYUwhwnNlzMS9
RxwK9IX+e7QREcQDNnVExmqgIXaC2d+ICW5aR40zLBhs1TXbKnFxBLmyiP5Tyl9K
XtjG/CgdL3jhDDT/VYZpuZ4RDs+0QhG6VtV62rTQ0FoWy8WutJP0KPtKiu2e75OE
xjZdVGiw22AHMGO2ard8ImdUJx75bW+kfau920U0adK1gnaoJCb2gj31XlRWvrlM
ww9EA0V+PoeUlgdtYNC89pIAyFh+pc5XJbu0Sz3MVE/ZxDzq8VzxTEcq4/elimbl
5Z4ExezLlyC5p6ZkO/EfhMiObUVNvuryp3n4cbpgxUimiwYXhY/pMxTbCdfhVM9P
og9ZXf/ODf8rY0HdEDcAdn64KeiAo+LDHHYqmK021IXFgua+NjpidcvTkoeejfb5
n6NZHZyd2iJAUrSSARFAnhyBIuBpw44wE8RSi0dylPfqgRM+6viLgsqVak+iLJkF
NLdxl9t1s8z6nVJxvQVzkDrs/4+cvIQWvNee7IV1Rl7iAI4bW9lI/8y5tVle/iTA
qlTbAMgP5Ccp0Z66I+G11mQEkKJypTuJkQf3Cps1UXU3NYYxTp1ZYx+TgNPiJSBQ
y9+Je1afxqQ6U2Nk7DNwOR839blKwR8buK1hAAOGoGXO63qp7ti3CYc/udgxxMUw
WOq8kaKk3YT238pI8rFXrB47N6kf4tc7bAAwgBcBYbDM6J6+sKPr+ZOJ1Ybgsgfn
G7+py9MVtI64M8l5HDCgtmLPHY11Wk/Dku1FzZLkwjqdoZfxdMZ2M5szqf2OS3jX
tk0/qNpnddRlm0FVQxNew/+0JdOcLijlVh834NCXzEiH78USRpzek9o/QEDBF2OJ
DAfqlZfJYIOHEyq4qi0BDvnDRwQmUOPs/UDjK6MFof3UkcRymKTrZmFWVniyNehM
DYN0A0xngCq4JA0cshYuquQlFTZSsvC5+EneyLq8vitR9XMWwuj2V8CQvcTViSu1
Uhb9uivhEgpfVSuoN+hFr0yNJdSONg64ecjsZu4whccE58HxUu7xqgMwMxydJqNd
lcRFYnH/9mb/3xPbV/05C3smehrzmt+GqNZW29meQY8xVD0ItZW4dvCwA3Y859bc
o4Z43K2hmasOA/UzQGtNBdQvh9lK9V7jygTHM4LEHE/BoUaHrjru89gy2n30tjva
yvOb+hMJ+oc+t4YVCtvsIVtjiNI3XIhBvZqFrSXgL3t4ZmkcZ6DD+PmOC37Y2q/e
puPsVU9HzH7+iAsiDF+0P978EZDDqdai6RAGtOgt2iJJ/xz+akOA7rlAPStucpBt
SQVGXSmTwEASYq1b50N1C74ZCRTG2wHX9bQl+WB954REmOUaUaOKSpaWP5nLpYoM
TvNj+xKqd2tNwzVluG2o9SPSVhxlziQn3CTg9BWF+s1y/qkmIWd6OYdZ+wHn0zUh
g2pMU5mx6ym0uSMLWotWqrpQuckXZDfoOuC1gvWH3jIFJp9KigwptM800BJd5PIJ
yMAOjGxqHlMZQiDco3YEb+QOy1GNPoGOWIA2WOoUE3/lRKxI4NK3xSoIdaUJoTxl
OpuBsLAkMViIjE0sOAhIn76Xxpo/T4IDvk7J7psFfRFze3AzZ6d7mtTlyJYECURe
wu4hrPYHgZVm0tyULybbvsAzxPzv1angRWl73qiM5NnIdJYZQZL7LlfssxjAtyFp
YvwgfWDmae/E9sNFZ8OfYqu6sgEmERS623XKiCzp1Tp8xtAwifx/mBLN9b4U92V9
zr0DmmrgjMrkX4jzFMMkgsGPSksJ/SaeAl8CI5Cikj/8yN8KwgoGKigUYLdhK0Gw
WII6KfZVzo+CS0QX+ELKIGHbauNhnUVggjSunJEbbaIqjXk2p81quacdWVtuEVob
D/gC6x75OhTiOmDTq11KJlTooRUNpcUqWNkoaaMRbV8BIkuVxqCQtgUDrjlXsAuS
NAluJnKCuYX61iFlin92/eMd5eSp3TCbgIblD9/HxcurJErNc3VFnFIZ8tHHA350
gByRuxeJCEsBizVqlgxu3L5o01ecSVEi3zxW5FWjsgXTVPVBmjdDEN/fwwIFR6KC
3zxVEjoQxaQ7h4sFm2HMgm9PXL1W/clQOtSLx0kat7pBzjOIk6bvnwam02yWW9s+
GK1VGIQUI0eD1tt77AlnacKz6RnsgYvcQrE/ezB/rudc1r0IYmyQlX4tVG9JRqBD
rJK+A8sezs3eymNmyjf4gzPkKbm+nZiiHX9F5tRPwZkmHb8Ywm8C0bQKBRumhg7m
1nDCLt7oxPuh/nO5HoL6NCLPeOGPho6lB3QhWNYMMXgJO8aJR4gieDM5z/Tccniv
xGYrpsRpKEnPVLwTHyvJv9CVCMlg6d0tQb3wEQtM8vYmAqdr3q3O25Icn/83xutw
La3DlS2qXTeQkoB8uuVZ1P8pRWzYW/eA9Cv3M3A5WX32UysuzuEWNCacM2JY+X41
SwRO1MAnD6xdHkTEXASTZNU3RNdMGmMBpA7xVqX0d9yv9Bgohf+44mgjWfLfvPWy
peu4iSyCVdRq7XDxZuYrMdu4YXlix8CeIp4CjVTwbgV86Q+0TPCg1hvJ0qozZJ04
xv5oPh94d1kLhFQjRQu1VwVOCJlg2DdOPUYFSJV3Y/zE3VjWX76hUMIN4QE2rUIO
2qGBxbtaqYSfbsVRwpa+QXApdH0DVxXo4bm2aPXyBM5DpolxUtyauUK2pU6A3aER
9Aw+0+crPQJmMCRBI7K+RQzVN3LjvW6nilSIxm+55Xg/1yyPeB39adlX8ZFBoxDB
1kAAxafaLRvKXWURUgoYAmrHUF4LftphiV5lUir1b7TIDklcp65WohGfD19k4WKl
+9Ao/cUX76QBueGQmeDekI7BjBF6vfDubhYj9Raccse/aPUCHR7qvYdd/6EqwawM
qOrJuErmYiVF2CASnRcHf0KJCgQ6gr6fGmW/WyDqDgSdfl0CHef0syKlXusQeE7w
xFDAQrNpSjZnNlIxTGAo6VxMdLNW9fUZUMBXo51in31nqhV1jlMCKuGRQIU9VZ37
Gea43EKciBAdJrkbhKgKyKU3Sn/4ZuDtq8Bz9KZfXMlS/rHrljgk0jD6L4hUKmBE
EbOYshwDJKl9tdgiyiuNh+dauutW2axi8ORRd1xi541eld1qC17yKmiIptMIuaMj
Ys1mGzPkMppg9WwmiLsyzi1VYJFayDv2BTdmwNhmbBCYchq9EXfpeXRw3spez+ko
qRwzMZL6pFnmclFJ2g0ToyB26IkGe3EzBOF1nWBuBNFf1gqlE5vupIKP+yPrjo60
Ti+uWH7tJ/9POdchSrGX9kkARoqwqNMQsZqeHVWzrAKboiFJiPy0zqWb6KKrRGLZ
DPjU81K5c6LAVLQu9exToOYtDO7s0AhwcFGEFJH1svdfoz2QjeHEfe3CAtDxE233
qLZNaD5Jr5XEERRGZCnrDv5gd8XhekKkADPQ9IzjC69Pv8Nkg9kSJ4dlARc5ipgv
j2sGCNr4MAoRgCaIMQP3StZeb5fS+Jo8PAT2JP4KzOIWZj5EqRNrODfylSIrhDaS
f/efGMPQKZQnvG2fVC59gFWeHDxcX8/gNyMZMFX3303oMAV1E5VyZKIEhxnHv5Tl
1GwVh5N+vIl8P1POsmHHJMCPtouVl1MmHGy7OhXiMH4xgH3MuTLKmj5pJU97qX0X
bA8QJHuW3CGqWbMkpBGmeHp7XXINzz/GoAfrXE5Xw6mbu2ZW03fcgHZ7RVx5a9kI
S5mXfVuEDMnLYSdr8Qgq6UzlOAYdKPG+aFIYs8/3xRs7gZcG3MHxdqpiNuExR5LP
7JZ0L1Ts3E8gDru0v5FjtifriZA2EQEAD8M53jWPmI2HoWAzT7U8HhI07rkIAMKe
hE4jbu7C95bBVpS1t4uIV8LwaQyfvco7V4zC1/m5UTfnDM069hGDEJQtJipXMauQ
HRvYtBoPq+l1AxPrN3y55uO1iTnkvRuD7GtAVPEnGUqbzHL9/WMp6Ky9/Rl2aHH1
RSNZTw8uFPmsg2RNBQlJm8eLVjjHYzuWanLWKCOA88+qrqp8VCf3gVQKlMOA19Ff
xa3ozmoYrswlRw+9q24NZ+RHlJntdU/hDfI4IfGPXvHS5eMbsjy2mbs8L2vnFxSZ
zuilZR47Y9R9zjkKNMQmEZy6EvK9+VfzbmZ3AwH3dio2P6V5B1IKzJ2gB7MvlsZ8
OPdfTreRuCTnGJAO1SK9KoCcUUM5MwiZAP5dmVEqjfDq7KC8T210+9jNibKQCJL1
UkdURztUFoVYULCvn6Cy1QO/0xT2X1VmFF1t8ewfUTefCViMTDyLbHvs9iYNEUWt
33YqQ4UKAyvlzm7yYXPwoKYkKoU+E3u1t//S5pw/PuZ/WGIsXtWWqN3jqsscFAwy
kWwUgS0qciivaz+7T3C5TiV1d30gPJHA75HJFAlLn6Envcb4MMqQyemC1p8+Y386
KxEiek3AvAl6p3NfjACbvsV4AA09J4zlbMPdAIR7Izlb5OHXmZR+LCT1AOLHe4xo
/xt6EmLA9z1YF3qPu3wT5Eyyv/zMG32grolbxPykuSnptXfETFSJQDNg3Mo+ip3q
XiXf+7hvDs0+pNY1SdQ9VMxFnHg+jNsVsRnYPg7T6Nh5jLMOD4S8oKD/wrWgSVKb
RWsrCIvA7r0F2FP0Zwa/MCtg8X1usUd+Iyen/+cwTdUbmLhFwplHVlTkK2eB+XR4
siZXzZpt3a6QrHN5L1wQN29sWckg5UB5jAhzEBLI/e8uJ+sedm9nhkFDj1pEQpYN
DSSGCs0+ECD03osg1B3ZlyQ6t+Zq/if/nHtVQX+OjYXCN0OrDpEjGSNd5fwPAcYE
Ps7U5Jj+v8j+21C8VFvgfMeD0vkv6ZBg+b/iLmH2jnSAuIGlPccd4nPR2O6uatbZ
yCdClFCUCSX9ZDcEeYR7R8RDRKKmZ5P2F5Afc6BVrC+DhOhSXOYpESFQEjjPHap2
U0f6mLUdp/vuIsVbiEI2i3syBPeN7AoTCmVx+4BSu4wST1rUzM2fl60LZm9BvjCu
ASxOILyJ3PYN7NDQuufS5ZqZVRFHjtookkPf93Zmcw7FkDoxquo2t79HtyUsyUOt
WxyHoPY8319hYdmbp68qddutiVjXM0vOrYeLkMYuNOsLLbEXoafK2781BdZ8T28J
bfFk1deBnH2LhhHgY4swsSNyjtYm0R1qf1QSanCk+VlMEanb+/gFRen1H0iy8eXu
/r0Yzljov9JWt6Wn8hr8vbwgu1e37pmGlHUceNxJQndtVxLy9xVKhg8cnCuTzCLh
oHfot0LBTrsZzn/FrBG6zChhk7nsmD6WzFhHM+Y35fPNSO3BeTssT51hBxYAcyhO
QoqxuOz+LDx2SejIywWx/wIBeRfKM5eL/UtDIbYLqv9dmdtIIpOhqN7LKp/FIpza
eBykYXH/Lh5p4vnTvhqJQmUCF7K4uj0RhbsZem7ip3LAlclNfwNA/pYQB1+cAOSX
MLLANbYbIgTuEhmObEP5/SGgWDcL596zmib3auLoAGLOBp9RFibhkxH8GaHcFvtP
dmeKNbTJ+HMadRuwY6tcQ+J4o6G1rt8x8ndLSraghlIxLL5WWABzUCtwmNANqVne
e0VtdR+TC+UyAT8pGCGudSHg22q4O4+Zi3dOcXYyV9CZ54XxPSVbrwDa7Lm/ik1x
OjYcbevkVIugLpUYaquDdMnuTATZ5154sy5qHQ9dVXjHshuZyYqA0yNhpFjbrw9E
FSbS76gJAvI5YTXFqM0EjWfwrSlub1EmXw1XFeDFn5woGAFPl2G+q7ZyAuE8Inub
TaCqm7VRokq2q7r2MpNG1csbuof4TQ47DgWVJimIg8GzXfaIziSxi14iXRGo+qnB
MbmGy8/miaBalpiMAApi9WuQnCmsESL1OW8OOmNFkgOouMxfOvlJePKcRNGXK80d
UjeLgFSGsewsnNrJsI1Edk1Dk5H4Ntu5f5VYf9TnFNPTdh5Qb6acNyk05MKwHcUn
YXZ5WDzDt4mwWnJqBd9QhpC+3WqbvvmcMnngzJy2baDPmrBPB/4mNEF5xsITW4ly
2yhVzMAu8gSu6FsIwgY0moh0GLsulZ0dmGdv3uUOArWIOEaDhKXp9eoN6ln9YbFh
FqNLu9z7RrNjGKVkTzCTuTVufWSZLStLkMvjGgwQBbtBBchAzRWXyVHbnU9RY/Gq
iOioA2Yi7diBf1w0ZxCmocwN9tO2DKPUAqXTvRazMXzIAHjUBaEaw6DD5TuJo6Y+
YyLhV0C8rUEd8HXBdToEyJruy/nlJ+LFwUa6M5mIibV2K2GgpSC18ZSo0yrpT30T
sQVmHucCAuGRXESrnP8dHibweRLSH1J3Frd/uL0m1Gdd9Zu5vZiu8ylJ2O3W9ypb
hqvqCDN8S6GVdJp8QH6eXYeSm2ZbMGvUjpwWVnu8VsUAA1z8J9I15F4pwwZWIuBr
zPctlU/wvD5F2Ys7HNyyCgJNexTvEIHwqTuu/Sb6soiLfmXvEIqd0xT4vE50yrSW
byO+Vf89lWG8Lbz99RcjRFV0U+Mq/esnTpQzSVjrzDVlAV3o8e4SctutgvXxmWai
nu4a05QZuxVduWJykiA8Y2+2KE009RsDCl5BIkdbodA8Z6mtgi5t4J4m+M68WGyP
x9phsJNIMDr/Gl3lkzQfJpycgQrix/yq8ud6srvgeyK1W7nf4sR/Ck94w28Tc3cs
cVzo80FQ7ZEZWa1qiFEGw3BmSFrrpggWStoxXQSNMoVxK0rZR9mjYPaQVDqDH0Bb
u/FYEjhqaOHJQzQ1RFw8rQR8bxtJGQskcl2f0+9Q4+QHxiOjZrbEx1Nk1wt+hl6B
G2EPjf9TVRtqkMrLp9uJhKazpmUtD/GyCq8STre/VkXEj9bVTOA0ZAtd7sfabvod
UQUE2FkYRTTBSBztD97iATFSlbYnx3sbCkupdcLQUwtlTqM5v1UqxtL2GJddzRXA
JfX5BhaZd/qFi4/SVLZrs/RlTgS9wDQs/RtJGpIFakoeRRIGhRcn0loy2RMvwTFk
8AIWxmfXa3Vj3S6gyLOWg7650ExyN5CM9VsAm8Jqlk/Gd2ARYVLYVqkTQr4LWcT/
xyUFCSuF/1oTDg6iZ2HOXat9s5NXqWdeCcpzfO24L8Qq4S0qWpjxibzpRS0hkD0x
Ly0JIZyk+j1rfFcsJPFHe9unv1Uu1DS3qpBVXTaA7u496kpvbh2mTh3ALcQ6+VdN
zQF7M+jA7b2Stj399gvKcPK4RwVF756Le/uZVAftqUMmomI6PkF+KzhuOObSGeJw
Pc5PBg+II3Z5CSHk/lf7JxmlRaN1Fh3vCklPTtG8sJpRk/jCCJR+yd9Q2EHzmVKY
rK3C1YqpTjjzzsNABoj/yowcuMfm8Rkcejlqqc1Cf8wINm/l4kKTkUgXUGhq/tp+
wWglrGvxxvkhpWWDwYnKFvFd+Nml8Pm5ov6UoTLimC/0oj88SZRLQI/GE4/jiVNM
LWZw5Sp2JHqfu4IWVqUBeckE60Mbv0UIb1Es5Fddi+QC+aOglzSqKui9dekHv4qW
iT+9wCiUH16jvi6nfOKL8wBqhsb7fgP9ORwbgxBayCEumxmv+hGVC05r9YZCuItm
EOFhq/TPCzlZcKu1rT84ugXY6fITTKKDf3k/wW5MkQCm0p1WHovd5ugVbSVMDwp0
sHuJfCHcubxOZhz7wRxUvOH+ukb2WOZ0vczk99isG8rI3k6/hVTzAMGFK71iXE+i
xaoPn8+d3SI4zt/1miVEfOFHpuiI6QluBVRV4jF3qhAT36c8HyuPrR4N871uuvLf
nyqmJhWdQrcCdh6VQMSisg1ArKQsMK2Rd6HRSy1nelYl+UwzHGXhBor45evwuWKJ
mp47o4VXNHktD3X4l0YuH+ZIywUd4pDwzrRvfokEFGMqAVbmFm0utkKa9ySu6xRB
CJRflD/5ZgqE/VUPwoZotcS/4wEBVGVr62XLxeJEZaMmOUPrL8vCGbghznIPjzzf
y37rjMx31K3BwaxeOx7gFDltiIqU+PA1p2mSEknh/3X6cKuj0oph5ivRO1T6MGvS
79dLd6iXvW2jRxgnFqpRk1d/JRmRzZhCKjqfa8ivYRk7uhiCaWXlIQdM9SYKhXTt
jc5IihQAeWF7WdIthLgcF7lL8k1bl1mcQ5TBLWQm4UMigMIquNPX+vRBhYfQ+lS+
O4JiWwlB6pD6natIFnbg/9YL1jWrh2D/fy7T82//3RhnfeVSuIzjz7guW0Hg42uE
jGWEBqzF4rd5Yz/ZI78rPJNDstBtzlDqZ4iBVjH4jl9QwSvp47QE/uXI7xpgYyVZ
zROy+8vuqc59mhmhxSGnflXAjxl7sQaKvHaWvx6f+k9BgFKmNXfxl4vxrjqGeTcd
XEVnSgt7jCTtdwo1OqwJuQuy+5jv23/tXGlY5Lt5/gkjXGbfp608LKaAbgLihXEL
cGKcL2Ax21zTOobK8JhAVYYd0vt7mX0TzVnLxWQfglb8usf+nOw/RxtWsf/dKrga
0ECnAmq/NcILRn7PRpT8ZQibSCKzOWkrU8bqHRqA8CfgWPUkuvCJwb5aWwJPE2jT
0gMCT4/RBH5+a6OcrfqySbBJJ+s4PbE47XIXKfW7i9i2wmsC1gPetaXpoLzIXXnj
V5J4UagwUd+aWu/ZbUgP12qfLGxfozkTb1N+v9XUJ+bEt8p9lL7aCWXMFlTsJZ1C
pM1IwbmA0yO0DQteT0SV0j28Sx/LpXZHHC52cGnobtw/4oDHP76AdVlgv3erCi4J
jeM+EAdH3ulVEcB5dAmkau9fWEPLVNmk9PQRTzhdHUOdqQvBvEs8egc/LBRCs7BM
aG++/GE9qKg9m4+Kebv63SFCafdh5h50Y38bWGDdWHNxnHnMfc3bOsHczKsWraN4
xEEIr5lI6IYGx7IK5ByzuBgF99xRYjL+RYC5sG69/+CzswSNoaVnS9qTMECkNTsR
AmsmFMr1A4cDRvAR/FpEy4dhpJgQJcq/1/kKlgrP3HKBQ7YJIRyrrS5KhhaemiJs
BFOY3yy0vAMeUUHGmQ+g/VXAD57L+62pHRK+/gCqolgKkuz2uO0ZgZ5fdCE+JWvt
kT0aAEymg5lRJfxr2XZ3hLYvyERRJPW5JjP45Fbe4s9EVGOBha3Kno21R0dXH6dF
A5Fs4fr12hKpugy8Y0JzUn6ykQIvUOTrSndefGJ3P7tztnv6XFlL2w1/skb3/wpJ
9quvBNkImI+9GjHJM/JghrNz/JY1FjttSfl3kBS9EJsNJ9JTw1DYhaSKTMampz8Y
VU2LQj+xyZ2cvq0UsaOITUgjJPLjMW262lUNRBq6KPYz1ZF+UPO9gDlFCcIHn/FR
smHg9lkadmdJyTRzAyjGMLC9QnZCLzTStRFQqoCuY/zwfsPj1GCYFsKnMdsTyE1Q
7G+IfCbBUwyuyz3c2fNRkAlD+Gy9x4bLhEUSBMr0DiZzyKIVSQ4PpZue663qTOcD
cDLs+e7rLHSbeKeva+u6h/dfev7WQDOSBRdWs3IwueJo6MdBscp4zCTYhL04C/oc
F5lsHccY0atOAe7V7au7C49SywYHIJmS8RgvaswVy1NhizVTJcFdm2v6TkhBnfea
wb/Wlo/RKakUcA4k+55f8X4kWMThyyoZJbOsEzonIH1RQTEqDtNrPiIaZTcHCk7f
wH1CuzgX/kBoclWDNtg8nJn/d9Xl1NxVWGnrT5VMJMTEP9Bj41DxpV83y8Ga/a56
tSBGkfLpVKDnnsYcjIbJ4UDjX//ppLDVd1vn0HGZpr5HUkzh0h3ksTCSWgIM34bR
FaNROPtM8n/1FBd+za79OjJmGbqaeF4ruwc+KMn7DUBCTKMFMJYA4ac2OAShcLgg
08yBdFnpdHfsHJd+hGudBZKFv9hOckLfmaPf0YeTjpAlFHNkH1Rym5G3WtdM9TXS
ZYVgXDbgn+uyqB4KWo3sQRZfOtbsO6tYaul5WBphFLFl3GlrtiCpmxQdF+tIwQJJ
xKuTTjOPNbe5+8TkuZwC/ObT5aMVK0SYNXDRhfdbH2BgI+PvEvLKOL5flfp90DLZ
Yil4CZQiJXxrS4Czo6HhEvYus8XrNhs2v+nY9Cibr+LhAMIFbGl84EWP1Zt7y3eo
OEStzQkH0qwlCzJPB+OYAwB8F96cI60Vi6UabTSjj62fwT/rvq4MeTw8cWQaNQF4
ZgAS9T7LD38WbL3PhtFHmZfoTBqwNXr1mqNfzGbg0nDCa35Qgz5ESbLagb5W05UT
kZ0KuxvlD+pZfuifQDIZkl2S3bGCYtKrRts4Ri0BMAT5hAfpibxq0oEm9s6+wvRD
l1MBnun8v/OeSxmqGzDQOeW9UNVtPOF9rMh3RBYGOJb3inIhfDXz/PQ0LQT1UB5J
/WvqfhNohI/Be6a0QdML/zKH0CL0s210VSApmidCE9GxhHjx5clJyZo5WGx2O29d
veFuAXIM6fTVU1GAU2e7ZAieyZMyOQR3wOHqdQSVNKdb6NvTGrXmsDu0h9eFyr4f
ipwrXXRwXnY4pm9/anmXq01ysqdNHiAc2hknRSXOFadRLydqs3VqJrXNHSS7ZHTF
ppM3CmcGFbYrFk/8/uT9cX9xAxvYM7p43Q1m5Mi4ejMDrr7Ru1fBeO4OEDfboHcY
SjrZfqZf/6jrJgBtJ/1KXGguyM/7XQYz2ph1XOmFK35FU5Ed14pn6/NxddxzyvAo
UwDjQAL6JhGuGQ8mKIzFi6+nkMIWflB46MF8bIntqcwjD5MOskIrGB2y0Kob4SM0
CODsoTfeJQQ30V5sQ3bYO/IPQTo5Rxig/ayOOpHOyVwZa8lqd3z/Wo0l48jwJFk+
aakP9ascIWKCImQe0td1x3yqzi1dXedqVST+4toniZ6D/23vu4RO0Pjxw4zjYgxw
YFrfo/4zQdxqnBuQQsZlxZUvr3qqRELb168yBs68eGLCwaQVWfnwEBp+udkSYfV8
LZF5+gW3cosp/E69O5Qeah8wPVDGJkiTYO6Fd5J8bSslEpH9GAl20rgwIcNLswBW
whAuqXy2IF+dE5U67inGnjaX66TvJX8c5pUMO4Hij9nXYL5yYNAj1vQ8zpVaMWli
BZHdUWCTdb68h8UTs1S3NbRUXeNSF8oIiFD6EsOMip9MiaJO1Nzo1Ni1kC1jwvFA
YCdqxgF/m08FuaTk7WZISuRo6X5olPESBeSU7iwdHO8hQPcCr24tvJlFMehwCSyk
tVl6t96zVzbJSrkWhsuC9+uZVtxTLBXKWorzoXBOT436CTK+zfgpKPjOTEg56NDV
gUkghZ9hohUqop+0UO6AM5iNYSezFBxf6FmZOGe5N6OhqKAtHl6ZCcCLfeRodcDx
J6nRm4TEO45CXR3YIWZdQZg70de6NkpZBs4WmNHUzaPApxLgknv9FGjqek88IjH2
HKxHfOcDC3dTbhA6gEiS05rAfQaYhJtGHbsmhVg/szNZWaKnmOieRpQ1HjWqX+dK
wMZ9SrbOg23+t7IeoLRniy2j2RIdYU76HbtJI/ZFkRWY6g7UW9LXoHVzdHguYcJH
ggW1nluBNNATerdRBZayY3ztcLZMHNHDzn1z2tn1ZHgUzHpILVhRU830evT/aX4C
lWVcIa9qdG4HqSi/kZw6nCSXX9UgIINo5FbGr90LztlAwWyucRTHXyMHe3+fU/H6
0eqxGrJpKF0ifSLtKgIdPlEeV6SJKsYUjhcSMWGR65ToPYBqzijDTRaRGCNH1mMh
9qOhOYFP4lSjfI4JSUGCWD+lPXygW9WdDouwj/IN1NaemTPxOefbCh46u6nWQKl4
8ir0O704VhQU953LGcvIuKUiHp3C6T/LMlGDSdqSLK2dpUDFnmCuROX9Bt5LUqWl
8yy1ntjoCS3k5OZTPCGzeGYZrGxIwg32/OfsBt3sIeEFzYQHRsKqciuLZ8J5imoj
/NCkisLFyL65gOO0uuQJwpgfe8hDUwlqxBO3RVuvPQJuDwkVEW/RDrkibyBykMTt
u/9P6PtC9tM6aBFU7h4cgASJLhTaBmHVmbmrpFAURW+LOBQN1Iwfsq9TbYeD757D
ekn49+/FzDCuys+qwz2SClUcU45OnUAjXDocAi9veCz+UozGTOdijNMTKBD3dby5
r1oCTXkbV5osvMCfn7NkNxzPZQbzpLvGO2j4xB4x2EsRBz0SxJVgcbcKglSJgZB3
1Fwu4Saa+MgZaVG/7NDxnz0u0EX79rdo3LoqPRPn7z2gwa76ewipNZ+gbBciIsFB
Acva52uin/kkowwDAC8W5GbVIn0aKLiOWgqPE2bNLWHwfsbduBTCBqeL8rWxc7n3
Kk0iCokyR8wSZPWuG+Nqqp28mUCgfMCGMjCkO+JqK2jgvjZoJmjY1QohLmBuhWcr
sANk4bTxpz3JqZwqppGtZodIUue6y0/C+ZZgPfceHp8am1PlumN/T4XpioRDHtMq
MR6sKDoeEHAPXbrR+8NNV87YYRySlhmtxak8uHd9RfVq76Is++RKnTWqKKQpE4Zd
jDjCH48pE3+/7qZmVbssqgIk6fw2g0N/nfoiDGbx8ZdXTLcSp8E+T1O9ndhXnKP2
dIe4vUlZ/uN04OHgb3Vi1tr++dS5V7/ZDIaH4MEMYHvOCZEzEqH5QwYxAtoHkW9z
imJ69uVL+VKoEWmmuDr5xMfDRdExSZs6lUVsVppP8jl7ysDZsH07arpnlriHIKQi
ko5CD1HE46HRmMqXmWx9lfAsiI8MZaS+w25wYfM0vDgQdmLQhSHQllWzhd9sbQtA
Wi6qiZj+cl+cfKHgtAdqJWTVy5tEMAwLq9AV9l6cO1uP0Bdp+hkfuiSb+V/qpTPw
7ceM37tlcbYyJWAdwpnjsVoH78kcFeNPszkJSH10oftXTy8iSgTD6qdhiRGNqf4D
a5BmQFnZ0adpordWfKhcgsmN4v+W95gDPCbIJmq/cbK7aht2OwbVNN4xBDvOKGZM
FUXoLZ2YXjj28GPXzZkLBalIRNYnDwz2/DPfsICpQGfeWvSBxgC3uQSf0mSxw0NX
zJH6sk8/RD8Deq+sPkLgKe+8ydKBwdeFr5OEu6bw/1xWpWE4U7wYmgCquYMcYnt/
bNpaQgdSDWqE+/Sjx85Re8dd1yQxxexuBWUHgm18fJ0hWZgxyC3AomsgZ46RAWHn
IV8FGHRXMT8FWLQ3acLVzHzusahQBTLiRO2DYioUughyzj+J94hrZWWESOvLRtzg
0tFuZPXPc705Y3J43i0ppkZC4nhbJtuycX7teZN4+a/7lzqmBxLW1Ri4CFmWWbgC
L7yOQc61sItHF/B8QsDs08lX/mJXtCgxV6do2OebosRyRQrCzSZja1pxSLMrpgDk
BncF/Tl7NcagN/fl83AXfHX1uG0hBAoV3m7Fc/DAFXU1GFUV/12ud2XNWLlXgu4s
+YG74sbwUxJJtGgKicLDk6RbB2GARymsJ3g4vyHFioc6WsamzvjTg7ghjki1EfZm
qH96C3WOnMeWoeHbZm13C/DQyXJePlBx+381kC9GtpC57+U3HeohgHuOEp0yrSPq
IjuCozPy0Iur4SVXvJsHp/1CXf/I5YdTy97HXK4yNAUKdApE9YcxmygfozV+IbFL
LWX8foQobKyluqkExCeuy2U0Kln/FskUcLhHT7VLuoBhasOHCEuG/+ztE4KJU0iT
6vOPpW/nP8hbHFsNGEdim33abGJ6baSpgIttBLuxXHGvY1KQOI1BDB+B/uAD2Yvv
AX1SMUcwQgbd8puMT1Dwf7LBnnOE7YpfZ7ZRwuriSyDxUVf14lamtfNN6DTC+DF6
L8gXulgAfF5wYsMdOmEJBwV373bAqJXycMnDR1RRQXOPL2vw6D/wwZe7CXcWnqT6
EHKquTzbxRTGfJBlX2+kseqE5Z1VnR+9t5cHl5m8ftNNIG8ylnsbJDGaO7NTdKnd
ASZtp8Dw0sFSb08htPZoA7qvSx5mIsmOL/mLJA5DxpiXSGKquyvFsUAbMuLPaW+V
LFjAgvl3qfvGPP0vxlCmAkS0F0R4/LLnGEnUnh8KT5FnL6HCuWznN501p5FHXAyR
mAmZpj6/0dnp1R4rwhnXX1/fOT7zr/+IgftGRzjq5TSyhtZT2CU2RH8Gv6vo1Drr
Et+mBPBLp4aMtFwFE52dRslu0wYUfhBOT72zCKUAT/yCfxCQjkPG+croCgndpFeT
JEr9tAVQx0zCWTwHc3U8o3YweF813hdzKnlxJJXf+XWSqYIYXXRUEXzfzax+gAtg
V+1vAzZ/Fe3YldP3K+SifdhZrIaJYnRnMp6Hu/AWY49SOXrRfBYGf3W2AVBkdYyW
EX8rHQOW7KDxUSlNRsy1/t1nQj5a89gK8ece8byv1Iffp27OFm51W2p2Z7HOPlO+
CtdwSUm4rvciAEkfx6m1MVtW7SVUSECVBs994NJO/78wOrteyNDdThq/XZ7J5I0Q
IWon8GCNQJBZNYNjvEbfoY+IpICTHfLIdEdRVRW9NGiqvPi3vrVqJvKAX5xBSiIb
89En1LI+APvyOMYDkdDHKXFaeCppQ33hCj6oRIocYSu82wZhfnirRgkBieB2Voop
/IS6qihw9XrcoiZn2R+685MRORZf0T5KdKsH/WwIznAIu0ypiZWOjzYrrkqbnIim
B0FpFfs80YewTt7D3LfcmM/4gse2QQ6kZPDieX+ctAHYun/58MsSPodamgl99sVL
/JxuuAIjLlwaz/WU3cwQa8mAdw8Ebyv7ciZBYNh+mAAq4pFvatUg7tBu5n3rmDDb
x6bgU7HMBzQFFJhexr85r+cCgOX4nzZ7DMj0zCZZyLZnHOxoYCCHLpYJEd+02EkH
vvvfMZQPvgp3Df51XM3YdnD0f97g0zPL8zn5A1d4+JpoMC4XOajHuk7YNacBTXwE
gfJB5M8npIESFtM9hxCqbCadYlhS44M4pTSRtLPH3yD9RptauGBT71eynF4NRao+
fsxg5AG7CMhIev9uaMBiAObOrZYKZ8ZoPI4TGrtYSa8RHtiG/aqkaOXgy8DwH1iJ
RI7URbQ9iMrV71mhnNJKs14wpodVhcGU1mcPziIckLtVSXnP1YnLF1E/xpymHzl7
47oEKqHBAvpeVs3nW3jicVsi6P0FN0xauESM1N4Tq7TmFiukB3w48LVyja2iaJrO
w2oNPKjvVuYwV81wcTGq6IVLUH1mvbrtghUbmBkqJ04rP8Zdlwy1Dmrwvm9tFkZp
Owk2OBqYB8CJudgrMdrpWZexPpQzGEl1Smgn+v0W/psQBS+tF07I+tL4fnujEOUH
C/Wii/InBS1DLln4QMjYoL12H+IV21BGkkKfrYiggKM9fcIYvv82DFw6u7XTk0uz
8wpD/83eKOj50XMEpIYtHjoPEyJg+oHP/1OCVEv699gwSciZOPfJVmmnEmuneXBh
X5HI8p98Ie9kNVAs4/W/1MZdLITEVnSxoDM3gWpHOy6AZVCf42oPLV4v0NBXl1LC
TlF45w9mCxlnzdKCQr+baEA5LpHOzrCsLr7BhnYbPss/fMJsgelDC2h3xIoXlxul
EGPkuAbXep4eq4qGC876tRTj1A5xfU5a/uttGfrvReuaed20H0Er2iigWF1tmncQ
GIM27gJi71Lm16mgbUBfjCgKPvZYucoZ3tWv94FRkbZGANwp2lbGN5H3RiOXwyjs
YGf5cthWGj6yGaytzfxnSpyWgWbtiJRv9Lj4+dUvJ22MaFa0i9dzPwfMiAXrwTi8
EaCmu28HrJbtAdhQwy9f2E7wfu7FYojsFLnpYMBWFOY6ocggbjn5yqwqbI8/6GLi
Bs3jAHUJO2dA/YORE4NdhUJzIHzF7OXL7A/Sk8UXkJLBliHoh2xCn5E3pG2OEeMn
w2QjDfG9e5kDKvNzp4qtyvPdgvXOjgIZQ/G2k4C0VGV3Mq7HTr6YnPtkGrT0l06y
grOklnhjX++N1tRJS9z3ntCKSJJBHhcXYutRW6cV52icKbhmA+3fjDhYlPKXZiOr
uOhuLhBo8/tNtgQASCEKS8eU4RmfTW/gcyB3cpz1h8yQ05DaIysSHliJRsuSjrQN
wtNx+sygd3SOTm0nX6u/RSNH5A48cMxC9ZoMEkAvlzOXIzZ5+STwAwm1wUIKR7CU
W2uSeKK2zB78/ZsZLHNZtdXfvKuvWXliV7WB6auz9K3glYu1+7eNm+Ee1m8+8G1U
TLc3OfSPf7lufL/iqwzudbkLY6wPEFTp+59whxwdSi6IeBfrfj/pccD0Os5ScWC1
8PIto54bQaVrP8qrYuON3nbDPwovaZOm0qSa51gVVvBnTH+FbKwRntYCflOf6WZf
mPBM8AfDL3PTfq9Q9M7ovls9K7N/ckL//Wjhlwxt3JbpIv6ZeRCroUYLcpa2/I9O
qN7LbTBmZ6SG0XPNZjbQ9way6Uyoq+ycbBvXx27l6VnxmZaBbxAaJYJhNw5ZgKsR
2e8GLvUhEvcBzdAC4Oqimdy8Tiv4bc47t/CkQ5adt0gDNTsMjI/gXVWbt+95ZHNU
WffyosDYnJ2/zDO3HpVrsbjb4gd72Ufc8c1kZFt+tADJt6rp4mn+zJpHIdC3jhz9
HjU657vaCwGCazY/12C9ZB1piL2TC6k8+Y0LU7SMsmiFzFQl/Y7aI9JggXwwxhBr
MYVnffWUpuDskE7WS2/Lo6Vx53l+0Df1BGEA5/WWd20v186gOtyyHYHDuz1cTgaI
nogBDX7fehzGTEvTXn2L8/XspasTHfGFTXCsoxWJDXl4wi346LLmx5iVoD4TokMZ
uO+bAoRQkGqDpWpQLIT+gvLqsIYWM8iEKSs4bLCd+3OTQeipqTRANbH92IF8RkPJ
J4AzqFzBDe4jYLs3mrK9e1py9Bt2RG2nwnfR700BddTqq9oUD7NDiUHd7M1B8oyL
KW3COX5CeFTO4fDTFQNufHIw1ZU6vjIMMLXDWKg0eDdLyF4onWyX3PxkvgAGmW5O
ZeDTQlX6HhpE1W23n15iGKpTLyuSlU65I7Z5Lp43gGPeV69Ne4nQ669HQka4n0lR
DPhzY84iGzseZLxWfPK+BiP4OF1NqcQpn7/+BkRkIkLokpSADEj35D9x9y8nORS7
U8fs8wOPOcatWOl/pbjOn/CbeeeL8Q3xCb9u00oFcIPOnl7L62jCpockLTaeQu/M
iz5uQjJ9LLHKGDGvTISAMgYUPpoU0UcncNZZcIOz6lQMjCDPNV+Th8YcnDki0ezJ
VOxqlYB9dazs4MSMr7bRAMzJZFw4hPcz4kfGSgtgvU7fCQL46y0LRjmu0yYqIpOF
FfOZr/kgB/hpDx3ksIFSMxri4NJuItv/FFxvxKvxZQOWo/RVS6Q0RDMHzB+vHWvX
W4HlsLRsWurmEvPvnbFHdSxi8B+SqugvpDRo5HNeEtnIxsFg0+L+uFgR0wnnWcus
POGsFsr4GmLucWXWsGpdXu7b0zkqsNY00u3TE5E0F6KjsiPDfW7PueVQ8rX5vkav
eQHUSIyNNNluira7PF9gtRZJ7jImvN3+uDYFb798AkZRX41ZFCOdFbj7omLcAfM5
u6MbVnzWJlpfLJkgemBOpo8lXxnkGV+qLFPTpmbTuOg7PKFG9JieIYIsHv9H4jIT
ueFpBdcT6k+mHF39irX/EzZfZNF74WOKaPXJQcKmQ3kkpdYgcI57tmyAJu2058ts
a7yFEkziuEkYcUOopFIW5v2ALQ0uWx/6LqJ3+G6cWPGUCKTzp+1o9sbtqaJFrnIi
KMBNlK7u2u6fKJz2/RLTyQxnqGPTh7wSlN6LXxCDND6mZyBsXLKhpy8FVdR15gtW
Dp+KWu9EepBf+4laXJz23LMz8fePfBfTwoOmnYlfwUMbF23IUQ0i2jL6skTzL+GP
GxYIgDOB2UWQROdHVdtIb44M+56DJ0Z8Z3of+tP5yxvPhQC9Ahjm7H6LKQl54k58
LUfXT70znldPNypOxlXH/is7fu8r+BaTmeTY1t7KerkVoRynPrkZ/p5S2/6yPaMV
WXrrcP7rWQo34KxG+jKxZxuzXFCEyVqrd1C1uO8eDARaHyWYVBDLvSpj2+vRWrJm
DVKXvYYOowJZyetTeu9GgLXNKuPzmbsDw4Ie5GaXDp/9jkisvkY3d7Z7e168lHmt
480YzV4tz/M+nNNiHjZFBDRky5+Dzb5UgUrqnaI6gEH4aEjJFDSpzCtjOhp/mltS
nplcho4qjnmpY535ntjbYnoRFEfUqlqLcGM1Y76unhZZCa7ZecaWWIoVHxRj5ns1
rKtq4/OPp0Ac033LIGTEbpdlUs7sIs2FG0Xelv0GXA8CMlokijEfmAFAandJYfbi
Ua7Aor7isvauFxqq2ae56U8/93TxFfpzWl+ZTt6J02/xwRk+25ML3/JIm3Xz/N9g
tcGskoTcxRXSQUZQnIOXfspJCn+EeaslYMxGM4GUiJkmlFm/YDAsnlCZNpMY9rMK
qDjudsGczLVaS0nnyTyW0+cNo/35PQtjDw5Ewouftx1oERmjCex6shQXcaZLeDEC
wQpqWZptwX+2XGAiFtdGGxwPCFQTqIJ7p0qSVAOscUpbsrRK+JPkhkwz1VQLTo2C
O+09gLtiLgzs88kSONf+5dyq0TAULtaDsxSIoYPDk+husRJhl658qIlGAZyOWoBO
cVBo0cEmCwXERq7cPtZinfhTMYhz38yFubIjDIHS6sJ6++QL/IBM5ouqZbNevktf
tm3giGly5L9p9T0z0hnv3kGMckaK8qKik9HvgJ7yYYngSV3s7sXKlDp42kYGf+CX
8b2eHgV6Zl/QJ5/NjoUny6UuOuhS09L+MH6yuS/za1GWOAygR7iuIFUD2PRSzHU3
WsC0+XiR/OZams1BoTEglFldDF/6LX6qcG1YJsfsRwxKkiiz6vzW9wXkfZmnHmsP
W2OUa43hUEKM8gzMGlJQhwZKqCKF0Vyr6szzJKulB5vTjBqq+buBqqsRcKotDwJS
EH1saO2R+wxPegg67ShQ1K2BEjm6W/eC+nxpYkkV0ROpB42Jihl6+/ltw95jIwM/
tS7Tf6YaTxEBQD1y+UnUbpLs4c1Amy77qeuxen5mHl7dQeUkyebtjHOgdHwvdlov
P2+GuWNhiu8d6ygt8qNZYFGVmMPLtRI6tvn3FxbZs9fkweOD02NRoFhNvhTL6TTM
EACzVthDqQKc8Pf6s3nAtM2WY9KhmWdW6Ckr1p7yOZXJDALlsnrlumXyAY9LPAeZ
OCwF0RclTAyZ3I6rFLB8d5AhRLuET9HlgqzYEv+Kv0KCqJrt1qUAbwmu9WqI6Uui
awv0LHPLIhrSbtCQpd2WUztlk+BiPCmuK3glJHyViJ3slozegpclqNZAVALdkjj0
2F06THKiQTWy6Xdc9GgwLja89s0PJ1zFrg+Bd1S7UEiSOq6wHeNNmFL0lwjhczo1
dliZpT2Reis6NssjttdXkThq5ILsLyde88zBp50X2qQFB6hcKIwHoxaYus3QJdnF
Lngf7NKoBUS3D3K+vOlhKSOQ74KrmLzBsnDpHV/kbPfci0mw6bhapSuvGhQrInYH
Cz5SxnfNj0vSsrBdq6rYCKmdd56JKXPIyr/InpbzSp7AwPDTWvfxP7QErbPQT/8s
a5IrezHUWmmKjxs7+FCcNOME05mljrwwmjpZMwcm5dzx/VADYw4TOUOjpTfrlfqU
cnuEJkyoMk3lWYR1Hs3F92bwk2FjI3G0tAWNkDUtNFOjU3/DLwixTun2mj5jBvXV
+4LQMc2aE8sJaHjwsxxn/v9vOu0na7j7NxQgjwDVann3m4HXBGTbPKDJ7dXZ1wLM
EKrg1mn2V+bHMlCDy511DUJtZwL6yDX1pQ3qcbk+dFkb0fKbd1dx2glbIMQHpLIi
IgxTZA6K2twGrONT75N0hZPIS0ZSnIZpU6r6U4mbtK270i2W4Xi9sJ4pbJaHC93C
gmVUIAl9gp8n9/wiNrc6hg+ZFGx4bVzCPCwCRDz6mLPSHpFROTPpv+aqOnHDRc5Q
BTxL83ZKbnNTXExZjASOHsNpsRQP7K4wqLmnP5jTBjpFuiVXUTla37Wm1cjUuN2E
3jPnRuNK++8NEmDi5WPXw3iRhdUn+TbJ7Kw6cXHi6GZscHvx1THHMNdKSebEcRmY
0beMdY3IwPtIvdvHWOjfpjJ7QBa1zmLQAYYt4gBcYx5ngMjUE6g2cqILY70Guit4
G8piRS2uU5CJvhygTWs62dS9uTGYO3Nm2ZNREaHlaglTE76T2ytgb5jrOIYnZQI2
QjuoHXVH7ZhHchHU7VnASOb4SH9wBZdTRvChnvXyNNdDdqlP8fwG43oRCTkMHg1s
oiDyDptN3PLJn1zwxXvTuuQijKmHKBngOR652mRg6CTzgNsSXBZwkcElOKj88LyP
RgycvDH1cfbODO40nTLQUWfsupFr9MVzIxniSHFVO7f0FCWYhfvDgJ/lPfm8NGBI
u3IvqBsaC6zJyyuCnSvHVCDfyeMMHXIhnVhkA6cjpfVuyj00v+zZ5ZMrLUtTRs/J
8wXG64XF1yBoFvATACCMAiKWflfbxTiGqiQqJjnYS0BB3DPlNxS4eD+A1mULpKiR
z+4cGYKdEJ7SqYwghqnzBq5B2OOFRgtNwP2mMGqzq+ZEHcuBKIQk3uWpRtVcOt+c
Kd+QaUYzWZ2Vkjg63pty9AEOzuHwklWPzW/l2H5XABvvVzv+8kaqeRxNzmJ4Ivbe
2SpCl7wHrsbgyujNE4YZHz1nE1wlCJ+Awz+mg6NtIOWSvhN+9YyeEHxJumT58Tas
F/PGpybwtcmHgx4SAUVIovkLrjKIGVT869HrnnISZBosCXcOO+otIZ/jgx36urff
wxxgmP4SjIfBv6YX0zxMv6y8sMXF8sGJ/rR5kIeGVXvkjtjBzelG5KIvIGrEaZMd
TyDtElTIJhQcBr8YHEOBVEW8nbnmfqL+ng9JmgsNQ1QmZCN9WeK9T9X80HomCjaf
qozlW24QE8Nso/M9OzQbDKrsyihwhoQoKwW9dA/WQQcdq4qnUQY2gEJvcFMLa93r
ciqt48UTLo826p2h2k/70+h4EgQD+rh9KsBPoMTpa4VPxEzqQo0zvcGFGLZSYgDv
oAYnnjUqYiweVR2rAIumoGpRInzujRnVP1DrD2I9TaC9H6f71H3KniN4HakL9jzq
nlJhsruhHEsdn9UMKppjX2X5wDIGPf+G+xCGvWQ/rwjZAPCtpTk18OdPSOjPg8yG
phNf2wAKe1wtK/zkI17Cvv6uYWw7LLFhsaQ3C4MTFrRJRYS4L+UURMF7r1w08eoj
lUquLt83LU/8qboNRFBkA6JIYkS5ahne31xr1adVk/kajv7FGicTP+h8GVudg9gV
iiUWVlzO18wOMbVUiof3meuZtOUaln7Q/eL8H9v+chpyoy/Nz9S4GhjzW6ovQF7A
MwAzhve+fCqPqSEh5zXfMR60uHAldOOC7VB4Po29yxsmxC0icM+J4QWhOBEMg8jz
7Z8BmRN6PH4U5E8L4aDb6kh5XwxuT0OBrtOzFfUeDZDCyAib2lFjLT0fyT7YCIFQ
NpN9vvaU+fhHDruTlgV/LKDUSO9ahrDbHMD2DgX3XVcBf6Mt7/IKlNDi3+Co+9Fy
3hOijEHJGkDZ4sEyzbQPLkM9sg33j3eocKHOSCCSp0DKR2DMGVx65L9NZQWH69Mk
w/40vGkfFq4wsskHPoiEATJg++vOqYeAVJHoJmyRdVcLDN44RyBJ0fHzmrsBucGL
rg0cLUADe9Mk9OCBGBKoGNW+E7Alu5YS6BoOGQTv+2W2hPqQ7ronUAKZQ05q3K4M
BkD56eT20Ws33o8lLpFGhbuJq0eNyRQ1m3k1Rvr57okdSYzxPzw6VgOLmQu3Dl3Y
s2E+PJpJKvyJAWPi/SvMCHPVkqLLKTsMLg8tFNEMUXjbbrIwRrAi06pS6aRhYzl8
kq4rSdsYnb32/GGPaxaporn9ndZjnY7GybXE8VNqCydhSls0po4cG0Bj7dqxOEhN
GqBswo56RWYI4nW7Oqe2sJOqLrE62engZhGyf48huuw=
`pragma protect end_protected
