// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:21:34 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
HaSWlsr4AJ3MOyg3Fn+AuO7NZa1VFiG0sZaA5JId+NIwdPR1l0+BX6qDqtRoHmHi
ddKpOXd1qUOS6thM7BfBPD7aPCA5rl7CsFe18R0yZx8HBjn/+NdZMdVtfYpTzOIN
z4O9DauzGZZpTDFR3dSzhl28MnURdzqb2OiOcELQBrI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 7424)
7uveJroguDRGQTTYPntLwFRYy7FO6vHWIadq7Ajpbtl/Ud0QeK0xr0I1CXWHT2iq
zxZHBokGJJ/n8oMNOrSoX0doUhhMNP9fL+7zy5BsnUkGJWF/5N0zds+O94c1E6pR
aT91LhkAiujs3HrWp+is8Y/Eov0aG1xP59SyfxQCh3ZppF6CAbV+XaMSrleGNIyh
xJG475ZScHSNxUIOUT3GMIXfUOwrGes8Ofzrj4hOdEy8Z25McoEArY4WBIbshF0Z
znenOdcmAJwB+8VD1DDMBddmrB5dhcddXlLcJYsz9rJ+DiuArvoJRMmX4sng6rvm
dByY88ZO9oCJHO+3bfHD9swiN3fAYyFvshIQnCZ3ELKMvGOpzbgAZokxCDR/kxX8
Z0096Oqd3TvEOiXlKWR1o2fgWCbUWguLBCjXQxnQFNdc4LKleK2ONxKg4dgYJZYN
ezo3CQhL9+0sMQmbfIhRL58l8oysGqG9QT8Mk+bpmKhRH13Lv3cw9GwpqRUY0AXR
A7uPAra8wfYhDYx9s0FQSJWXH+v5EcDHsOXYDtlWD6SGjbF3OnCq5iR6/56UkEDt
BSU/fyA07YU2/1IZbzOD7vlrP8xz66gvTugrRYJ0wVs0oWOGOUVo/TFukVP6T9vb
5Cc0/eaTw2YiUqX/4ETQURIXWsIsIOiFbAeoPF9mxb2DFxUC5ZC5/9igvZCCnXJH
6spGmfaMxhwGh6jcxnO9bEkQ/EVB9bQovVVHuQH/bkSxSl6el69JvlQzRQ68O5ld
5VQhVg7WsZOmM1Hm0tXlL/1fGqiZoMi8OtlvjT1SJKO/1bcOVZ/WAqW3hS8WF6oQ
Gr6U5okWkDzuRNF6EqhgHZ3waa0jIS8Qe6Bpkk9ijlYGrQOyNxJtpXEHXuSGsT5d
RRJrR8l9W35FusLlTZdZmOC/0pefcwC81kKbpk95lbUIgxjS0b1gDDyz6fueQOVt
PPiUeT7COM0RC9MqoaXdwvmar/9o8t/yhbghoplhIMhaDUeNAS4oVDusre0hY9ny
7yN5c9wYJRxFpYGGp54JoKwcvjXwfaMi41nw00V7cqveSQbzbFV8EevqRU6hNnkd
W+ItjjlMBOHkcI+EC9Z/T1RIEuLvVYMDDH398CXH80mR3sf7Hqhu+vzn5J2H4jE+
t8YMp6dG3hsOJLza4RuRts+qRSiJgLTpAb1el7E/QcS/J0dF+4BSzM1NTguOTfeb
xAEaZOwKRxGr3R/782pFJpaoSYuuTdOAzFzAwh7lON42PzMyujQPvMmYI6q9UgxU
EwrgEnqoVooeoTuoA4t2TVrr/wk7NMItwDdAHxFDJvbDiXQWlQig0ztoGKswA5mj
7myZMTkzzVDLOYowFrfSXD7hrreWBLiyIWj1PRIoJA5EXxrU2r4mkxsEIK+At4wo
b0EVEDyjEH/sgATsVoWFUsfuMu8g5VbOGxXka158azXHnu0iER0CzHMZUbgxNOPn
mXpEZdjC/y6nkzmUzw4X8OM9abEMFWoqc/g2ldY5pMV3GB4HDdwQTxR+eJFdI1Wr
7vcGZ/WtqXyvsPa0gurr7mVDNmQIMZc2BZVSLd2y8zOU+ntQAJ82urR7uiymsbZX
g/e+LYdoIh/Uv2m98eVoY0xCltFRn1fLq6hKE6h2NQ1JIMMNshMHVd9DU9Pbzu2a
DYbDEAc3dQO9nw6RhZJiaQKWrOH85VCTg2jYWNlg9v4pPdPTGYIBx04QQ74JPUzK
B4KR7ioX/vXy/7EiSP+MfOPAzXGnfKi2CYjSpyir4mkQvo/HP973We8v13sR/mTr
6KZfmiC5G04E/l/SyVFk/CEMXM7A5DauQfG2umNW3PG/Dkq0MuhibU2WgxMkvJHz
3s5s76jhYd/ItHlsUfZnz6KzUv0cGm+rOZ6I5b3dQWtjTV0C353toE88Hb+mOasy
zdlGNW5gfxjv7llaBDEylgdnoPu1KiK9glyBXpWv3yl6l7WDWqoecdIv1lkW2T5M
cjK7D9trunsPy2VodhRCAqRPA7UIgTQs1hghSNj8HilnslHageM9CEv43uBzhRt3
ugzpOg+JBFkGzV6mcrgZ9NEBQEn67JCuwWwInNwXbwzB+EPXFrtAt18C1mAtPOHo
Fr9+BPDUyFpYnBn7HmCReS5NtZZCgi+BtXP/jFG5JyJEBCCC+2H9jqIqUigHRlMn
l4EXWZz7lds826MKzLx+FuZqiYy5FroltHu2nLalBbohMhN0t5IbVOR9guIsmkuJ
7cXg1qCsVHIaqwZPd3FLBvi7RVzADXirf616qxfSDh+uKjTEfVoM/XKcE6J4/2/F
xTYhYtJf/MjbEMPD63fttF515Dsjjmd82/W8qoD6F6Ew6UtnNQz+Ep2B6pA2SkU2
IVJaUk43+eM0YDIv6FexNHdMt1W85JS7TwnUYyYak7lpe+2Vr0WmYtQraz/bU/qi
B1n0IYuD6bRp5EMc4a9a101t7lMKgobdSAisVDHQ+I38UDW/lkDNaNTKQix54CpA
Zvh7sK9WNq7wiDUC9mDjpoZ1ggMJi99H+n7Ho/WuvXn+N1Wt9vxlL+yRaNqvxBfr
aaHrfy6hUh6GT5RUOedIduCARsiZ/f+M208o4Q9477xkXej+9u48jrxTkt14q2UG
owntxo1FXWvHMxfCaoViUcRSm5CNJTgRZ0p24Xdbot4JJrb3L5ofGXhN/x56okH1
LzLJqfaj3c9aR74eYp2JlfugoLUt8Z8NplSzBOym+uPoy+STUHntdPxeOoitoBwA
Eetr1NIJzQw55aRjCGRhdeoDW1e5ZhnrZXE/+gGVlqzDMxcBt0oYSNPtepR+iCNA
eq32UM903TSPlec1dZLo1Ojwoef4US43KlBP8HlK4Kf5ytcSnDGZlqP2UBjTgIn/
fKgi1uXWVzLTVd7qzL2WHdVRjIHGZVkX4DElyMTK4gntOlbJDlFaeyHtPyOncvJk
Sbdf8aLtRvm/Sm4O9L8zLnphKrhiqyH/b+NWtEsbLSjPbsBw5UaKsmYNifgFeFNg
lhNJ9jsDobDpwPBwXmrMVuqt6ba29uj9kzdeHGD4rpbbkWuXSliWA0gs+8wZ/bAo
ggVHnfPytQlzO33CBo55bIDliwM+LO/3lpbm9ePqqaef2sWhvc25ROr1jsLtw8FJ
brCDELFp9KvT3QZk/m+0qZ+xlPf8VolB0xN8pvuy4udqL/NvEP57/dmaY2TvieAw
LvsseI9FBhVdGJvVqP+HjclqJM3YtAEIPUka++KKT2XJIgjzbdyp8yAJiXj4DkA+
pS8IJMw1H9nIWXJJwMrch/MRO40DfUB7HMpNTAm0RxYs/BL0rowYPZImpzo6wkg/
3n2VgUPlg1T2fPIx4fKuv/CTWv3tKIkdP6dwUfiVJcgVeRWEGgVzo25cW2n2/7KY
WQqmc/YmtZxw7sNIkvLsuzXpcRx8sswzf2oQDEpo7u8kkcPRyawRl1El0M9cggkX
dFovvYJ21SC42MwycCccDFTMI1b7mbgBkSK5PrE54F74fSCjDpfcfB4cagE6bQ+/
5Y1fyeiIEiXh6azvq6Shy5lY3ttIkXnT+cRFSNe3gY8NkvULNjOII1Uvyq1EHEta
NlFb2FbgdQMplZ1KA4K61KraKkJ8J4F/pVqKew1O7VWVk/wy+NGbcaXJdkXvgcF5
1y2Qzi6tduyvEupcMETtzbgoQtTfNKujA6KeHGZw+ukKMG5UkjTNSkQssVCuqBPT
3JMROI6K1lsNGvL9NWo0VhxVZM41Em++k62PAc70Pa2cFeVWJ0zUEkcEKZgXmGoe
ZqDUCYk5tA+Pbjo+JehROXTXbXZNAiRDJvfwpTkZwZIxXIKK/TRkUtF4oGVdfeTs
r21z1MftnO3sq7QRqQqNQsNPCc3N8aKerh/QAc+HjCBHnf4w34lqFJw81WT+6IBo
Yhqt/r6Sg2jCT+ys125yoIHEISnYXE1B6Pe3+FZ/1/ND17X7i5j5yWmhHfXyMAYC
oKVWaZMhpgUJQsuheMGx7kg9/ojYQeY9pB6OHf3FDQ091hMbmI3s5zOQ4Z0cdGu8
rR/2JVQ7Uqx04UFM5LyJmuOuZjakC+xJcaOzd5yEPtUMXQbeaZxYJfEep5qg75bg
baYg23gxJ80sBQotEMT4aAoSiLKrKfMmdolJ21/CuzwEFHpWz/3SBoeRdArMWQlB
vrSOlwbP0MHuQUd9JvRIAAmtVLoiPQGCG9po6+Ehi/gUnqlWoRI9NwoLzFsovYC2
rMODBTNYEUpiQfi1INwmy2nAkcowBr8q1UINhY0HbXAeaKjukmCJTygyZR0pZG8G
AWu76lsR4EBuF85XJRO4uOMh4dJfflc4COa2mYoXRdSRBS1Rpj2zf3tWS0cAvrj3
Ax5YltUBHKanTDL/OCEnYRAt6YxDdXSuAqnbxmBwCInzmj+SBJPAFPM0DSzXTLhm
zit04AToL0/gMLll6zjs2MJuQsZ2IOkWcwNyge2Jxt7ZDex+AtT7JWgPiR1OlZFL
zIRA72mQmSENgPGZRMRJuJpkvKyI0vpiwN8yKlUXSEym5Z3SCPidgrWVtbZAKivc
PATpJdFMU0fXnkE9lHUiyfiHFIVm1DCZih7Q5vkcN5NrPEn/ZlTT2+hojIwEvY3C
kQ4/wmZko4KnJ/UkBFVx7Sbf+A40Q5JDG/yUu6KAKlVli9mmKOEIxroGhzojx1ko
ww0t0PfOAP+IVgkbnvZ+bNJcakhn4axsVTbJjYAD2l42WM00+sCCcm945XzYsbt5
4a0k22K8rnMrgelj2XIvbyK71sgyTXBcPEME7DRFq9ExneP2/XaBCiRh/W5U1ynP
adrprdCikEJs9mxri3YBfaAB+Oj4NgX//nOLnkxsly6bPoOL9XaSM+Sf/GLoAnKR
xfdi4mWn64wrEvIh/QHWnCU6WKd6WcByi1WkPfpsjJ453MooBD5j/RSq0Ut7wgsX
xCC6qiZnh96j3fnlRMcfIjuo/JcpFS4eny5wXWlr6bk1aZvw131SrF6I6sFf29I8
ptc1x9r27p1Jbv5djIyHGwRURHlAWEQ5l0ltduO7SapE8iup+bOQXgUifxxtcLU0
THPAbPB4+5SNXI6te2ZdNZE7CBMKOaq69nmKd1y5htd8i03QRUVBbBVxSTKtpjis
rlzfLdgQbajgZB0okuXwKWT+Ss8YUOJZcZoQ6RUwpDFJV9I6vd+4G6CddQLPlBkl
3Ja8DpQyMc7pbMCcgZmNZymH5ScpX0XPUR/8dL6ut3//qdV4haUu23/SWF2shK1a
FDMQx32/N1I/00tXzbH0M+FTS/26vosPw2WyEsfp0U/U1SKH+HWeDe7zdrB3s1ig
LopPKAMOjV8e5cyivmCuDCgR+qk2aCzaco2/GfbYBBzgfCYmZzf9OuWVwT/n/b4A
qJMIngAt0A7zInjHlK1bOMJAnO08H2MvBbof24J8pmMnzvL9JCCk2ApAgIcm8Pys
iYA71wETn95swpONFmPYDcbqUAf+WkakU785H2kLf9Io9bJ4xbGnggE/TUKNsNeZ
IJKs5RlY/7doGU9wWCqzmQHoAanFeiZlngk8pHUlLRsvrnXAHowjQkVBkFO9toWf
xrzwI30Hqd3yGAfffmoO+D3ttpPN0s6z4k+bt8d/OjqkgfjrEguIsNXiUgds9Cag
FokRIL+crG6LwK7ZPLa8pi6gsJhNkD6UBl+4bu4bc99ohqVyAA3f4cCBHKKrdD/p
ny/EryX/74Dzl4aCyRPdmkbLxipiY3PjNhX+AD0FBGD1S/aoVdS9wbRcgbe7eqh7
zTsN3zWUCkyLhS8v7ow3auon8jmzUnzpHqfCFc1id6XCS4CLH26fdVozoOJmS9WA
Kkiw6IkgPq7yaOcbLUPWV3EkUsXeFO1yw9+Bp4kYUAGXALPuy2mXIw0IVjUSg2sE
0HlhQlUrFVxHvxNfUq2tafeGddB7/JUOtMo+7G9Ybwe82gjcGCJGBotPo/CPzRZs
Xxs/q/EqBZ/I7bYpSOveIJIWb8LdiRaSjRpedkfLfyJ3e8GSs/gjZDLQ3nV9vYNU
hbLBYU1hodbn51ZizRUjumvXMtR0+qCvZC7xWUkIfKJyMqAvaSysJV/MRVQpzHWs
QQE/x/2u/lxw5H0qAyzvj/WVRsltJ1r/36XlpPpzNtWPAM0PXmuMKhBmH8g3TGk8
RIIwKM4LCDcFBC17HRcmaaVchycr7HgpdXGnUXy3NvPXhwGEywQILFLroewOFbFa
mDx9Lz670SAh6Sx6nTYa/VILQryvnKU+tnC9t0qz1YzRU6wYCdtR+1ubuuzxSOfu
v9S2np5WCNeCT2YBCQWfa0Clapf/5t8+CHl/H8Qc46vgAAdG4ZkcnGgxqgiUEaHn
s3OjsQU1d5VEb5oKuxb5uptk8IIoDD1d2jUZakwMCSB3qv224iOtjFOFsVliWG4O
R2K/NxrVrQFKEuGHno2GhwexsaO3ZoPPKcCcvn7msf0bA/PIxAn1eVMcugjEqRrN
jjDEi7tgH+2hkMr3UfN9LItKNgffGKj3JRyTjxiqB7vJ4o8XttUcG0jE3tRLz12w
WMgcEzfAafIlpaDMg766yz2uK9jFzkV0JF05R2li5NELmgFUmODbAeFQFXr9CmVx
TIsMV7UL3fPAW+Ioy14jcIbxZin6cyvTOsCr7NPSqt+G4YxSHEQsgF/42bbg7lez
tpycyWyZCJrcYXrT2SLxWyMOUlOXBDaPLEDVD9B8cPUxbFWkBOjs0NuZ6F41B+Q5
9PrMnfXC1Zd172yr5voUqjJxNg3DVhOze5NZxOHRApaKZGd9Xj/ESkMpC9rW+Iav
eDjXUnbl/zlcCJflsP5OdxRmYqw2nK1LDoW88qoJHndcubJYzAks1a3OELcq0FgB
6JsvVWzdgWo1Tvll/edZuOoUdhsoXEOsQxEmAl+g7DWkYM3ycyE+4wpd3BkWT4UO
OkDyvVTILGDlRg67TkSOzDhChZzwn8MhfinMy4mh7JGBUh9zqQCSJRyuYhho5+6d
PwAdkhDU4IGnmej37nDV7qI+JmP2IVfIUjWYa+erxFb5IJ3HhfvV5I5p/KbLewX9
EMm4Q5f4doPnZiZDGes5UHAqh0wvCeFaVFzpkahgERnRCFZ5Ipgo/bdhcb8vk8zp
nrOrT/TZ1FWIPNLDgfTUNwoyBYOLuh7uw+ebhiKXGHiAjbL3nCD6rXu7zorL4+F7
oaq4tw+BGVKjLdRBuDq0m/v6a6nsGMXj0nCq80SC8vmQs2nbf3dbQyWg4b4fVDI4
wBKc3q7ucMEpzHkzIziLgcRXkJHS79ckPEbNGaQFSwWocyePSwKtppbTXm3MRJLK
LoYE4CWz6cjWSYuh6/JRy3R2eNDHDULsj/YjTFUF6eUFljY3DiaJo86wQ584Vrmv
0lilfuCZnOR5HA1Et3CZqxjwpCaNfL0/XNzJgk3dFf6d4fljvI+obZkIcDRJxQS2
U660aOXTkMr5Lz3d2zHsUY5/RIXXfsRYeg/fOQQwWogpAEz+JXdgbuQmaCQgRrRL
Ky8br6YL29PHOmaMW+BcqCWOVY9c/+eQkFjwEKmBUBrPSU5HbTL69wVslNKSOeBn
G1WtEMGneRqEQy0ZhHx3YA6KLnSayMU1NJwv4xaonjosmwsJZJ/mAhIvCrdwiGiw
/tqKmXPSjBg3kFvaZwhmiurUDn9E+Pg0bdSKUcSk6E8JkCZxE4DD3oyypHUqrfQb
+Pz0HUWwKGWZDT60XbLoA3556K9zgwFGyP7ic6WwaOoFZ0zGhJi30D6bZEoWWvFi
SsaN1FvfZm/djdT32M8/G5EfCQt2lkdRKjBGG9LXTfb5ui3ojbITHVrBntHQMD/u
uR87KtUQBCtBv7IigTKzYsA5ZHDPoL4D78tIXYV/ucDgvwcLAl93vdIEPPpHxoGY
W0nehqH6WTx0w7MH5QhqBFrZTXo0Y9l/b8BelrAmNhoRNN7nRcioslV0nGbgeboy
H661W22RPRRIgwBENJ2TJqdD4j4lGM+hg2l991uHiXOjnc9LLikQE0/qKA19OI+w
lh7j5U39yG6Rv3iyA37YYV3ZJiz1+iBlCDWJxLaQe27EJWYRX+FExMQk+gWCXCO7
DZnWY8HBnAAyX3vEUWFL9G5Cb/04Q/TPSS1Nj3cazKn9tSmU5vH5tT8v+K2iCA3K
zw5TDTLAD+UvL4V+Fr55tlUQjbat7MjFiY+ZJeUeyEh/rYJgudWOLTWo/mOvxtL2
cvJPMpvRsUXwPuk4JY+UV/00z853wbSM9DSPyliu+iMo9VerJDiTMK/oQ3DRVa40
PKvzwqqUCe3QD4nF8W9TRehyJjbZMqwJVvTs1r2c8uhkmqwtbiH754MYNw8jsZps
Dv0JVWbs1I587UTjheyUi14hrXT/mYSoymM0KaxhbRGOz5ldXhXaZt1r6dSBF8Op
VPK+TjQ3QLmJwQd0b274wXswAVYl3aNCXxeCK7yJASnQlDSDaf1Nq7ccRDbROpbA
GynZ/wT5FSsdpFlRq779GdGyhgQV7/VFX35vwnxMKTSsoO7rRKRtbvEo6Y3Q6jv2
xf4mtIiG2EJZW/OAyhKCvKRPUTN2KxGhJGRAT7FtuoRwuTGM7I1YnRFIik9J7VCc
ddjk2vEjhzl6CSiZa3lwzs5dsq0Oytg4nDrVEe7qlaTaDoBcfnsy95IpX19rSmJ1
X7ulcML8pgJsgL7bywEcZ/CcR1wS52hilLuzGjsyZLsIPuomhyyLJ10fQTEEKWfS
ubNTxv1YALNiuEVxr8ZwLJ7lnfAEw060mNUB1Sxix8lnZN1JQkeVEbny0QSCR4by
Ln4fEU8rcAqoOBpWH3U79vPuXRJkMdqbPvb6K3MGBnRE7Vj+0wE9xqq5+sRrrTLi
VbV29itzB13VrMK9Ih3X+++hq8ByfbWGG8twRl8hI4XK8Sq6l4qYCfwKJV6c3Ts6
QnWz6xAQz6eiAJqOUhaKW2rzWnXLZRIjC4k8WosYJ+OhJ16Vxh7SHVfFx499c+Fc
p46L6P6Vo5MnH3bBtrnDqq1I9FvtOcfcM9zCexAo6D8eHA1AXg51boBlUqLiYkKW
Z2I1gZGaLo4vfApOg7Q+U+cZPuefdRTLF8FWJnCrAzDP/f2ne2RXlZ0whrNM2nPn
JTMFKh4gu82bF748Fi5jYESOqzo109KMJD8WREVdVpSfHrQOOiNYpyC8O7B2l0Xq
OSEWvl6nxU8DhxnIJ5EIYHR2VSfRKSFSjK1CPMw8RqISpA4pGdsFqQIzbwjPe1GU
xX78nIP/yCGF73kAZaEo0sCd2YsIw1cEEDcYqZE9zRtPXrJq8CTKPAVRoeXgzSWw
92aiwN3i9F2jrNEB/SYf7u6OIIgFtOMDhk8phom8oUY+yNSnE920TmTzSii2eVVo
z2k1LKaV5/vKGQbMSwjGiTf/l4G0Ej5b/fl7PvtuuozZQUjVaYT3YFaJOrj6biWN
aebukCmRggwNurGy0zHga2J5fkDp5P73jaHyKi9CRo8jOg/Ib40iYj2M0QBRTN3v
/jFNvfYWjJNwgrvfLwsB5jdWGHlyPJrMCnMEwi4xEj0ZHIqZees1HFhH//CPmift
KW1BVqNkLJET5qEqCc9+gymAdtWhrF7GJiqSHNQqEU61CQVgpB/H21GDNkX6vVQq
Pld2LbZ+3venYteyp724CZ6sTqOW9t7rNzVF14sau+fOhaO5faVqvoArSyMp3R8R
XKzVqrvZxbUiXJIcrvGIlkkVSRTJQddDSFILs3skIhAxdIwyE/YFb/FBnK0qVFba
qflmn+y4vwCTVtbk3ouPoz7RBYcD6UurCrKBudnQvByKuhFFkslJDjAxV25zCEeB
Fo58q2h/hWN2pYkQmbx8hw7Zd2hqzU///6O0KiBXG8EHEfNDS8i0q/pIbj9LsZwl
Z4EJ4Fcb5YzkvNVH726J/u20H3lAKNI7hEQX6e7pCo4=
`pragma protect end_protected
