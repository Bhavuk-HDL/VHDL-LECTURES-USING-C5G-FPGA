// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:21:29 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ecP4KcihwAKEvIzxEeMwTApsrSNPLMChAj33oAJ42fLgmMwsceZA8ThlTlRlXIhk
k6qixnrLUyrnoQtANQo/HB/tIZDt3GkQ2mG2bAFd/mcJg5m43+rCwkL+NytFI0Bv
seyFIV1TtjjOGEyWhKuF1vQXmqXCJaE6yOZZhR9NJoA=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 2816)
XFXCMcuGMoRTbhmY3bDxSMEdLsRhvWvNLMaG3GutGl7kB4mrLFw7v9YXN5l5P/r0
YekGc8dEHdYOwrrxhnnyYWmPlKvs05njNaGD3aTpd8l5H6t94o0cKhpuzps7WEga
eFA4Usj5gurpfyNM5uJ6DU57DB+YHVvCNcJgtxBMcwg8bbYPUrrvt8FQUmosb4hM
qT28cg9Y84Q2eJZmUCdWmYoxyFqCaIcver3PlWUnv44TBOu0xQUFxV0pA4N6VTA2
5Y1nSaJBfnZ3K1g7vkUG92SobYo3cxD3bY9OqQc9SI1iVpF4Xq//TVxynYCwl8OJ
PuKWT7NTsvDYpl6U0OAyGSVKxU5cwt0lESc+KJ/Z1Vr4HUMScpm9PGG3hAlIa09P
F+QBjkkJgdDx+OoJuQB/X+4ECcEDaz1jwi9QS65wenehdQprE9srFYPBaecqtc37
lrJyQPut2I1f2Ri+X35xlJtLqbfnCEjOLlVCg6kmZByTs1eYotLYMD6E4m4GY3mI
xNsIcys08NM53bky+q8/tRqyZsnFmbTCLETC69RDyXlFcNLXm7DpxYJcf16kxr63
JkLSpuK9oVnRLP746Lbi+FZcTX8jvZmthSJvpJRGF7/9XmgtcO2dE2YAYUifWH3T
bADSPeIK2rnbtWXTUCJTU6NOJK8Tb9cogiVLfJ3Ian/Uj+DXzpup8iHWr2Mlx18a
yI2LCH8uMH0W1SdayxMqIchtqIIZWP6+TN7L3EBni6xg5AvCW4yA0OeLgw4icMXn
ITkAvKsEif1Trfu2OuTmhaOOFujqd/honcmjwCBzRL3IoQZzI8whVdggBtkWSLgD
OQflQUWH2XUJlbpZ8iTB04bfXqNkUd3x7sdNXeeeRUR+s8NppjMz7wqaUl1/5YKP
GsIQHcAwpZW647/0/dsh2UDjgULCEXFxxdz51busxn3i1Nk3gd23Rb2qfLSnBgp9
GhWGjfPv89am4JyUgk3NkztaXF+uWkyHsK3vjy1L46XzaAUPb21rmxJVy7/Bg46i
pFFJhC2YGAFkjt5Ue9M+WvIgxLXdcjyieoZKpNBtqinE8uBHJDCshVJFA6keAceY
WgyKaxclfK5v+gxTqll0IWkXbw2o12BGQXNqBYL8f9YRvCn771Z51fkY2nhcg3gd
+roOvBtNXnVSUHLxYHj3p193q+elRgSXgMh6/xT+8x11sAKMx+D1ANgX1DucuCzF
+3ywc4RebGH9lSfECmLEo2tWtLgjSa4zvVgQzc6UAt95Gcr3iGlr32FSChHTj3o4
z8pIY0XlMTvHVo3yL7cDaUFYzQ7K0T4lrenDpaRPkfKyClD/aI5jFSkHrhIZkLjB
aan6Gyki0HINuIW6upP694oBkH6byHGDd1uWawhMSenQdHv/GYNWC6yit8KU1TUA
IpLh0DGD/d9l8I6LGVpO6TSUyqUFTZuEUKDHyu5N9JsDz6K37C29bU81O0m6nkQa
QF8uZz3xGTncNTgEMuPoB/sj7tfQOvO+eo8mUV5sonn2JQtFZeUodIGgHcOTNSNe
DDnSP/XPmPl02+/wk6LyTA5MkDAyPe6Q7S1Sf38zUm94Z9nbVnQvi4CFnCN8kKhC
gCemV7TJd366oXwfcPPDKDPjdTBb3EeQfm+xDsHGjWSJvphgPuO4q7VbLvy50Umm
SssBSsdTinnwSNoc1xLx/IonWyQoKNbp+nNprujDRXIc9xNydL9+AwHVrbwDuCFz
D/M2T+FZ4waVNWrtuiym1Oq6wenAbMoTKOqVL6kG2w6P6tNXcbfnPSRZlOTeqYI6
ILYbFTTYzl6gCxVoaiJUHwl3vHFcP0VuFdfECnTGcbyaHNEAkXBNJRKOlJqYgh+6
kNbPF+bg5W+qujQYVQC9NlqiesH6lBbROt4HKB73hVSmCUPlT0hm4mNhCtIZB6j0
K2MGP1ZKtoY1lois2RoZniH4eVF9BoElrDyc41UJ225BwGnMadFxnfCnu1XPby/i
ncgbwk8pZD0oiY+SWW9UZuv0dg7t3BJZHuZZdc7BcGs/x0mo1NYO6EdsIcIE85qC
hiA89CXZxeTApu+95he9lfYuT/sCjXSZKevYzXO60EpM0I2pmlaPfcUi+jog1zIm
Q6mvrPwgT6dM4CwgTlVokmlBovDAwKzjOfrnoSVZ3d4RkfheKwDjvlvWMR7nYa+q
/phAuzut39nav73pEXpfNKCDA/p/2yJAiYp79CjF6JHVZ+vfJhSK9pGX41y7cg1n
yBXWnFpAPuCUtaatwRAiV+m6Xp6T0TWVgCQGePLQJxXt4K3RyJ0+O4wLl7/yjCf6
I8DiVcZwDl2Iah4wTcbIGh3/S/+JdPLtOQAzGdQwz4toAuB3ESew4X0UP9ns7yA/
vLAMPPVeX/L8eMVIQMYVkzBdhfJLN9bD6deICpUgVDvBQejitJSYELtAeYr7iKTF
g62hr2iEjRlNXtpOJh0UBeU1C/WrE5vFXYcqUEAU1Gewmhsw0/Limjr/LFgbU/Hm
IeXsQAKB37WRMFmts1i+e57kqTVnGYYdb7qmao5fWbmFCV8GbYRfbeEnU3G54oH6
an5WOrx/rLVief4yRvAw7deMloZvX+UWPY2qs4hsM6ZfF3rG9AODSIBGtUDqbkOS
tDzx1RCYjcWqrHT2C5mdgEoOvJ+X5y/kEPWCZvhHAmBti9C+XBJzEBLfDmDi7HSs
FXxPpuWEWfXyOEJHQqTjUA+COhGl2Mtx2MmqqfpTAYpb/4icrZpeusZcEYyhrGGc
Z2oe8CHyXl4ycZrUjQoW/eVqD3PIS2d8FQhgkYHUbIjT/Vhf8AGfgDUYcp5VzDmH
10wAxLcfptaMX90YunVOjdHDiF0/SKMFzTmH7XWM0WXY8czA/MSixp9LhQGJj45B
J/0Gt0xb3BEGmTi6YCIZRSyuBgOGp/5V2eSp8sH3eeVxd0f5sWt5/QcSoW11Erg1
ZcBr9FBhNdsAv7ITkol6iM11RnjyPqoCkbaTzJzJ2FryBWqE0VmuO3hPLRuP3rZE
qXzq35ol+f1j8JtFM3GxYzuzWDQezROQSO6Z8GVvqk5SOHROn0RAhG2uwYBsPNRL
riNTQDfoptKgG18WyWEBKSkn/8IQHzzmEhn8Bwn+JU2sYgYbaN0cQxHZQOoan6nu
cg0hNCRmNy+dFsi44JzeozpYXcKdlHyteov/RfQCHCkUTwYu5ordR0lxJwa90jaA
apSo1mX27ovGfNZ/+NAES+NTDheOxiCOz+JS42kh33N/ukKQor/tUdZwOXrIYF/P
i+DuanS4NyGtpOVbDN30n3UMBARyc1zXoOSX/ZF5KGyZcW1kbStzC+BMdLfO7bbI
DGw/oZn+lRDWkjuDeCluIaRCbRl2N5ZLYCrwzxDH/NtJqm1dKezc9wmqLwG4a9hY
7QCcVh+6VmVqzvDtx4wAAHugWeBnjXfvnO1N2qMtyMqPb52JtHsRiVE9boD1a73N
7Z4dYq/OROuv1ADJPq6nHWMwvvChaoA1U2eaxLWS5fZiMej7fbQ0qoJN5YvTYCs0
7dKN/rkAVHR7H0ibjax5u6TuJb0d7BxFFiP4JN53pGub7RKVUNQbDatvcMbsC+SQ
+b0M20EiOm1s0TV7AX6me5vcAVmbF9RMGz7vWWFYGk1Dev0u+z6DzzbGCq4iEuZW
9lz68xObvyI1NaUFIOFM9fAY/i42SHnlVheC+PyTNpL36XODpKXmNEkhs3tyH1De
ucO9ZdZPMNXwl/WQYVyEVCQMw68bfQnRR2kQu2NUVGk=
`pragma protect end_protected
