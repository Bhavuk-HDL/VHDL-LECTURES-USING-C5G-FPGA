// (C) 2001-2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files from any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel FPGA IP License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
K5Pr2SlI7Dw+88CpgP8FVgSnTFZeJVmlSz/ArZk4ySNHCRooF0dERiJh4MC2Q7GQ3/sghIDuin+I
qBZKhW7JeJ3KRE7hLOj7+W8/dqZuPxnUJ5YTLkXrDUAbDciwpZ5WlFtMMnkp/JLCPBkyITdsBp0P
SCFZH1FcAkjl15Bysb+s8m47cypetFYKYNRc8oTKY2zZyLTtiztqK1I57UV90pQepORhlWhupTLe
6QleK6XHFN3dHtKGGa4etnCLkvlcGhjr1pH846JvKA9oB35Zjnr1NFLYKfoXqGmKrUln8ENI2ean
DFHz9yIpiBcA4c4bFNGVmU5pbMrdmeQNOrS0RQ==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11392)
aiRp0PKhMoYca0iooB+GYVPYHGJOStlla3Y+I+1rePVSnDOA2pitG9C3kv9f5RJJmcbWEMl4rL+/
gwChIEz7vGz12w4IqkpG4obPeJP5Bv4EFBDlkt8xMrO1+7qGQQJDTJLJLJU7gqu9HNNrsR8NDZBc
l0RqWxlhEkyfvTC1IV20dOzaN/jqtnp+izWgRktkUThujSupowVrFqA9N9ltD1YKW5lQjpenbYpx
EkDgSkDTfAhpp7NLm9BelFVpYfZUGDGigZhf29SwV7Il1OskD8P+OO8DyMAlM68hyBBWZhrrI0sM
wvpReg7ZcM61q6BjD2xIEi5ymXQMjJ8H9GQONoy/L/Kg4SJAgPYgosp67ngbZxoIPZ4nVVFA0f48
Zr/ATA+O6hQ9BE4HyM58ZvUrBstvP7Pl2ksrRn//qGCOkZEm9Jpd5zOaDbGoVsBRDQdIr0Cgl3PP
7RyNXaP+Ozd0I3SycUvYUHjH7sMMb4rlB+8f10WmNVnKmUXk2AHDPmAcgxBu+BRCUeEzC/Kb4+td
1JuwmIVHZpZvdXGuXIuu/UIQ1eR49A4JYgHpSfgJcOLdXIUtE1fsdMjMFlvtq5o8CRp+Qqqg8lIR
ZjtcG7i16lyyjX+yk4MX9OObhWL9co1l03zWmVK5PVUXZ6FLGHr4F3dM+W7tG/SKFd16I1cf972L
sjcuYZz6aIB9Wl1Dsh20Et+JBkXH/Epof2cl0YzSE0NIArbMrcQsis4mfEHy+cakGviQf7wP4fsZ
BJcTWSoYBLg/zhv6VHcpcvO1NYaZ5uIjho6+ookDQnlOYVa/GnzmqZa8yf8TM6+8VV4h+A1/Zs0Q
g8UqpPzQSg6+vUipsv7GfmiF79JoFBo1xRUpBpfRU0tWcpXu30IezgOnPfTixZlb9zlUHSaOjYF/
pZNuVJQzf+FMWajpsAMY6LjXWfSOobwlHQeN8GCuz7o2lLKoJ/WjGJWjUeZo16wQAL1IGBBdy9Fo
7gcS77YjTYuJm4Sk7Kniz34cfdanUxDlQ/Y7cWlmJIX7B7M04uSSnNeoBonTXYRyJK6Ui3IksC8x
G92+HHgxhqwhOkf9Ek9SW8Y8xNo2tPegWTysQCbWxDczI+jXeM0cIcks2M4esLcstnX+6Qa6xlNP
U7WvLg/hA+EYsGkhqPUNymXLIZlL6ow/qXa6dZOmFrlJzsdoYt1i+O00Gc4KI2os7SuQ2w+qTVmk
A4bZCkz/XhlYsx3S1Yrkf5Fr4xckWSZQl4rbh6k8AY6B6q6nHOp6UuJW/k3N2I5uUIO68+lymaig
ABrvA62T8EaaICE03XOV/XWSOgt6ayJBjAWykogbNLHjpiwS5/yufbUkG+fEWqtPtj1h4GAIj47x
Xc1nOaGdEzhwM4bXIZs7ChkqILHGSgO6zc3P0Ble+w45D2wgpfHwpydF6GncsT6N5iSt+AwdKm5V
w+cY7VSeJ3gzvktg+nmfz1AciCQMxEr7Awe6RPW6wbbabqHLXWn3BmJHABEnEz4KjTRpGKDjG/55
dkX8puVG2KJxSN1lvgN9OKqElEzov14l42WDAdEcPOvSmvoA2DBxPwZUcxdRNqSm8ybdpH24xzVa
j/bXMAJuQRfDS4ewFv3L3pFLxXHgP9tMsfLoVW2vi117ZeqJFp4qVBeTAAIfxv19cCNu1DUng/vv
jeaTZxj57YOLy68+TgAOtUUubFNn9AiSvav7tZ9g6m+SxE5D7za4vhhgDLG2zSsi5cJEcshXWw1h
BDKFDgf/oh+3dmy/IdXRyXbY3vYm0q/IOj/BVay/vm+JlUibTCI1FTnoHFETrOtnl+OXVGWAye8f
hNpxuX0Elv3OqRsSnzHUMm6WoKLGBFRYQHEV8GzovwZP1ZlXmASPDsrYdIO3YIUA6nOA2WXaMBXu
lJBtuCVIKZvZNFtdTWMRmV9A2dMXKaS/zKKQnQ4iNFtpk06rgs0s5jKCMqW8mnds65avqsua19qB
tdxqu2bkODK35i+zGnezmpfc1cqmOQV2sb6z75i4ovRl91TgqngTvV29lPvE4cVkcc1JpBsmzOIS
jVPcBLqaGW8iywclBqG0CxAxgYjtwinrwGfyP4qKwhQmqHDJIXfDbwMRJPlEbEHn+I/blwssB+Ot
Vckfq7WW/HmS4wHgyykilXZwF3X0rJrh+SM/F4MxmxY4Z0sau0FTdOekrM29O9TYXmbwZt0rXQpg
kU/om7T86s5cqUGFzN8nhTwCuLQRZWNg7IyGt/yeXdAKy1pA2wByyXBDwtJYQLQX4YzKZjaSmfse
ZKqG3GJJXCGXJjS2aF/lQuYdgd4bW+J1miHonCA2WDNNRU/fxd8aT8geItJWPeEdTxp6NXfFVpS5
KbxHSE8lJ4ngsVf4sfBVYlA6emCmXUrN2U70IlcRj6r/xAGy1BvviXM3Rn0O8mxgShG3E+rDDZbM
noR60GYTYyGYhpG+rAZ3mxuA9pR6SakRVTYEz2I5OMNgEjGkwoP0aDq7xyCSnHTCZID4JEL/6Pb9
278fi7ftrI5axXZ8W0EQtVPka7kl3fa9bl4g0WTt1KoPJIqBxofxmS6WguUj0KI2TnwsyjBeyac4
MkmQ+BdCHG8VcQppY0Xuq4p8LLQMnB7o+Q3l8jI/fU9wl1g9a1QwjrtuSscaIffY6jRGMWEzJEDW
U6drqO36XMFcFVhROevjn1y3T5nummWw6ZFb0XVFAn/EgGmIZt/nK3r+ZCcFZJjaSxmxLE7ztcvU
6Y/MbovBoXFAA7WfbubQd1a0NoKPUWtMI2q3knxdbGVkBUw9XcPGRmxGLmokxOCjPyfCARZHXM6u
xWsuRXtyj68sA6f4G7yOP9RM1Qa9RIC4NkkZ22IAC893W9pCASuiB6olg4orgFtAJpt85kgtHpbf
0/cKmPsT0+oia+9/oY+1zMLvHUhg9TyAAAA1KCMUmZaISJl2mCsxQAAMWHz7er0Eeq2vNmlS36px
52zSNYRu1NIGp9dfUM9V3g8cZiL6MZLqD33Qujqch++HOQDlsgp+D572Z9q4flZ+EcRIY38RWan1
gIWEnRfSmOWlHVEa0mRo03Juuv9XFfx1n/PBRN9jNF/Q2OlNbJFYHdM2JEA0HTxMCDrzRU6Dr32B
aLuLc+jzzonYH3Emuywb6Kcuo0nFkDytQZvvoUrUOjeeUvMUkM3nda3PwYehkEW3iLnE0Vut/nTq
geEWXfKKhcJRKMYYTYmz5A90fZdY5RgfcUJlSguVDHmGPU92OY4RckFqSIbltdpddN1aEEzZM0gS
00E2g7Pq6b/C2VfLq5JDtC3USCsq0agE7CL2XHKB9VdWPMH22PMa887i8bVl1ZQVhfxxc2smDxNk
7/OgvCKdURCm2et5hFQm4uYvfgIAzJ+0qnIVcWVlvXaQhZ1F3Y9wMJdf+FXLvjw729wgyVhIVzvP
dyRZEnSnTohwZpZNd5Xszrg9vI5qyflQkCJjEEr2r+6HmEWGeJ1yMOdu3JdHk22q/VI9zt5I8HzQ
pF11P2H5hrZDPPxf+9LK0XxxLX5g2rn8MwopF7ZwiGw+GVAKpzjYvViT+BSNYU+1FsWnTxaQR4pv
Lz5xXgnIr+b1hrp1SkA35JQnbzgK/ehcaHyeXYTNJSZv528dIdtclej7M1RnJIPE2W4GrC2n+KMx
VF9Fj9uKq874wJqYQKfETv/q1jU+/72OXmR+UxKuqpEVxKmK+rndRkFALuhGz1FNxCKLLCEl0Mdm
8u5iJtIr8vULXxxjcJtYLu0tiDB+oG7JLiACuNP/v5N9juIwNaZHhL/0gECp7yYSDlLsKVpvmIgh
4ZQRE3LKR/qIdjIBctRXJv8l8H1C1ig9Nz21F9MBhkM7iXgH9BLHdNHV9zKzt0hvswWTOsO8V+Tc
hA9iM9SVojV4FFYVhceUSr8rqwMjEWpg7cky+QuDKUCJ7CfFLGFDwwKB26+lMQPAfPnIg7in3Oof
QnFXbEd7BkNus0Rig5rd3MvHlY+F2Hjuz2DhRGRaeH/OijPUP0d6Vexr1VraCOyOWIGSOz3eYBsV
iPCnHLjPYoMOM7BplltxM9lbp0viAcHGre3sj6VEXCTyLeYHrG/SJ3XuWmuArAkr91qe49cXKWA2
n/FJP9Y7XpWH5o98brX3aywOJYD/CSXI+tJ20WI77G+wMw62qsMfeSaQGs6ByyCE5RgrW/70rfyi
FSBkHItTpBDuDhEefGwuhqIt23ykkoxTPj1ZHHStnKpAnLG5LAwzkjU8Bk8GRZmGQI7hBgGF5HBH
d+0L5sQk/OU6f65LFGT+FGfAD4nqmkeLfwx7U8DFW8Kj7Y7bA1/lx0vQzm8MHvnclHrSkJQi8w2r
MtQ0kRzuE62MDwUW2S48uqSm7idK/QFmxKGqgMUpfF+BBFkrSmqjrj1xfOJCYBODc35rP2q87cMv
qRJokOD/TPdItK8kVagrS+05/528+pqJE/kNQQIpQ85+OJ23xy0UT0UiYEN12SMCWMdwhZv1mq3m
PiuLaBhkcYdp3AHRqNLitz5f1rC5BmiyeqRWelD5h3zD3TWa5njviKGUa3mI6DgK/ZbxghMPXn5y
QJEWAgTHwAKxMkCOm/cHxiQZnVkoz3i85aoUSAjJeDHVa3FqpqaJKK7hzd8cXqTOOsC22/a6EMqk
T1uUPcRCq0+15wCW67aVymx5f3EyfIcIddpY2t6BOj+KqgFxHOS4hfps8XMsTkKTe3/wsFzY3s4K
lAEaZiGL762DUM3zCFoaFbL9yHdPjnk1edWcipbSk97XahpJn7zbI5AXAd83pi76ZdV20gvD8PGR
3wVBbu5Wzl2ubLl+2Jz0RwWUwsQJGY/1zh5cJ4EeR7AiBegs3Fq2Gu1wcgtal+NmYsvOQi02tRme
1rFlXwR8HDEGB0B3rz9WhsnuHWjGjC+1YCNqrlcCUF7ebKKRUbmFDwggOMhIpL/LHK4eZlQxV9ta
CcsIzFZ4WYzrDJJeb78QHuLXfPQoOeMrwoBfM6FHhj6M4ltQDiVZzmAXvIisR9YgM+w5PpwIqpw4
KbV5vvhK+IEjYTw6kPxDEb1xiV4OPn9oKs/EgWkAQRgHyNnZ+XuQFAA6FyWWUqf2LThyaY1m8U2c
mxssnIr4He87161YfQEa23+qMt1ja1JOYtIKdHWGqcFsQUttppYaAoBQeG3UOxKOvLmSQ0/cu5K1
QT27kW8CYk1sCJPWrCfno96Bd82T2Meu7BGS3HW1BTfI3lQCSj1Xg+FtDUteb4B6xskETaPREzqi
K2rIbaUsr3IRcjEjH161dvbN6oTPlJYk4rTuLBNpH20MKU9bGSIU0VaK2LO5EJBUGgk8dauPU3DK
p/C7Vt87EwAydDc+ITH7JJLN+5/qfIovFBrLXqfiOfZLGALuA/PmCg0y44fSUux5/dQxKb70y8Rs
PKXsuRRlSxPc25+4Cs9otf/+RSLNr51wyvvwY46Rp1qAh2+forkwTdK6luQkhgq6wfe+4xr3LoVn
1p3AMSqK/1jwzVfXgFTIAZE4fMy2HOkWV7/e7L3t9ZbX4U/O8b+f2iXulUKDNSY4iETQfrWWEik+
BVAweG/awvD3/7QnFe3nVfCeWpDAVu0PHSxRH9Go1W6AbwajJ65mbGNrM1Pqc6E4ATXnJwsHmUh+
aWWjJf77VrrlSD4/Yd6m6d00DbmqZotyN/p6HJVfKUZUsG1fwvrbqKaqOk2WoqIqIEnze0pZOC5+
0msc149IZLuHX1GHxZfT5+dV+mDPz5yxgYMxLNQtJNXi827l++THAcPH/Qu6w+defGvh8V2qB9qK
rAAd8B6uHYt7rWJB0bGbfU7tvK+iB/8gwJK5BpaOlhoPJcE4mcIMb4wjzIoPxW84yN6xygPkqwpv
KBos+AK+P7vKfh8eqIZ2Qd249QmCWEM0Vd+ZwifkOxuM5E7ZMXzeEn6zbwBRMm3Icr72YS06/aZ8
qe4t/TVbu8HwyqeRQqiStHt76pR7QY32c6/JdXKbMna3ynPZHJXIqzScbcXY3QdPjGYSIfW0mh0a
cyjxZ0ZTIFoAXhJg7GIYTYbfO3WUxUmJ60x1kLfYBnlYRXQS/ysEgsGMyRFgfbgrzlPtmR/Ofi0M
GIHBBeZyEYUl3HG9pTdPhJYOTxzls+bXSiC4fuEcartGgp/h5jFVP2Q2VHJRffQwrnI2yQrRAv2E
kLywPd6HEx5FKcKiBjC9uTbgYInFAUd9xFYyl7SZTj/+yfjHxvIlLByUmiIMGbx1cybnw2OTr1Qj
WWDWwufTEh7zlYWQmi5fXiiPV7QjdnCu+B1dq12zFKuvwSDUl167IM2w2pKUEdK647b0DLEs1LIK
QNrPJu4Z1xdWh6ye0Ib49MLdetCe2C2A4AXtv/m1VIu+cE3nL8nfKvJZ0nAnTirKbshPXYFHduq7
rc0OeL+YioSFKGymLoGKn0Tr3KCM1nYefYiOT65fGc7ap8H+uD4+WIO17apVeom/tiYzHVGKd02Y
8G3T50IKmE30fx0eZetwgCamUq9FUEpQM5/5PQM291Ks3ugmtSDQWlIFcpQ66tas9jm8WG7O/9dN
EhBIkb3uzYnNje6/GupKuPddSQsx2PxfK4jmSEqlmx8MafALbS7e9yJmhspjTfsFYJXuYmXLXYSA
LXVx4T6ukK4oAwuxEWBaamwkWk1fbnHeexFhO1rFKsO9x0wD2PF/7BJU13HihWiDWqGA4khdFp9O
oiEOsjniLY6xSc70IsMnKYXN3ZHvCA3I6i/7jabBW1R35DnfHBZiSyDiQKk0m3KHw97h4kSJppBd
qRkHR7PU9KwRUvvEZYJZW1SM5atAfrXRzpPypgp9o45RXEbs4PCGZXHF9PoZ6T7AbqhWdorxFBXy
dKPOcciF/6w3eCR34NyXSKRO+Jxut9OF4DI7j1M384HgxXVa18rleQ4NlYrNQ0tCnRED8Ipzf7EM
DFaFp0mnt1GpXZ6hsH3yhGSTDflhjTa2N7vw6r+H2rerJdjA/sIuIeXbhpCIHabnGSKOMdV90maf
02obAn0FvIrXhRrEDPlO3mt2n7i9wzMnAp1xb9AcaeP1HeCIggHKF0Y0sUL35MvuKk6iy+wyArVG
KyVyL5QORthUwULGxssrWC0ZQ7mUgpIH1JH/dQWl3oKiCoH+SonQ7OHylyfK769JGhDMgLBemCqx
R6WpnufNc04rHF1LJuoFxJMvDzkPV41NSV1owpojKVCNboa8WxSfwin2eNwE4x7WBuECLMsWlIAv
WRuhtWlV30I7jG1x0+trAVzY6nL7stwufFrXZw+Up5t4GLOJ1PRDdWWXqnN4P7w/xT9Tw95P9NVY
wk/WTWHNA/DX6/FCCzotfOWoO+Sp/L/hxchC35pXqoBfRtQG1QJcKlmcylw8Aoh9B0twYDPL6h0J
8gu3ejYFhe4MigIm8z8gNa75G/K1JX738tf9GVUODZ9mK/sHUo6azZLaZByjWc2AhZGYGHzUmFXy
APWGcfE1UIjnl50pQP8NcxkNSNy91EMjALfjFQJwi1EjHcpCYDrellLXu5wBh6SKoFKT1dxdUi/J
oCSJCLSB/fKRtUFGmy8Vdw0pJhQzVMiyjBLHBTOepxzz/AMalilcRqdbt+PbKZYTWAbRRAJDGtOc
RtmlptVOcwI6MfT4ecWOe/FnW+ouSa9d12jouY5vq6pBPs3kOxWYMsf8yj91efzlJhwPnwkvCZcO
YoWiFn67H1BqjIZ6tk3J7tKjqERs13M03RcQQbpX9jwSe8su5noUblDAZd8oNcdl4zmyHj4C6od5
/vBjpLlmf67wUepcGrACMHSigt258b7o4WTS5Pfg6xyHSrdgZuftHRE0t9yntycI8gV0YUjsXc2p
AhN9XsCjnEv5zfoImEA1zMmktwe1zjz2Z36XTp4wtNLE/z53CYj4UX4tYqBba0MrNIlXde2nieeY
k8+pwRlWdi4aoyW3dHmAIkYLSKiFp+kWTf1jrT4cH0+vL42kaU0PdmSnF7IUwMDBUjDvOkHCQ2Cj
um9KOMo9JanybdmZ2S90FxkIIOzL+R19U7jIGxkty5nJj100gTxuepEPEhUGCOU6RXEV9hpOQ9G8
RmlQ1Et7xi0UavPmTEFur6CGbBo9QoWbEChHl7gCNKY+Xx4W04qIZXSrzZ3rx8IN01Ocrt/nmQ8w
aedkH5uaGy8a20IZrg9ImWvazAyWQX0jiP+/kJkZpRXUyNBfdF3I/IsJRkzELL9HlhMsFluD7BZ/
YMBSwYs4Imw6JkgjhkOtinjlPV1mEZmr/TmKcpwfuSYbdbaXNdI1RJBsU4DSTZQhafNSm53kRD4o
FJCHmYnAgrgIng+mX5mSEEg8g0wxD6DvlO9AOtVWWbyUDous9PtZl9RR8lrl4r33jpgwSWT7qu3O
PhJS185nFHpgklCH+3MrWGWb8sJutnn4iMsB4xNSD4zt4ICpHYlIKfzVPf4IxClP001Tq9M5pkMM
sgojlYy7WG9I9yOzHEVj6CFWGjA7XrQwgIhyPLr1JPcaHdMuWpmm6WBk0dK5Lisv+jeyjKvcs6FX
N32ctCXXMFNJBDYOoyw0c4KQvnEPLhbu2v2je2yUi3qwnf/Gr0edHYsjaR6sdUjgjsRKd+JfWXs8
aMOpLoDaKuBWBIekSLwAyWt1vt6Tj+N9p9zNHujZh8ckbHNxp6jbYhsfg+di0qgb0+/cs5t42h3B
/QZ1I+QVWvqRMHlLdug/S5nlq4Fk7QUD0X7Z7XCBdxBQKJLaInUrk51sar+ddCM4+A10XBCkYw4r
gFggEsulaGg+T08pVjWCY1WAZ9iyhgv/xKZ4WanTNkZ8mWw4uVgbJcNg34r/ia/L7J2ZSGGl3Dv/
/qz7zp3vNNQLCfhHd2GKxUMefGGq9l+D3F7HARKgYVZp0mcKiOXW8QIlICao6Go6QG6LL2V8QYKo
H9Vzoa55CaXK0klDiXFhJDcHGKu43tMOi63zhWnJZXlo554e641m5Y0/F373armqaGDjelOZMaZY
u91ROv1p+YZcH7BWUSn7IDxYZspuUsQ7/rX6HIW4fqRjPhEtgNY+cmp4K/g6dGdJrPmZpgltuIgn
tJIh2fwFHPS4g/qBIUeUnbbgKZmEWtKjEE/lskpDDKUiCmgMNgd46N0XjUspTStlUKd++bitPLcu
NO+RcIuSi1Xkm1XDnH9ZF9+NMEPCSE5AIoEafftZKFV4pgJtkPpYv7cNkp0oMpT6G9X8XFRdAOW5
uj20IJpvBsUhryi82oXHe/snWaUUA/4e+B6fiBtTO542rniD80OPxZ07x8SHA5yTTM85wxJpzIuo
mdMTGtUqlGOCa0UGMAOaN9pM68mNoES23+oRFUYAaj9BOpend3OmySsFl2e7U1vXVqI+DI1erfgF
6n/mGk7U2O+J40Gj3n92yA4d704KZTlO/gbLarXPzK5Po1LZOkCOQYKh8v9ezTLJp3PO6+LcKm1q
iMLmZysif/PUYv9KJoDB/U6KJTYDjy+zJmlKfg8HEEWeupgNIUMEWdHTCQE3JeieyJAkq+YFGd/2
y8k/tzdwiT9XJKu6Ye8bvA6rOz623gscyxUvcz9jszqEYPiUBtkOqMBQ3NWT4gJsG08BPK6wuGYi
xU4lZC4HXlfgGNXrznYu7isRrL2fbDFTjYvQCBvLC+pSLWNZmmkkOHqBRQo+sB6wvILZZ6XYP1fD
6oWfGSmS93rXXZ06A25R3veTB2Hi+d9FZeW9kp/wp2AvbsAK5NLNZPIQYzFNnSNZ+XU87ZV1zWQw
temyQHoywiGivB8q5LDZsAT6Sw9aqgCnXQOkvnjRP+8sqCmSTbGMf1qZnFxRN/W/1vqOJ+DZ9oER
m/jypqcMRP0Prr07jcAco026Fe1JXX1dJssUSUAVCY45em8saDI7LCf6/G3wo5L9E+IIGYh37ZnM
CIvAaLdd/0egfKi+19lS7VAobQ0/37gjyDEpWLNHvw/8WIUfvz/E4mSjV6ckWw3+vuKs3bmlGlT2
jBDr3VZamgiRSA8k1jw/iTHeFnqFj39GsmAh667M1eWAvb3uLlqH9g6LO3V9FzGpXR+PP970O6Q7
2Kx/p/63S1O64e9isLMumRS6T77f4fpu2roeGFDgqq89tzy1GAOL+2SL0gF3TRQVUiJWMqz2oukT
nR+jeFJ3wsZwQqDtfOjdm3tWtdxc2RJbBqdpmyeo73DulGcVigMH3kQFwoCj2qHPZz3eF37QQFkZ
JvI/Hc2QFhi/Pk3lgQIEqLWDSa40JNlXl7GrTXhMLZVrvqiRmeuLounBJiPauQVCDq863/CXhVfl
umxmt+VQfuzkkd2XmHrVUIg82ja4qZV1XR7jvGxFiT2M+6EmQmJrqqGsk8FOTXCfRz0EeX3Pt2pN
AvZuTnicCSp5lD0ad3pVkEBPeeSeH1RxMumBr7nTdI3BEfW5gWsvA9NmGhMQxISpkPq4T6/gHgWv
aX/1Z5kZLPPd7YtsLrcvbUFaiJhYP/NzCnUrPPREBREMGnSQ2WdhEsyzTACE8qxJC9x6xsWzdnwf
BvmPiKN982rGn9Nn9xK9ZreMf6WmMn66oM6uVnmVMfFDLlvhcXAfKz2hlrU07Jy3JVNCQUSNOFUO
q0TPnWbGrtCMHMZ/XRP1mX3SxAUwOVTT9O0XHPWFROv8pE8/pejrxp0tKQvxuSIa74h7VuKxFDhn
VH/SZmExFNK7siTWqLJJABV5dVSJk1JiBVA6JOS1/FzHu8PO+RIZRcjswvv3pTYkL9CS0i37aM19
fjl5BgjsOc7n7nPndbfvRcUuzrzQNSCkAXV/MzLVGAkfeo6a9hdBFlr8ojAuoEgb3WKRq+foiXnE
Q6Sbz8bkupGzjBWUIuT7ArSrrFa4nYYd13rPgTVzqQ4LwJZnvZzCnaEE9ozmUKeNft4pfBgTnq3t
U+l/N+MFE8h3Q/zK2XMDkrDnJ+sR/Pqzwb4yZ9RmTPk+AhQThVWR8VA4RVh8KOExpuXk5oeU81gs
iqPu8QPc3KFSnZwlRRZqwsetMjFkXR4H+Z1gPvU1mh9kn85+n2GDI4MKgs8uhbx4ct+e2XMcngci
Uee2/eZI0H2xZNMZ7g/90B0Z2OUzvyIZ3/tJks6fi1mZvaMRBTWtiIwaVzITDep9dRWzYQDFkHu/
aNzmFEoaP5BUc/QuCNXmzkErbxvSRwLEY9usq58l9FA/b800KR4u9U9TXqbWIt6sJuPTTRf36T/L
wLAxk0gr4eT/74lToXuwAdCeh9d5wdRlrFzw3+qT7dB033N++r800IZQo0oogFww1FzDjRp5ZmLv
44deqNQfePegKLGmZ0knVBo/RqOV5rHCOTZpXVqjtrX5BKqD3GqUmAkZC2fX6Vy/A+3NbpB7uQl1
mTmontCJMLuycgfAyWKS18t6nBKwrQIpEtyNeWhKOEGE0k3MUGXemaoN6hLRHT++Vbq/grEFU3u7
XQB1tumFJShhbvtIkdzygViwIAy9EPXV/fZsWEWvmJPFXz0WfuM669YwASmeBe1ZVtdOOwxXRMHa
PV8YCSCxEZKfApBGqkbK7M1qVWUWaMerjQ/heln3QMtD9DZBQvFbq9QTglD26HHbt4C+raa+VFFQ
5c2VZ1z1EgkkFcfGNnz7teRe+Q1wCephSY8MKfD78Shdww5csrKqZEbI5WtPB7q9pjSWcXq7O2n7
IMTFYHg9KsMHwr/W6XmLXbJPwcjzIbjaZoFqeIc4gUPEIGd641vyobvfn7BcmB+V8MHXCaTZ6JgI
ZNTKzx6QkkkvuV4qzg6PmkDUxgEFByv2jtI3u9pO4prMEoGEhsB/btjHou62lihd+NNiNjh0yq1T
wG8YARgYzhOJSRK98V4w6101wgpexccLQEHwnEcROlHd2qqHpRxRg6bwF0UyDur4bfyZyZEK+JFD
8PzwLH5nZgj0C0g6wQnebeE6Vi+LZqJs4HKbouiAUvak4knFeAQ2WUE3YK+21Kk7zxiZtjROy0jd
U9LdvuvCKcEctHIqsD5wnYCc5nfM/mKX2DljX8LO8JXt3XwK9Ff1iRhRqaRicGGNiL/FiVGxd8pc
NDungil3P8flBZ6ru60g2PT9krgAgLgL5UYJM2xJ0l8jzjlHJ4LFGP2fwoNE/aRxo459SQiFKzFT
23DzPqfMI6vlMmDl7dKkxqIQYkYHzVe1SI8r5OYS1UcAJY8HtzOCQHGLDPU8yXcbhuIm+Xh9Sn4Z
bvJOKeUzLIdWt6PhAcAnjDQlrBw/z+089M4s3Datp+iwl+31rPuOU9GpS8/385CZ+0qNozRcgRN/
twmCGWL/yopz8Hq4BvBgPeVEsY5KRX0OpXvSSwDCjI/7EUrLCKZszfeC++2M4gL23SPugAOgLdmA
AMwf1fLzBPwcSxVhDsT/9lQXFoK+p3BUOQknW5HnIyG9wQFBV1W/9mtk38dE6s2vBxVxv+h7YNOZ
35v8ciqE2eTFUonSgJaNZutUJf+LTQX4o3L2buRKcYf5sR2dGfEdARg2/Ujrn5nsY3SpefgX5Rzr
1DOPh5I1F35vMrGUrLhRYcRtt+VhUnnXnLclum4pM1wZ1d2RRn0BNX1ZX5RHqdLaQuetI+nyfc2w
OWCmYoebpeQHJDVyd3nyMk65aknHNsXN50oBecb9NZRrxbJqUfG0dFFk4rmsqMquzT+1MHyT61nB
uLSjgfZJJgRyi4gOCt+L81lyqcxatUv86yefmkktxsTkbIediLRiXEy3KjoC57Wmro00/T5zXE0h
O2nZVgUEwbx3wCmZB9RAVA+7VBJ08ef4jHvP9de3IocISu7uXeOdFK8kOopPInRFzSyaqxj5S1qs
o2ibJ0j1E+gJcoXyrmjAMl+UthruUbgVDjAHgG7tu72J7wX60fcdE1Uo8p4fe730pYVhH8SRH3Fe
Dlo2s92V0X9J8PCQos5VdRLHZDpGSK/edMAsVPN4ZTFhC/Uq9YSeQxZ/b2rnCQmYNG6a0WRQ2Osp
Zlg5Zg66g0cN3c3SrGrz8i9R/9HcdTaAQfQ9eGTdHW3mcZ0v/kNKo4sDMOfy32q6bV58suZ1c8xs
yHpt8UGYg4uc8hXzJqpAO/qyZgMDGFMUkqbOGFColJsbPtnLXrYLCkEMTLitPLNyUy9J6aYnHX+T
deSr+EjwZ6QXdPI/FZR+oG+l0NlrYpYYZt+9vV2MT+lfw8OimDC/+d5tDDErEr9CKPvQq/wRr6ei
8tLCMNVSuAbaVZ6C9cpuitJBsmAoUh9n7jTpIgsotn+XEXWfnt1olJIQhzc0tFXjkZkPaE7m2uWu
X2XgddibJvBfHxdkjdsyq7+iT9Pdst4/W/gx7g71LnrM6pVMwdNtBZI71LlT4lNBbHDxRc2jk17v
J0KmFEOvIH914dKnV/siQ9jmGqjMKSy4sLExckxUCGSl8g4uWTluyXD+vqEAqxOGdfFD8z5Q3eAr
MXWpahXtIvbm1HlPRxwsfVS7eGscao0/2jHwDUsFOSixw08P5FV0aw048NELQoDzvUkADH4DpUsJ
2zj7WsNGDtFt8ayIW99lbVpvzsz4Dk69ySiLZ7z4yslgBcMcRTfDZSwE4lMgwYGlGHClZPt22QRC
zK39YtiH6isP6e+I7guWcsiYGff2gPCZBsTw1ylj8aq1z6e6N6kHw306cHB26rVhq+2rI/suecLl
3ehkiJ5BZ2ILw+rssfpGXIkXSuI6KIeU6kdB1AaRoqNn3AQmyNjSyvMYw/QHJnjvBj1zXN7Dldi8
RRUP2gZeCvcwyhQfszIeJ6ujRcqzzPmhVtJrSq7aF2VQ3kgKVbBPdliuOFiOM66ul9W6IdH40rzo
yJMFjdN9tqyznTrPVIGavsFX7cNmch98uzYFd84uT14qVpnpzM6mZQg+KjV8H/AzVQvJcFdPtQQh
wKb4HegiphNI1Xh3q8Da4Nxq8w00QbXA6Qzbhhl8yAu1n++MbTPJQENseB3RvPmKv+P3SRQhXMLI
dGj8g0/5vxTxREzGrFRreJp6fGbVtk9eKD7qpfsE3maV95qdt/75gE3vH0Acw8pvvwGWuGKjX+YZ
VIUaFc2kuIri3mNGE2T6EKw2t4oL4/Hlhbap3FiIshiijQvfXwaKEiZd9PIrO7PGpl/ZEAmTWEGz
goLNAMSgPE8f9BYyZELluxCZzJi5JpANWSzsPdYdjJFtNYmqkX0SxNHtyTGTLzayMe/1BbMNHwYP
LVT4Q4FuP+cKwsgnZIm6/E+wDKeULJ8rFSLhRZe03tX9nbapfn7BPSuUsM0FxHduf3iThebi0sO8
Bo5lP6vl+s2192f9c9f2oeZnhNLj4GDXiC+dQ1/RwPHUc/xBSqDOW/he/DAJRzC05kJT9tfl8iKt
Alrz/WeASAM9cawZbphEP8LqnArkCRAyN6QZ50k5aGJeY3j+RY4rvSB5Dnl4/88P6eAwCfLBmzch
fRDQT5BFzELQGdyqKB3poz991bi20+kCBeqXh491qR9B4HmNXdddYcyWTUI01XMJ3retXvhdKiWc
in/CJ7iJ50FuPTFT96xuDCGA5jy3zrgD3MxX2gOBB7QDqJfK7VHcK7FuTFW4QrWybuxNffvDgf5Q
jx81uemqJIs6pTEWMbVFhQ9P1f6xPmH2S3FP+qNjEcT919eRKViJ2aMgniJfMvm0zqXHgkH5l+07
paq6yWkGzXx9lqVKofxWcbYp1i6Ups9wtcNWJlSubn2VvQLPCr7rvRAFBRxEUFGTqi6d5n80Kokx
3Dd3QD/+dJ/biDwK0qJy/D/3zlXXEu1ABG7HyyjZY6K9OBkz+qTaxUYuBz4DyU5oO5X12BxcAIiG
ubIx4nYhGGOCpD3os5XlK+vAkagfoYTRssfxQ5UfyHq36XAfPnje1kJM37h1O//Q0b5uV2gqXl6b
68Kpug0w+1cxGEV3SzsdMhxqjmWiirEh0c7FsQeSPOTRdDakxnf7r8wSWzDIysencA7/8TuYwd9C
xav6qQE7zCWamw56RkXjH4aN+CqZSY61eiagDSy0ajp6jnpKBMHYiSU68UuSSk+TctCT1Brt58Yt
5QKrqJpKE0eypi6mNQoz1yOrBPIYTw1O91MQG4s5nGfUHVaevjaJMylPVTYXkbRc3Bu40FQW/WPo
uJAlQRR9XqfhR5ueRU+vtPl1FfVeAuMgCrOI2O57PEcx3DvMXupqoIgzXT3gcfsUyCvdouZWTMFD
QtDeVLKAv6X/48tqY8Fk/7TA2HW1pEeDtMyH7HShKdf5qTY1RvCgp1Q0EiSB148wMA==
`pragma protect end_protected
