// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
rwzj8aCVzjf/bcYAYrScq6CGSbMD4qiWRMK97zSxA6w7GftGorIKupwGshgbXvQr
Oq/4+UD9RUDTzE2L8s8NL6/VveWSwI4Oc3n3wntdaAXT76/1YZG8zahbmYZzEwuK
apmpSXnZ0r02YnFqejcN9/GRg4BCZ88NsIGjRVUcxv4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11488)
2yM4Dxs9Xz8eJCjMVxEHIhVeGaqZITopdmin6V7onHmNU4zRQWT5O6B1NraLzGaL
FxzV5WjcGea3L0fJ25o/7TgDRpDqToodIwGz0ouH5RwfZsCVQq0To5HBzjAdKvN1
ZFNBrMswK8RW83sGYWv5Fw2/Rph/CjvCpdOAFc4CakKCD6S5geOZIhcTDbNFhqtY
0nZZBR3o3sKwnupLT0GFcBwCv6Ft074LFNcedGPk+768PefqmTwQiGoqFPIiH/ch
9AV8qiAnz3F51Kr8WkWmUAQgJnPXPDm9L7Pn52cwsD5n6O0jeG5eieQbYtcFOuV/
oCFY7PjpJMBp7dPxAzdInUsuF2xKyWC5jYerYwHU/cmdjbmHkW5/nV2J1Km8/PAw
yfbCNF+fvGoCIAoW0e6Iimds377lJuxQpFSIlc+oGR4JLWpn/NctnoTgAhBGeIp3
FSjaS2XEaKmS9cy3kTfRZVodH8j3o+UN6Yd9ps+ZP/YK0eeD6o9qT8v+PJqgtdME
O/j+DmGzX4K4itTubsB0S5OLqvlon9Lez2hKoBI7U1Sc3WJik7mrelKgtVCAl3EO
/WFbeiRaL91cUCCi56NChrFNkoPQ9LjjHjDiaNkXlF7SSHJ89ntkl8RFDTYL4Qqz
e0TzjE2vhrF4l97R5ncBnbX/F/keeUShe0cuvIo/OCFFOZHRHzv9sXoZXqDN2WYq
eOkIyreeXwEJVyUuT1uBN1/RJEurbJV465pXLxEkacnr8qyTKjjFT0kgScDUvA+M
z1VPgDJFKcwXweGs+OuEh2PtLvaT/eUpoGNRw/pSGVBZljMjrthpXjits2yIe/YE
hypg8XeWdUpZaqSGUPdaRRM+ftqXPu3jjJI5+eZfVTsxeQURleWRYVXH4ryoIzw9
NdaQEUFP9VTH0T40e0ezpmo0vAHldtVGYZn3AAuQZ1C56/ltIGcl0c7JjO3BoW9X
irOKqrRRlUSQ9BX27UKnqma+SGLDjIKVXFcaOSWhSETd1iSjfvsbxjjkxSeWT8bb
7gWVK5Jw7sb2bC5zBJ21tsOXi67+UWGFzdGBnRSlb1W4QJUCbHnLy+lln3NWzgKt
hOsdT1comTWPkSNYCS0Rva0nftmQx5rk1HKvTfjSmVhUGYJlloWJ9QlV/5Rp8KnJ
TW+HvQsuk14A7SGap7vkxV2/KhBEC55SykQmcIOdbped0v1TRK8+7KxYxVVhyg6v
+HCCofXFQt4/vGCzD0ngpLSB7FJpNT1TYJD3UC2DVJ0CmDUG/zqjnrB0Tg9X3QtC
40v0PCA6bu30WwPQ+QTnK1bnE1XTlZGwioOkt8c04oRbR4GrjR7qAR3saLxPtyMZ
qL+rsUEoni/f7Sh/8SLPSulMmJENCZbImBAwJnqa7j44msoue1+ysuQsVTKiNJSB
72kMjURehl5HmZb+8O+VFqr8wishhfoUfZZuz7P+4I11WzZ3Xhy/dP1qw2yajkl+
K2w6SbrDNLWxMZlzPqG2x1mn3CLI3lTBes5qz0GvHL5ZPQrlPcdAJLYdkOX5cy2g
/Bo/tz9/yP3MqfVmnTNniJjy7lLJ+ug68BSeflBVF/uNGMDzxdpxptGk6W87SBC4
mALVcgGpNumXm0juLw3JQt++skrX5zkwqGjieGCkgZHQyhi0kE3OA04DYMPksjT1
qJeTm0cO4CFTESaAckL9LHprC1pHvonPwhDrADqPcYu+/qgmWvoYDG2hhhdBgQxU
4h0J8TPesoHxpzxlPsANiM3S8egfEFGMGrCRBynHeuERQ6RmdA0b0EiY461FwZ6k
GIehp6wcx8FqYW9/7BbDSodeZe+qrAYCvwtS7NzFoM+QMkzGMUDa8/b1PRBTqW2E
9SDlOZaPNkYVr3aOK1yuGrI1yemDq7hAdsHJzhg+hLBTa+8vdj9wvLLrRnxetRk3
UZUMh+KNq8hdhhQtXnAOnZhBehJaRTiix5fS7VS6kCOYiDlsXBw8mrrjncdUesVx
CeLf1quCibBBtfl2ilL07+MJtbUPzJ/o0pC9QSHfmlkF+5XEg89w55Warm8yNigx
D8WcVpfDLj8sXmGf2wNDNzE5/D6PefGJepo1dzcBk4OV8dfWq8khxjmb5wcXKAkp
OGK4dHXqFeAbukBXbYiLpjvsCJmtDrk+cTO4L3mkRKiVYYkH6sMhx7YrvnlP3kAY
BIEWj1PqoR6GTG2wdTxsiPnIoq0TpAgm/yJHAzBCGwKio+cUtatGDDcFmG6BJ4kp
gTchvDF19BUTemH8tKLtTV+dgF7prbxt7JfzsnmXrU5R3o0Zp28+oU55tBanH4LF
kDF+4YOBuh1i+tEVAKNrZIkGroq7TiYBfsTUJeTy6Ge4QlOGVU8VtDmixvLvkzeH
DYBOv05nsBRky2+m0oJK9FF79oVCglk4jWJrTFI7HXubWHWp3JLFHmmHZyP8G79e
YR/0YF4cVqUHe0lMuRhZezMNfR9KZyQyfItU8t/CCcRQHtK7dqrZZqVoOGuaJkak
oq+wQyDeOi7m516AlBf/AtIqVciw6TY74+557X4MBITRmZL22175PaGTzfjyMEsp
oKWrWhz/2hi2JS6RAD/YrYZ++Z06kKibQODeqqpOhah8zSEX41LKzlqLri+7HY5n
A7qouTLqwvIcYbuZrzXVVhNs/bZqbL7tayzr52rL4dL27UdiTtmbmQ4QUMhNQDSp
NvZpvE0vbZ+4bAtbDgWQyPtDXxGLys7JSFne1VcRjzHZxx9mKD1NqqJikXq4uMdU
f06IHDtv489dvrhtMoCUFvF51eIAAWWKh7/U9EfJYHZ5yONlOdyMtoGwo/C8TCrK
U1WZ9JOKPiRyyCJhaDFiAZXHyswO1YT95cbJDFs5cCC7b7Wtk7TzIMaYQINnFsQG
sIeKB/8jTnKvfNZHW0W0tivrVk/dcUnchuXKvCBj0WdMwMB9H9n/OLRvZXbexr9w
so1Fqg8Tvtpmf3pl1zqpcbMd4fJX0fv1DCicjY7ABs8gwCz2KAf7MRwh1dZcndC7
qRx8x4WkgldvNLCCTErQNZYNMnUhDVnMqu/tzp7YPEs9Ix/Ea/rba7JZxq5R20ZA
KBdH4Jv8mvAiUFjMIUhyQ2Lcn2pSdT0f04DyXwlofMTfAGXJDwJ/peJ165L/3RYw
4hH6qsg032C6z72SHTBI9TxQ484m9u2W2LyLPatMeGT4kD2ykoV1F3BtlyXzYSSd
qJc0FSY4gqymg3MITm8+kFcgWTPHxmildEIJzknrOLlUQ3NRActytkct+WepNwMP
uRFJ78X/T8sRkvEqbOxUF9xSKBaEezx/1CLKjl5EMbMaC1vBdz0WRbgotHfnkJwv
QEi6glHFqbvAAXYFVXTj/MssJ81cXMXD793CC2YluaeJxnVo9UrXItG2FrWSquuY
jojtPKZERt4uLdwxfyMWC6FawhGI+frpq8QhoVD+eJzRH56gpvTnNoL5rxTcCak9
KHzkEy7ldKMiHce8nMQzbC+2NATheFz5PqUpBnbz7tu4+aBY/vsYib/LsSdRaHo/
f6YP051NPC6yyai9uQ1hjy3zGFWGImGSajHgJ2z/kfyOt/xmeW8P8eGNj/b6qr4+
a5unJSrU/OBU7pG4CxwNLHdbNcvpjnY2czL6X+BRV4ZFgbYAVoCE7XMExn9NObwt
gBPa5GdnakeYAjaFcb47d1ln04lXPwpjSPQRCbwFH/RBKI7QED/PGQr8Cv6W4B0F
ZhlvsTFUiN80YCqAYxC98gjgSziNzA8TkmhrHLrY9O1Bd8da8+Jx0L+Ks/QoPsPM
oHM9YDoGH4LwtwnqvJa6JR352EvO1ZbLc73nxpcjt07Vap4KN7abFH3KBe8C6HZh
wCcEaClkr4jTpzsG+xf6G7LeY0ceogIeeahgFAazrZnBzLpHHig5zLMVprGIFevt
9t05K/q3mA4aAGs0mpCAX2QOk89CVYFvO3kjY2LwS3ojw0ADLiJL+5zUdwc/XMUZ
Ko944wBdyfFSK8Utcp05+NOm9ng4067AKwOrRJ27coNO/9Ov5tKQYtcYLGsyXL8e
01Z9HXsV2Qij9/KwZrNxOTRlG3+8M+nUxAE232lnmafYtHCRlQ8sf8pYhDsrUFK+
1+4sc9dRYZZDV/EohCeFD1Ebfk57F1ZeIqzwwsKMHEpw4PsETzRI5zRa/ABA7lnr
oqlgYte3gVjNRrO762j9jlQgJ2V+BrMPL8gPIXmeAVI+NvoCtwjXe4YmlkWazN3j
GoYbp74QXY0MIVQUwK6tfmHzbAp4Eq/ecsE6VjSeRz8Qi8LoR6OldDLRvrwX9QDr
ml4dtbdBtG6yswl5llmBDngWNXUzkq23ks+umob65eFp3F+9FlgajW2aSR0+NN0b
sFwKT4bOtTN39HuSVKktXymy3XkQq66UUnLFOnzA6EERMpiLz8IyVMOaJ3rxn1sx
xWmVfiDAFVHpIXTbKZGyFJTjiPt4zJSz2JFQf3C9R4sX/kIclMk30QLrxTuO6+pE
DgTS8pNG4hJfS/BKs1LPcf3ykWzzhyNAmwWm/U2kjsUiJxYoMFnoom1GHGlpqMNX
5EIeAdAtw97tHs1FrnfF+973Fh+sugXGXgSQgelfpdaoB52VVuR3pPh2D59ayNe2
OxUt77p428gZ9gqnTM1nj2gFnMEoJG5xeZGNbMyfZyRBiZzJMPaSb9/23JqJlRLq
2HTkPCP0+6uVJtGgufuko5A5n0uBNjyIu9zd3FV/cSZ2zM+q2BHZfH0xlu46CfMC
jB3BHE99Zz1ZkJYN9vipwQexGcXtSilCHt5GX3n1D0zgPXWsFkRYN6TonPss2wBF
zLI2slaSpBraXzdtzuTHRzVgqbMSI3XpcO0SUvKxtdvNyoABeMXfs/FBVS6Ec6tr
hownWqUrfNWveu8thYRFSGmZus9kPyMxMr9jy/oQWqt2Rp96k0/NoMYyxeIQOpj3
d4bUwbEFM17izBHYhj2lcDnM3dabGTASYzDOS+6BhhPVm+zVF9SRKxRj+jbTULY3
1IQJIcUfAIWM9qdpyj91vyy5FfoeoAOFSLTFYPn43ommKaYMoOapzArV0EWrbwos
+tMo3IBrwXxu+Ayea1kGHhggguNrxP030/EZPwelUdnwTRz5QVfQpxcVlyMNQ7vK
e/62B7dxPZGeB5le47JFFlkDAWbdFwzmStPJnKrVPvKvXBPYWmaSHS8I7aADiDcK
RkVZIxtjppM1h6wsMxGLCZUvhYVx3hVPjw3POn459ooa9/MIvESfxeu4FWGUdc02
wwG5oHPnY2NGIrVozuJyHt7Deb9jrmDtjHwGZYW7I4k1k4sG57KkW3vty1sECn5V
pz73H+NcRyJBXqkVm8hO7KtLTZdqTYjtPyV1S+v1no5mQrOO6pmIP3cPYZCsUlzQ
Lx7Ryo6zDPvjkeTg0IgUjFNT3LHalIcWK+UW6w8dyeWzQUJjxWppF73F1MQf1Kt+
dcq9XFgA9hESzPUU64JbFs4ZA4eNtRPejv5rAUI6duSexxi1I68vyZz6Lum7WC3Y
WL3WwWNlPIU9Z2ca36nG+xT3y5T9hxPhM2d2K/IddH5ZcQBToqqOe8X7gIs7u1Q7
x7UKoFJ4lPOaZazYU5ap+wee21aFgF74Qt4C/V5mzcH8/62q0GNKgSDOUFdSUHnI
6v3i/4dw8pfqXoC7htQfJkYqAeXJwAJwYsX/QgzsDg3dDEONbi/2zrpK2DvL+5jg
sUg4EvHzj2HieM0oIiOsOYiRpArl5LwmXu37TzDTLa3FKfaFTL7NI0EmwEdZm07M
uAZu8ZB5yUoEEWRKLl6XoFquY6dh4j7bC+SNhymAZ/Aa3FlOYmhiYbDHN87/L2r9
lymKkamJltIVNer8mgEubn/0xNeTREzM+tjSh5990RDyrFRdVxKu6VO/JWa8gcoY
De3ezxDJY5F87XRgyoYrHlxnw9Hh3W1j+fqLNr4N/BKHWNJCROAidjdmKims9vhm
B1Kvy+Vow3Bfd5f6kx154p2igfZCyXtpxsEZrXS5liD9a7Dd84lSvsr8VHyuOGnZ
oEbT0GTRSHF346KrnF811gaVjUPDo3Bo3ceyf+V+i1cyYWLXk2V83UjrWXaNHtqO
iW43g1SAbgc9UAshlQc2ROZFecs2ymK/wTWnLWPuJa10CxeoY2SQeJalRF003IgY
BW9bcvZSyu0dPydFwMKTjwh6zgan4YB6ax+tF54is3DpRDPavT7yI5AZbyrR9j7x
GdBobtdXWJskbeYiZ0Q3ZTVwUmU1DH9q3Kiize5LEZPZ3TEsIHY6ZGP5FrlrStQS
Uvpx5vyDsm5uyc9brxdUFkT1XiAAwGbQilzDuL45RwExm4Yey1i35UqbNshrA6Du
c3E51cLWhPDFmFsIm85iYHC48MeDXtQSvDdcd8MYzHoY3PQR9aKNVM+i9MInWKMq
fziPv/DckOsLYGFE3QY2v4e952J96RGm/pAzaUi9wgNI5OvZmybLIkb5CsHE8x0q
PRcl2JjwbzMAlyr4EzqLLUHuyRSiMjUFol0H7UVYPrXgfNgc+bjS+qAcNCsfNACH
eY0Mq9TBioKZo4O0J39ajDdncEbTnRhvhbn2vGri3VQMK3kqTGI0Vnn+zkKUnSUI
OmnkWSfcC7b6lTNR2Ge04mM0zdropSuC9zPaMTviKk+zXOPAXj+WJ1RuppKyvZS/
llz6qsM/hYCZ0zoA+is1lr2qcO6IlDuTUDvFWaXHHIqdYCGOTTppSdHKQ3e8iXRj
QepNSmDWKW8beKmFH6YzslU6HcuGHfxWw7bnuZ+KSLc9UETus8eLCxOB4oluPhZT
ZDtvaxbQ8ao/6eXGTKOsWzXiQdVr9iEkY1B+qQ7BvpAnh7lHbrxU/e5+ctfEvkwb
FpPzd+HtsPTpLufRQPhw8Y89FqWS2Ri8w1kgbjeWSqXJbNm6Il/PEa7pmu/pHtB6
5XGxG9VZ+gWqQ/n1ilvWf94mLkpnfHFOCDCxJMRgBBdfqqb1zmxlTf4JZnH9zlvQ
SRyAv5zUFigsk5NlWigrNDSKRtONKt08uz0R9kk24jQ5m1bLCF+usjv7xATQFm9n
oc9JUYzwWOQrrBOVc4riHmNafgJRZZRPFFLtJ5XOf9Nd44MHu2lO7dGYnVBhhLBd
AVyryW5JmxfR9LhM/je2mMc3eoFacReIlmq4djtV9+RYAFUJ2iramB+7ymhl1s22
aBgDg5CqhwVid2v8XEgwxiJ19ju5y6smbMIhv5ZebNK3n/978+DNb2UA4ONLKgql
BImVTExPh+c1Gqgq12dKyrMm6qqMQFom/7Ghw+eNEXnW7LXSPPJ/QvthVeJ6rNWP
a68/Lo1OL8LHKttlCJNxga+4oGVezvf+VKWcEvl+unG6Jo03tVNqtVE8qn8wKvtq
MjsRf/AzNncm7f61gXfYJP7NboN8ql0ougZf5WYeRQNSAPq3jsoAtDho4aZ+7k9I
SedoFSPGR31Lfkj8XPmbtWfvlzVYisMuZUXTQ71t/gUg90EqQsVsZiEWFpEBkf8i
wfpf3CyKJKwaLlEf36o+ktZWF7TNhK4HkvNEBIkocF4BRnisBzu1rgU/mGkF9QA6
Ky9Uwt9dgDKmC+4lXSTWLKYx1UjZMqyb5cxPkhZifZbahXg4JfLqMYrWVEnaTV+j
AfByggeGpKhnppiFTMyYMtS/6eN1x01nGNQlOPljr0ZZCZhgjG/xQgawzAP4MoDQ
c17M2dR+KMaycLfyrYzITWYzcWLwn2i24BgWBduAA02CAcmDtxqHXqLhJXZPDd+c
UiTkj+kxYQ+4ftsVzxW1vFE73A52/R0Qi6oGhvmK+/nanWmBaYUl0Gz5PEsrtmss
m8OkvkrBrhwZFhrtzejKPJpi4c1yXX47fdmP4IINOrA4spQVC5FcH2r6GWp4ILCS
Fb1lDdndSCf39c1CUZYKQK8doXqC1wNNV9C+e2tsTqtzc41/ck8F6Lf5735xy2qR
/gO06XnN9g1h4WRkwxQg4CMSgz82/wttSlNOWilFbYdD1MQ4dM8UqBtqAsfhxVpq
0GeppRMYh06l3DGnV7ZhWH1I1N3kl7nEVYxMrzzZJUK5lazn9l7+YJ1k5iZNlRf0
RgimtDfFubwOhGhw51+epcPjFIBerd/apqtQqVsJAe+5q4/7BrHvg1YwzAzq4cX7
NFXjesxeVCjpo2zIHbDoxJpTTYEzWHVAnbGWp8M6PoYZhMTaSht5eNLw43DBOFx6
9gl05p3B4h+MjVc+nudDFlWrrE2eLZ5Ba+JhLpDBhz6fK1xKdO3kVRK1EdphtF1z
a6iBMQc2kQJz9pLgHU19f3R2OSWOSawok8aQBfwcrWyRc6fUKy2SFGn07H4Mctqy
Cqcd+NU5HGPeKQ+VBt93O9YGlccgEN8TphDQDpSNsqDffVAXoXnRcdIAh82exvAN
3ywXagUc3YTH4UfdlUnVS5BS4UhnxuixtQvJ0CvPywxgkzDU6xr1TQJ5GjGpTZOW
7U42KbNyryOrLKDtUEXjO4zPhWKQRCGWXibs974l4yRWVFG514OdzoDQwC5gA6tJ
WgYSn4uivGQYSu6xGF3ly9uSggHyXnBRdtWM2tqTjotac+RefDtCLQKQFJ61UsSC
0lko7pFfJ2zWw6W6tajUgvsafCWy3jU13qIY1stfwzAPSfQ9t968Wb3EaSH2v51B
HGf00Z0HjxzWiICkNNLcws4NgMswl5QuURFc1OsGWqBQqfcz0zUEPXiWmqn+vcBC
+XMhOvu8tKyjL25Y/mo5Xuur6vSOryOx1f4Qa97708VUXApk6kYJ2ivcPgaTr3CO
cuOOJPFmaaeLsasxEejruFmfCdalLT49Lt5TN8B8M44JSlbtI8vcWNj3AFC15t87
p6zEPSbM14oFGFFpYyE1j4z8NgGBIv9ySGVeccnhUR46ewTyqVIh8DHujqFcCCzV
OKyo8X12SZicxbOLjutkP1dmmQ3p6+TNoqE2HdPhob2C0Nr9hSaQqcuzCWaGU5hu
BNZPmLC4I7TgBs2cnpkncdd52nbLWZgOr/HI2pziS6lkmsCz2qhZ+HoaoSjI++wu
cXojlYBUseeeYsCO9sYleAPqE3ZY1kABIyo2keDFbz63ofYEYEKICWLJNc+dOAVC
SzrD4/duCiHTtG3vE1apLccwhwDBzdZxbjOk3vtijJzgWuEQL0xwhiI4Zndmb/M9
9UOdef0NgQYqH7yK9GMyYUcPe93JSflyKO8JNY+0rdQFCSBohCpcwywWZrM+3fBV
y/z+kshT8gjrwJ/e4jCxGarNM4f+THywFR6WN+IWAvqKAxY2WuHIMK6BH863Xldb
O2+0aFpBXmlEfX621F6vakkBTU2r6b9QTAItzvoGRwL50zOdRxG910k2fWY7a4Wp
WgzlfVnOYoH0oOWG35MRcmtbpj/exPP5ckR5syaCGCREARM3Rkgj5lYb4Fhs2wcE
gEOg+/FdErxaqcvnENiT+3NEaupVbRLhqleYxBRdLoIiB8ZMSFZybV8mcchx/x7A
qN8hibRZl89mPdpjKExKxMmv7BfxcAUSUQmN1vnRzxRK60/BK7AoFpIYzpBPduEb
NgPfGxbp4unICLjOmWfa7R2RWOAgR31uZi4+AE+2+LXFhgzyOx/E5tZIKkPjqKsX
uHN8n8DkOYXf8c7/4zddyDNOaBUVmVdcD2+HLwPZxuCv/6gpNbPm50d2wcbXTW59
mpRIRMWiFtTkoTYpuUecucY56PWkxbIaAJYL4Sz9UlEtEOFpxIKuEFeYfFYgJSZ8
FBNXs5OFf8GzxhtlNf1fZk4bKh+97mgBf8NkI0eO2pwT9ydYVZcRoO1dRKdVBKGF
PAFsKxgIESUhr/h/mc9XaD9kGH5WUshh/okJ11vJxFhQND1DJPM1JpnFXAs5QFK9
HWI2EjATalMR+jnSdpGeQtdbRF3E390K/aTvgtJtDkKqpzem6I5PSt7b9WNrPlRU
npvdaruhwi3+m8DJy91Dkc4zwm4xwzg76jDsht43OSvVVZSTa3Q3h6iaClW1FmAz
QNdLl8JP63+pXY2OtRCKGhIpqaKk9M+YynvE85gg0DsKzgOFIqjCGbZShQYVGvlk
fqE++6AhNtMjjMlvXEz/c7A5Msa+fTHKsBleBIDFi2CAGFNU272scRjeaP0IC1w2
T5FWbUu9fINNOg1xKoWzYaqIZtykJR66MGgmnb9/0UgwCBsKBFCBhnr319FW5Tf0
FxxX6oI0AKmAwsDuGvv4fwGyJ3MsIwp1gzbM95phTYUiP6/heahbVT3IvxQENP1E
/ZvU+BFu29cAW4nul7oj1KWrlmGsJ97M9rwhYBwfxgBiUcaIXZ2nCkWwH0M5lw/X
ivf8uK//zezGG6cumLclL0tEwEXxyI3a3zBbF9h/ss7xzfRWu0rKt8yafelh+yl7
9CLX/0smR++iFzKzprr8em2hMEZl4LEwtid552Vj6s64kMBvlwxMp47JgGDe2m02
T5yC3B4PvGRIc1I0M9EojjjFHae2b5xtWfScxRR42VJMuyCk/Xg1DAs6BJ00Sqfh
edvb2ql16jxjRvZmGjVr3F2+uFTjrtPSpjeSh9pPIEWtV2oXSyLrbHoBfjbyMZqn
v8vXk0AOzvq9wLxTyMkx39yUbyzyMAh9Ov3GUfVLOW02RVCTNIfBQYpE6shdXnyO
5HABlRugcMiuS2Ng2j0fMrtJnocFPVRs9OVClQa0qxKl4vmSVSfU03R5tHG1PLg7
DJZdc4iO9FbSfkZf2IeOwi6mYHkgF6VMVThc9o6QEOxxPChSs1A9qQEBMbyC/FEA
HdY+zhchW0dPg1WKeiRLG9vy1W97znvAI/zcTrlyHUKD21LrqaoIYXH0Ci03hdF1
qf8sY71JU9ewt0an2TTTAhXrTNGydUzpIA5j5JB8kkR6CtcZwoFzrN67R46YVBUa
EHbErTFTKUzSb+k2eyFlZ9QUTjPN+PD/3Y7TINvQFaXbHpgWFv2TNS2ca0mLKZhO
rMg1tQl+GcnCtR3pin6W/jXVi8VbtcyLUbE42vZgOe2F3dqIEEX//kEFnoGEXyBC
5+X1b5CFoVgULyDms2BK4HvPpmr6/ySMh9GMmyNaBgc8373Z1a5KMTGK5um0F+PW
6h5HOoEUfnF+LKqHSnhMHxtBVtI6MtrPLV7Kk+bhaQqrwFuTV2j0K+qmeMvkIgZS
/9m7XIxkKYNI3zXXT8v+34k/x2Ts70qvL2j9lXOklR7SEkyRJVO/E87fXbsbzXi1
zu9gDvkcDwo40RajbxyPLRd2i6tLZsGqnuG/8eaPh9kw0op3nVAV0OvXQBJ+QijB
bXM4dOitIrNIfIQzKfXXFGSoU+q9Fc5LGW7JNtG78EB34dkqnnO0sXBqfU9dj4GV
5Kq0HZ6Uyg09I/iQggB0rPKXWLfti7HQsOGi7TH/MjI3XeaMK9dR5F4WmzVJ57w0
rdekAlqSpKrwhgVJ+9FUzYNrtUmV8g7Owm4Y0TvHe+v4jByFG81/qq1+Q4QQ/Vks
ZMUqMCs9R1gLE9h7etiY5cjoOhQT0KQYVhrCpUwecCL5wCRBmaUaGZrxEGPiqI++
Vp7Bf6wa2b76x75cYlU1DTV/omG0XKkhECtMYsF4bHgF3yOswApGYKhwpP3YA6XV
9S0ZpYDWzL/L6385yzdQQMElHfyRqoxl7CNk1vWn85O3YIW5HTWm0UfDkFtawQpv
dkHlLoKtl9AemiKtOPyGya/EUW04d8V4V4Y1kGZCrcKt38iEnTY46lAs1lWZgEcO
Dwt+oVKurVW3v8X8jzXMBxoVaXSj/G3dN/j1dod7P3ocsQDsxrqpsyy4z2mAZSuE
+zD4DePQA/fpjgfvlqNTigGqZaCj7DdDPogqDJNySoiwkCMASd/mzsuNITAD/fzR
VRNB3olA6p10AYcPKmOLu6IObphbaSM5mRm0Yge7oDZGGP2Kf9381oQNK6LIEPfd
QDBBED7sGvKRls8wpsV3AplUJaOm6xiNnPzqy2iAdyDsXLiSWnIo4ux14h40X/Qj
ugt/RRBKT7UFMjX+zsm2lHF5JKi9QgCwjwb1CjnIlOQ0QfhFg6pDRluI9WUyQ4kF
H/fscHrdbcsr1tnLCfyB7j0y0KfokjJ+ZnXte5g/e5cdjWb4pnXhHMxcnvNdh+Xz
KOHhWTFmoS6BRupxTiK0+wJaIiroc3omsaIflccF1VCkNzWtU5t6fX80L7TWeuvx
U3wAgIIiQNPfmqepRJUgtsjH4wikzi/GLfzw5VY+3PNdGLv3AJikVj/pgmU8r3lX
SBBL1eTOmqUIFBy8qbT6JvPl8s7NPsb7AjkhnUTULLBV8gxlwTy75nlKigZ3jhan
XlC61wd6piyqnCdrZXvrZ+JqM2gMsY8wdr/w2IE9K+mbC0HCYxyfgePXNn87AikA
D7Jr0mPnGTLKjabP0oUdugTv4cwnENSJ0ycQ38tnh+vfsizuhyjOiICT32FhYuIy
k/rnZMx/+e0HPnHswTdQ7YckI9V2Xq5CXQJ0frKkoNm2K2PGSnZ0ZRZXSg5dbMX2
pasa4QiXz7MwRu/YhWL30aDYL+B5H4beptn+6B6XxvT3osu29t5c+4GWaCfAL1TF
tV1tcbDssN3deAxJ+C7w9hFRsvYhkMPxVy11dbwFhVINBpNubXIOzY+it5IffLFp
EUI4v7cE4Nmyh7KRz9c8mOIo3hL0IizMqfuIOEPvfhR27f9DQPVKS3f/LsjP9IZn
BQWQCP8DKM/W14sA/pYe7XkMGgZYatA5g+Bp2ECYphgDwhLbWB47qn+FMYs3IVs+
XIOLXqZJJF/BtKYO3XIB1RBG0sGJuM+aJ5qAryilUR+Zz5mDr8X39ycXlmHg0bh5
ESDQG+DhSgklZgpbJK44EiHIqq2G79DiCdh4Gw5SGoZXjHtPipWTXpj1kW1gzXCp
MyJ/CrJzeb8bzhyc0chLYCXPehA3VLhzqv+iBai+ALAL5ECW5T+HWiVLG+x7nzQH
JeeO+QiOOEILY3UzATgi+2Lp0z9eyNcgmoGhjBUWA1k+OH4sFi2X2BZoX0erSUpg
0HkSfCthyLldI3YnFRc6vforBLpmzNfNH/XrbZP+ckCt5wua0JEVzlB0P6PGXw6S
f6AwoITjF0Ag56Asdn1dIfwIFiQWlWy1vp2IaO/YYLAVE/tZjyrpVhdlH2N1UyYO
d8iIaW518qy6UdyyElxGVPpdTJIUpIxJsNkAVOAptyL1JUZl29Rl3pdgI15Rl3bE
WjHBGhegOvM533WG49KNdl05hdipae8cFjKdoKj6K9+drPELDxfFJWE23LpvAtQm
2wfbYRxF58nDHdwm5MMdnXkx97LNXdlHKRbmxxvXfKslNtd1zcz2mtKuDiuH1we5
r1m2UuOhn30nSXEnrvJruYvGa+17aiTQAaGGw9GJmIW8EC0Vv+JtIGzeanAACL4H
dYyMtLNFmPISjqAM8vGw68BWqTEtrA3Ojtxcikad5UpS0fPHJZU71kw2Z8MpQVO5
suqFGPfWvZn4AIdXGD8+QpZvVG55WGo/f/kYM7nPYaFN8fD3x0uhD3stFPm4z/Iv
N47HF3T9qTYwrkrR2I623aTL9YwP6wF6TyQQoy2FRiEG7U1H+Eu7jlzNo1uk8l6C
iCxUjC7jMJq0ZK5Nx5St+tj6+/UpITuOdWgo3oVg3JGOsOwWrgB6aC756+huoeIy
vL2o5Cp4lyQFVZdUYUzk8Na5FwVMggPRKlK0AbN9ShilQhA0euGFsyRjM8Kj5GYr
7jEozXpEL+zLeAR1zxFf0KJMx90/Aa9DZbGn0Akc5olZmaAc9cTdwIIQhgkEvTli
UbM1wfYpJ2O8pKKSPawlGjAAbd3xgo9qDR2os0wIljH5iXkNES1pZ+lCOHe7D7o4
5Acge8juscH3Y5jK4rIhAn9kl5bdm7fF+/+6C04Lyep+hbx/UkQjnmRBLuJJnjui
SN1tCgnqlIojdbe5tLxLUMWq5wrx/2Qau2XkqNq5imAybX7Eei/8+U+YfkkTBILt
AezsctGAqaRmhFY+VhYnILV9f8WZrHItZ3GfRBEn7BF0Yg3+zdrdysTgcOZtFvBk
OfLupUqnwW1Sr/NWN7QVBM52E/F3xFztIKtOA4lo2kXLsKtzTY48Nb+Sm6OZRExp
nKdRcGyJQMjTfdp3twVvpYgc+evXAo9Y2xETnEPIajTexFRnAXNyR+rW3fca+F31
Oihnz/yBJE9XfCumVYefhJP1UZJtyZvHbf0bPJmBy9SGZd96MA/lpdA4NzAyAIXO
BR9eaYOEBwNdguAzhrwgaLcRLMt125hPitoU/NOx18zp8IqGbzt/XF7SHQIAX0vB
0CixHgJ9jRzvQeGzgkMD9TW7qqg5tsDAXrE5VufI1kFgJNUCkTO3uBwQYMHNPd6E
fZwImOA6lTvCC9ALifFTgk/UxvehFd0V1yAFYNe+805bR5g/3P9n9NXLwCg1ciuR
dNl2bkVweUZgiU+zTrIXLNMgWY0uB3bPdlph63zQsyig1WUEuejdGo0fLin1dFVk
PfRUSgkH7z+A0Xg4YRC6XakreJEcCObZ+gNtO/sL8qGlNtgKB6g5ANOs8qF3RFI+
+g7JyEE9GUE9c1tzr9cp0v09IiQHpbZHuizmT1wOb9xMg57JNmED7uFMx1vfjZ2Z
X7fWcx+gSYO4YIUfNOu6GGmBquXWcfR+36Yn4wAU0Lhil9W66wgyvUjAT+07qdnG
L51/5Z4TtZ/EsbiwK3aFCjJUAnzHlRNMGoFTH+TLSoh8Soe5fdvEaCrbihuuQ3CW
8JPlz6VVNlLHeU3cyYIA6gQ6oUOROQkfaiik+64wgX0nDUwor0Hr2fGIBat6pjR7
U8I0iUVIkd4hLxOqVbD+rDTInVBCLsCK1s8+/G2skfGL8Edjo/Tnj9GV/yKfyXEg
yO6HBHEDdXB8+DmD4NoZkLa0pJVhLT0AbWr+y4QbSkd9vZE0L9Ph8ruKKvYPgDQq
dmudgbM1HOZbaEf1BSEVkLeYs5o9caIOqVtQLOi6qdOPJN9Xna0f7dVqxOa5Lvqa
uCqIE59kqQ9WGBdSBUQHxHGNDuCKhbonkMtbcJKi7mDlMwQvBTMdyh67N2D4Vvef
dxd9Xf7oSEUBt+gkT2kNlHq/1DW01uOSfbyIddN+KEGvbNqIA62hUUC12Th4+8HH
gO+/z4BPlv/yycUHxzF5ARRKbryU5Bq9us/CIvRa7SFEC3sVU7Ngie/EXQbxrJOq
ZwQOH+AkQqcQkN3yMignvO7ZHgrtRQ2rvYr9EA/AJkdjOswvhL3t5OPRuYaPmXUQ
RgIx6dz6vi/wgbxI72QmHZt1mOTaMl5Os5Q/X8h4jD30/X1NngZB/knjXio0N6jt
oIthjWra9UAZ8Qdjfw32+Q==
`pragma protect end_protected
