// (C) 2001-2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
X6eZYirHrDqbKa6O7OuMbrMNKquB5vlBYjiJSjVzA3HI4ixbIjSqGNBdwskqPVOhll7pi5IbD79z
bWEsWc9/p7nVOu9SdD7D6GOLVLTCdfJHiBn2TrzZKc0Kuf6lj+055CxIXXaRBQebvAbybZWeQNUp
XMZWWMnZkBjyI2PqqFgzzb+aLXePg6lDg9L8vy5lkM0dH/qnd4rCYSYHSWvThbH645CVMbDSnkBn
SbRNgg4upsqr+f7CcFt46MtUb/j3YfA9URywnXJeStPbmXDyZvoO89RpvmsYS2Rvhq8D+L59kQiS
va7JFV6Nr1g+e7+irgigWzvcdN+vw+1O35JOTg==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11392)
zDyBOtd/2Xu4L/y+zHVQ6OzqOj3px0dR+jFw6KiewjG+CxRKXtXKxqrBC+wEPSGiyTseAiHJV1y5
MHeLE+Tft5zInpCKNqoTQQDVA4oE26W5q4b46tSkMcWp2O+t265C5i8wstXh4X7pO9JDT5I1sQsr
ttuLsKfl/RF4zwgk5kFUQGWS8xnEWcfM9bGhDdb4OFe0+9lXbwhqPl1gqQ85V6kSOa2zXHl9tFYI
GfAGxAMf9vTFBprevUEEqHSkiz7F35/l66Q9RxPa94eWZSjB6+hn5/6QcVUKH+SHORMpKAUDjhLh
hTtep/IACfcqMi53J6TZZDawALdSeUpTpIAKFxfsS5W55b9/eaInjy/f0Ppbkz9M5uwP4TxtshWy
GdOe1CcJoKf/V47ptYKTJfQ9Cd1TF7ZnBCvQVjArHMexQVCor2di4IcFitXnWoyHiaxoxN1Td+Gh
E1hoQ3Y15oxzlwse52iGQRVPq9a7OOTd14nf2qvWY3ceeX+YJxBm1mmQ27fpJEoE3i+i0bZmeEfD
QpUJEN/Sidz/FSI8dNxWZpLWQQSraGPKQouRCGg1iBggWeH5ZRuXA32X7PZ8iBpFNCCNcNVmPP+V
4HU8Wxaw/CipLPQZ3tVZanhmr+HM+bjl7bsokSUa9nXk6NVW9QDAPtHrnakop4OIz535m4gq0+Hs
d/lT+UtabdMMXP5R7nqbGWxU1xQz2TMYFaFXiu9Xuu+mQkHCnONZlTHIk2P2oKoXcvoCoNDVDl13
hNIm9pAjHErVW0gYGUi9JKakWFHnWtcx3joIBylSvVzqZBhmRcbWATd35yPLSQLCJ6LJEyfsfJSa
TjO4rgSs0UlLvGY4QQ0N13zGv0zi+RNgsH18B9NWl0pOc6aJktuNSNCg+E/xNlY/UxROthkGzZAu
1LJd9fTYV8yT6ZAtCL8CKgQOWxSq9VpopdE+cpd1vjg653GQoiURlyMDI9pchJTKm/uCLHKxgWV5
jOwvuOZyO4Dfw5zMt3Ni78H+tTruHZjJBdzckM+3IKNlLwJv0PSdWAbv9gVwmnzq2k3VhOkgBzue
+MAnGVA54L2if8LDmUd7uBH52w/ab54arUxWCs2NstlQcUZmhGJBQ0JaA2LeapbAfhhu574hx7VD
V/VxE818pLuAr09/N4ollVJ3L/HjyBVne7cqIXenPtndO63xAPUa4g3KPKdQ2cfD5ByBLMg2r9s8
E0HFicDLJZwhgp/Jd9NqU/CNUKGFm3/a/aQGdlRVylVoyu+lWQ+M42DvfL/ayvHwS2yPjiG8gBfj
BJa9odeFnLd668ul93Pi1CbCRxd7xePgY/RSSfomtTQWl7lyQdY3HPBSmnlUSSb0qW0G4uRoQ0AC
YL7X8moytFjhdApjqN9YVvNJIlO4XHnHFd3fXpXlYfqQoIC9WlnGYOz55D/XYsOdVFK3ZW5il/H8
itnbXilSDz4RDXXE1MkxGsvRlcCxqf77Q2LCpTWcb2oRI0Jmnc11ucoS7ivIgy4PauMm0kxFn8Kb
hTC46fm78gzffdnSAJhYjTs9wMLg/CTDAOpHnKGDi2jlr7MFoFZk4AEnLzubCVGlLH/mIuj22bbh
4tlLYbqIKAGqEH47wA+to+czJxKY6oMBvr+0hl53/Er1ee5Zvaz9m49on8JyeCMqn3jX7sFdu3Zr
UqQX9z08KBEcp1TNOpuqsKdR8xmm4ivY4caLNJw0na8G4sSRb08C1HtDlIbl4Son3MkR5YQV+m2N
m1q/fJ9Yao3dSuaixSln5ZzvZcCMNd4RPwGsL94INrvMWeWKojTYeS4wLu/MTjBUfI9a3iKp3MIt
8QFI6AdaLSprkbyBUaiStO0e6GxhpPhl09kxrIhCM6cKk4DgIM5ollaXVSvUMhaio/x+73XPidRP
6dKGFDz+AlltcZlsaRESpFzWwJKFwc19OmhhLQcTyzHb+AnauFw2FjqZGNVgiLSa7xPuCBAQGcmt
iiNvnVcll7PJgeEAxJWJF1G2RX4bLl3koGFtLLxU+10TnLls5Vk8qlExhb/XcB7w2xQeoF7O+J9B
2uQwqtNVnS+udsO1kBmVNcGyxB2CsslMx0dL67Ue6ijDjm9GgS2fGJ/uOkYJr68bvP5uAjtLZgyx
ZGmKQDSihHM15lK6gQJ++66NFsD4rmjWibmzWOXmSKd9LYIWYgv6NckvBB1tMxL8IkyDZkoxkoXA
wZ3rcE8Rd3BxUMcRGPgDyXt72yeUuspYsq+Os2oyiguXZg9Kk7vH1XDIwaTWnUCQCeF1tinhEddr
FkxKwmYoMEfBXZKKcV46dVvkN4w6WUQEREEYvadX7UVoCht//p12gpiYcrmlSPHkx19PuWp1B8j8
LOWMRXFQytGeWjy0Hh9IbnHcb1CAeEG49k6+SV93/4uggDaX0L7AGoi9NxdrwAH3yLhGf9wU7KBL
TuwxW08NsBLvOqGnXaaHd2m21EVEGtk3Ii/2Dm4N3muFJp4YSXPpZiz6B9d0W9G4/S5TcLIJUSjL
9PUaLuOV30+HOzmiRolvF4989iJmCZPnu3fFt7r6tM59lM0RX64C1eBCvXNFw+xaS4qvRe4FSjzg
aKlCnRfQMoKQAoegBr/Rrqr2whSCX7BF1GucHQQDXIpSKnjuMOwyfCbv1gI5UJzvQgYG82d8iUo9
yPilaDjsHoUX5Zj7EcZ7+/ThaHSbxVIv29d5GvVYmED8eMBeTanaP4ecyYpmG8SGRgHnWQOYDEAC
r0hQsyKCZAjnl+d1lRCZIUGl6pCvAsKa8C46DXhhVDm60QX1jmZQ/Q6lFAaZkNw5DqX2bEoeD4BA
1MFlW1urEImtSvVw7gJ8//3fgcLcL6AQhEWcG8GPmi9OYKs0UF+cU8dRFrsj5skrz9Rrnj1G9Qne
VpEQIICl95tCRR2fovADj8Mh8Wv+GnfQTCtBTM0Qup4rODYOvjsL8aV90p7yVEJJgfGiTR+W8ioR
6WcoXiFuWUBdUkjw6c5lCrJyT6Od6J1LUYpjTENRi6p1XJ5FAwD3/L9Ci2PXWkbEuEjZD+E65/Kk
aHp+/6fNbvu1R+2254vnN8pLe6sOpA7+lndGvbhtsYJ8YXi6GfMu1AaWHMMmjJU79XoeTo8TgJXh
evG50Odx83CgjB7QxjOppBoOHqoqN3KfvkF2GM7gr9KHiLUCmP8odWLYfHw7Vt36S/KS+xInrn2u
Hsp9Djio+onFKGwD//q1HKBUCXhuhmmrOXvtN+xwpMeIGzWFCDnprxwdU7lCT9cIEBUDdiBepc/0
HW9AbS2xuc/gIJ4fM9eE3CUMZKYnGg5YjESNp0s02MTjdVMGzUguO+iFJyZP5x77dgPeGwr+5t2f
hz4HRpRSNJablFnAKV14fJ7HcBaBdVnMeACWWKn5CCxpP7zRYK0tUJY10L5ylBpHo75/iS7Gswtg
qObV/jc6TPUtbgMeYbl05dym+3oq5QD+uDWe/R+zPdtkZtwxWJPC8GfZk54pvPbqb/nSUjc1hKr+
WlIekTEGdJaCz4gxqnZaIITqlJvG2fPEedzcVPSaJFgVHeMXe+TWicbBbLv9wVgW8kDZEheWLFLN
6r5p2lJmbmJ948/i7ejpS3LRdYU4pffsERSxnXwZsyYkPFIF7UoerkGby1DIGYjBfVgyh1P7EaZL
lhw63n5XpetfJnWpAu6Bo8pbU7evzTr+LWOeGcphtd00eY9YMKhOw4XFQaxohKDl7iGdxTUze7ue
455AoNCPeMnyvjGMxrS+DZPZA6gKeain/mk86HKHIelz2Y76a6gPOyxin00PXGV32g7l8j10E6/W
Zmxczu/WkRCGzIQM0LMZqhVbPCpMxbkwjRGPQs7FqARUcCafB46kZE20bY+Sb+4rax7p5pYNC8dm
MNaQai1BrfahyHG514p1hvXRG4yEjLAf6nQmTJrOpNUoiO9Td4tQExMiutqm9NEFN7hm5bfH6PDl
04ZvUbjgoTp8ltFjBJkfkKBrIO1+xjQCvnTF55aV5qknYT8fHU+qDi1gLecWpWN4Q7yp4jLON9Ti
XGoeV+Lb8HZo9oUh3wyYP3dWYrbEHPF74cMC7hL0Q3baKBRis39eqM1f8+fpUGyr9TbdAlU5xhpu
tTdJ3hszUcAcLmShomxgv7yHCdu0P45d9UeVwZ7RMyQml1aGaorDWgsHOBC5HLtWLk0ZvRx2YB0C
3P2CzliXqrlsfQco/pidYADFEDGRml9N20kxw8t7XkKOPu/GsESrObroK203sXXPhFbjicqH2X+6
zwbpvHzAk25IqPEIiV831aWHSqjFZzM0qiHCO2ZNmt2HK9GsVbi3sGA0v3wFDyEa/HcOM8t9KxQL
bgFlVhbN1mci67qV+TQuDJ306MWHgWRRSHnHkLvuai9TWqLGLzTNEnwFGzGd5pncUlqnltkYPYa+
qeGkOlXLlzoeHRlf2ozf3Y3THyUn87k9lbre590UX0gh/LxNeIXjLPdg+wnxchEZWHHAQM0Y+h4V
hCPt2orOcDSqKKfuF9K7I3LFnhz06+SjhkuGoGH7hP1CPbxWwdssJ+WMXrfOoiIb8YXf+JpTyUIW
6gaq58jXoAt8fD5cPe31U9LUvIzzrq7tBKNjrlQBbgQW9fSoHpOvnsLc6/6DOXQPANWzKaEq02ij
1Oiw8u9Om+FGBgzfAlQzuZNmAjfuJ3wH+Qs+c6pieKf4Th7IqriDEYMuQXQGuKn2oul2XVC4L5Ka
x8WF0/ppNDwMusLGCsktnPPxb1KUUxSrX7CXNJzuRKb0N6VBUoll4RqkqACZHXsj2hnKCgoNrxki
qMXZZoQQHGMY8awGAsNrPLK4myDcZZsOqcDfSMaPDYkt2lbjmCIF9AthHjEsa1OC1qAXCkDQAz2a
p4ynN0rdSQRAX5W3bLVIFxy9p1XFvY5mYdUMEZ28/czfEWaZJx26fD9vbeE/2iO7clJsSGrHcheo
gOVO1kffQO6yLfVrI4a9ugzUb4yeK3dQWCPNpX8sYIOi9JDZnFMrtY6EG4MdoUhTNVZZtsM5SutG
pb6oszPAgpSV7dL+LAX4m8DEaH/upbMollBxj1+PkAhk4wE0TToeM70bnvMfBnj8vX6L4QG12sPS
fvHHXhvlC5xuSKlxGBdWn+2qXuHeVhF/LGjBailjicSzOIhUoAb8jt1fzcw3CoIW74bY2xqSO+ck
cpzjKxjajoZ6SVxeNIeCoMG7U4OgVKmdBVGpr1YTahk/VlpBeUUJZMSFllPI7X59g+S8qX88AXmc
S5H9r2r0JRK0/Pk7RcVBMhTQR5AOSeV9okQlfKuTYDb95LGQG5l7cL7oBGzFwykzKnSHeBrsyI7O
5oabjke2QD6rcvwKgcmYCvGX2H7oq5YikGKYxci1sLsHpXEnXdNTiCOeyNIDCd/4ey4cCwlHVU96
4gdE80ttVl/h3i+gJ8l8vo7zDFIxdMNRTiu05OvTUkCB3tZIdKDKGD+afNWdGzqKIbM09Ash1hwL
BGFH5Q3Of6ksJoikxVhjGKviqQcrely0fwx4ArXIWyreicbNBZuYI83yVdslkKahTmw0I4aOkwOK
Dwm5vXO3aEIxz4UmVfsOfGUIHW8YI/Ws/0aUoWObS5fEQtJx7yMmvH1rhcWFKcM8rgUgcuGOIXBV
hzXOasERHS8eZebcPM8LFUNHyuXGGKt2hwDw5/fG7HC2nptaCh2uzpr9PUW/5CdkVgLEgZXUu7eg
tWegAWusrdCap73zjB5KfQOn5l1CSiZoi6R+ZTV24AEZtgow/0H18B4WZVw/DwLZvDgy6MVettto
u2hb5DqEgAmbhRyymWS8sjnIiESrjDrlQaKZUzlCoUY+nXjx7AxjuTCDTfQs1zAlM0RthbVH5vpB
w5mRIKnnoVtCMAX7DmOlSBQGihRP+DPf8z8K6t8DRGF1ydOW3Jt7ojEzbfRFcPC9EyQGj6tfG3tq
KEBtFyNhLVWbommqWMd+lV/UbY76ZlsRhqJqFurn8sEZTZCLQ1Ci0Rel0ZREeVk6iWCOt+PXUfVv
n+kD778GFLFQ3ZfEU49gUma0AHt3J3bSfZJazaZyC0hcUrQKEYxUxK0EVB5AGWY+2wKG48YtCJ6S
13O4BH4rLB0KvK/rIf2t10HxGPqIpo/43jgwEltDvlWbSdK/VYJuHXCBx70F+8Ole4MFx9SpqzCL
DoL0fyPabSO5kDO4oYfmgWpLf4pTZHfmcCPdLi999ZPIJHqilnFJoShfvWhS09xCE3dp3lFcLp92
AnI6BrJZTs+Phf+uBnePtmXNs4T6z902ity6QcR3cy1g2pInJiOHOy0LxV55e08WOp7LZKDn1rfn
UtZrXqz62iaifik7pdKlgz47FOqjbxFKYcZwUiISLjfHWk+XrH03dgHIdCrRTDp6rzhfjrqkJuBy
Mq76SfXmT3+n5Yh70ZhVGaXq5+xBCa4HWGCovVtD5zcyW5w6lbbqtywHWHMbGoq+LNZpaNBkyuTF
rmgA3ntz/Unm4ZPChwgEcgezz1Yf02+bFuiG1e7iMS2LvJAGw40Zznlj8P9HDhAbIw4yKMiwyxjg
MGUfScQvZ6q4IQYvs4EikKK+U70PfVFguZRSek9eFfJ8a3I4yzNmUftmhacli600awKzUwwMbicR
Jg1Oyett053ipDr245WmeWmyjMng1O0KuxVOGZrcGcrvfuNUTUcosEW/ufiBE0ZP+TAKLDXSfiWI
gSWbk2Rl81vlyzK6h8WR0nVG8DuX/AUzyj0alj/9SkXNiBxnHn6UhwO8gUstsloBMpaYzjmscd75
xkfFPiFYwm6ttFp1NF/bvYuyUNhXmBr1hnFbFCaxUnjD/IwBAQzgCzMSJ0jL2UQx5jKVT2p2Kxpa
WfUurIztH4TPkJj90gA2LcOTnkZlNJPm3GpjNAYaE0Xppv9jq3KrOqBSrpm5VkTRNOfmal+hzxIz
WyKufAEfOyAVoKGRR+zZa46KV9MiEQM8R2warWsy4KRNkH2Dv2QC0KiV1c6yFEfI14vHMNZ48doW
uLDUhu9fvDEMirbnOzKgEIeJUhoKCY7jOBlCRywOLcYeWOucsz4ytBLYccjIBJ85WWnq2QLwp2fa
B/XdC7Er1V+VRhl5drilOYY3wxOsjCq9Y2ZNBQKCy5qyLsa0aYCvgaV2fnntf80ULHwJedD+rT5R
UX2pYW9lmVZ6g5Y4SRiV1+iXCPctwiBP0vUa3G/httgVshscgWTtCor8yUgLo3fLX2lTpcHgvqFi
YGvpcsvk99AoMDhmpscq5h0WNpDkRnFideKs4zjOVh3qEXjXMHuIoDPJ9pe9ZZcryxuTUJwKq35v
frEzLtaeGkGaNBoL/um0dSYXd5eYq67wYPx3IUx+0JGxbQEOgH0EBsUiWqJ4uppkaMspDyIJB6S0
3lguRKkbpKKLShZH6MNcLcKOqDze20ipCIjM9Cn9yq1Jc8d80tOmVkXSiTay7XwLlLXQ/r5A3OSm
UEpt0PC5KBF0sK8Dwt0bry9VFzcRxMafNwwYjKCjeCZWHWxU7QoUYfl9fy2QeEvNsAKC9gxR5qgC
ZU7xAZct5pEp0HnuxcZEi7DHkyAPzF9RO6j3VVMhO50ueKuohYhCiSH2P37uIYjEnqMprgBFXjSq
T2KN92lSxS1aIm1VZtKt+ee4+ZK7PrTiNHbyGRc5oleAhIoiWeKplacp3XDyWP7pXaEZgdYo6AYZ
5egzrYxBlFd8NoZOtJAGA0ZA1xYWo1gN9Z7iU5nG7XB4S2y3AXZBxZP9csI9s1896wCSd0rMfZUr
loGMJk2HnF7sWag1LldlLiQ28uzJlEoRjt9NeIWVEM0IppawcmDXdX6ZZUYSTbrfajdI56JvAR1c
gAl/9Zelqeeq/HCr5+6Cczsw+74RbME/DAP2E4J6mgnPnpDbuEdx9npw3Y+v2KFHITlieGSv7gJa
yd0LFtqNjSnemzAw0SUOpkgahLWtnrypVau07C1g36oaCp3mzROorbaN8KJBSJnzB7ipGKObyLtd
ehAWhY6GkcgMmIuIxoqOggaIwIehWws5kA0io1u+k4+4Kt5k8Zt+FizTz50q9BA4VscWu+uxA9RN
fAWWNaqkuQHevBAbniZd2q1Ut/TTUHoeq3bWqn5gPIrGmE59U/IDZ4EtVl5L56JoVVfiFc9AR/Zt
9l8Yx0yfhoju4auNtcVESgn21lwCr9gNQ978K/xTEchNezunYpinxg94oDR930fpYorLZbjASet+
tAXZ3om/cGHuvyjNKxvo1xTBbb0As4zgTX9GP0qDMPx+bBlKjLjOwE5dTLf8a9f3d71byd61Vgv8
9GLyHdL4ChR/e0lTV5ZOSR1WWm3ZTFwIcniubpRcyukaLY71zaTcq19q6BmJ4otJ9iELBRSnFqzv
0KJts+7FeKPFICWQpQ2TEq1+DoD962fOMAslJsbh8fqTrQP2NpEsn8CUdl63tqXWsz6CTarwQHZG
PDDPXy9GRrbsfRQd1jU+bQKhLOZhVcqXamJx986hqRFbKazqNqja6g+9c/LR1b7UiOSi1FXKsfYw
P/C8FIcvV3sX5do9IkGmZOomjLZXltuaPJzWb3zbhekiJYV97cPQbuJzyPr/vKgjWtV3xgh0IZxN
cQ6b9WNAeHnj9dNSJb1Factb7M2nSk2jAMOPoYPORY/YCj9gs/RLQsK3x3vkZ2RcRhV02eHUckqv
cEPAcsRDyuauro9DwCb1ooHPGH1chYr0SA4Oaqg5LZKSI5ZURmjRbIUZ7aOFlVFFl3+8wJUvup0v
1exi4QbAiesykh3stvd5989Djp7mM3S4g5bMdtEY9MTkgKSfRqsCiAB3vR3FWyU7+u5J+INdxRDF
zI7d1wOebUcGar6j9XLc6ulUltDY3/CgY5BnxPwc+ABgMkkLUgVb7H66AtCUKdiV9swr8JDRqK+K
TkYYIsgDstvUBmgP2RRtx+RdmDqj7Qngq4kbMpiMAzQS1UeKNeGMg0nFW54P7okf7jafDvU6eNsF
SGuITBBqVvM03PzVT+DreOI5Nl/Aq6WuEG1eyMEf4+baqb2s2U+k67tISI6s/rsFEPOXZMjryHVy
q9Bx2eqyPOUqWNSfflrx/1wTiZN9HTlPeQtiFB+YguRuB0KtwSfIOSCeRuW9m+mibvrBXqM2+ZOE
pDa3wEKOH6Us57W0+znvOfwDOzrSgh/5qzP/jDJcy/NPfHjHwJ0YPCeekNSk+fBG7dg4WWGKdKRS
Wi2y9Q9a70bfxzHFqxJ1C4TDgW3Y6pY/2rXK5lc+J7GtrRd+g8rP4Jdsis/e3mezQuTqDYzvex8y
x10YLBM0FsaNJIq/zDJBD/stGgd5h/UkmBZGDORXW8mNcc+eNUG7h1SpE+DYZefCLk1JgJ8WIAi9
/icZW7Lw5jjCQnE7e2xx4KEBQMwwWldjWV6WcgGwMbuu4SBz5y0XOR5uB1Z5d1oTjw3UNdLehy5P
B+lqfUQGO6mJbhlp9XII55XDCSSEQtNz88Mc+0/gUasEYwC6EXQDR35r47XH5PjIsRKcNh+68K0I
tg0ESZWQ9i24utFs7MqszyM4O+6aYE9OYRjAailPZEJCqQuvklfBsJnhSsPHDOVRFWdP5jcFqwpl
wZtsElQLYbem6Q/H/frOtatTpbQI2kDdNZ93SZ8qHCQwwt60Po8qmGni69GaasWSVaUUfJC/J8PR
mQ9VFJsYQnP2g2ZCZqtyu7+xzKTzjesECwIee4Tfjb8SUus4OvL+fg8WjnKUWXC1f9COWtkrXsCc
VEYvXziosII1DqYqtAroQMgxCOpvk4KQ4k1nR/Rn8024J4LAHx362dnwPTddhtylFCPv1fKGx5qz
Od9nwESY7TyFTI67tfWsTyVtTN8BcVb+XnI4ve945TeT77cz2seCkDIBe7KzXuj5aidmJbQgbUPK
wJjBV+VnRrt4LdbSabNEEJGvtNluTM30x2yWuJD8anBBTZl0JMzwO3aaUdXVtxhlRufNsCpFjtPC
h9xTwHXXCNeObdDyM7BZ5V5l+tsfe42KO6Ux6vCQejKm3qkmJDT2InCp8Yk0UhK2JN+v1mSGhOJM
dHEblwP5DkPfpzg8GKFQLpSsIl8mTNqJrIaGNoevfQmsUfoHcpUZJcLZS3FLTe4tM56q7xzv2BpL
OKlEG75/l/ywj70nIMFfhh59LAYfJirR2WW94chi6AwRe+arG9riymLEKBRgfog3uW2NL/Q5jymx
BVeEs43d3QvUZKTALZYaJE5Xkk2R7E25VA1hd4wJKwj4PG/NDWxzwgDdtpN15zm+uYUh5rgJQCx1
hwAUA9lqcuICyeoN4D6sDelOAXHbo9gXmbr1f8O3g9sl9QD6Ej7m8OZJQnfJltVojZlnPbiKhHf0
5ilYjPcGNaYLZzX04PlP5+i/2hQ0abMFon0yqm88UjW4R5lX8EuaC6bmIqXjgrlGs7fcv/9jMroi
xAWn598vOUEjPmiFZ529q5x+4AgbbeCfPdboYSaGwMb2mh8mlO550NP9HPsYXBqnh2+ruXkAuUf8
jpbqwvnt/zyEyJCNKTiGEmNM6ZAckCIko5iu5yzz5PhN7R4529kX25Qwdw9TjJJHov2aqKmx/YKf
heoSMNh94svB2nC1G5v3dadz25Tgw2JTesb5EGmSvw2iuo1MxOVqLS7zgbi2HHai8ayFZxh/cwt0
IupQBpVF9s7dDfGtlbwW8aRuSzGXe/xx2A37bxKCfjy3iDHhRUipTkDxMBnXLyEE3yY0mXCQZAaj
eHMA5xkl1fsLPAidpO+ACvHOvR1Wsu1ASBSB7xNaVNoOZBULrRhaaUSCFeyXWgVHZ9V1g+1xDfpb
TvrelRccde3UgElqfV2Z3cMfHpjwuYNiG7XbPSYywHmRf9okxOzF6vx/6x6lQkiP9PZjncGyiopb
ClSyD0Lv8w6HcJopcDLcosBUYrojtq1C4knbPktjKlmUXu0usIiOi8dkgTPtlN221MBGkq6wR7vN
yUihF30gyVhzQQkzPfzL8NHyfQ9GGKxaREbjht3ktO6lfIlyRvzPpVu4ybkAwJEW30YgTvaV6wng
G0YNKC2IE+m+Tj/HU82sD96/MYxgm08qkEOosZMfL9Jum1bt2viGMi2K0EAMP3C5evzUOfSqGfIF
+06MulvsfyyzdfNXhsFAlTN/937NCINEKZS7Nk8cHch269+QGzd8GkW0m+Z2jll+k/t5awNMggwQ
8bGryv4+qIcTogKShBy2SVWulYBnPTHrH2ru49U1gJrmU3P8eQnAr/y3FLUEaVbc8m5UKSAxUOuU
i0j1xbFZdv+1uXU+wQAzsvMHue2AneqIyULJVmdVYbO7qJgvFFrkqD7OZcV9FXyq2V1qyLQTf/gK
IQhAADnQBqFgDeol2jckFq/Q5EjRG81vLK4Wl2AhOjQsTPdcn/x+9hUznouD0nAfE4qPm+ltYU0K
YXKF90izPhgxpB9vEt7orJhTYsrViPav77mBPmSfdEU/4fSB+G4IQ+HjDwDHuf85WIn4Sc7yVUiJ
C++Kn5Cp0FSjCLsGH6FvCAF9PiiIowrQ6PiMisgouQuSocEG7DVQvq9nbcbkUQicQOab/1wtVf2i
Mm2bTgKcOAA2dS9P8mkeiuM3QllXh8T7524U99aUZ0iro5Im9gs35ydyqj2IgaHL3m4YhxJL+lij
SVGq5J98cvCyLsMLdESzM2cASWTC9xr6AD8k7DaMu2n6bwLMBAaoCLbrmNbCm7uK6fXo7AAcjD3z
7GU5fmVa6i6EmVmogW08JjUwWRByS7Zd3hxq4zbMC7pDWVlx7LZJvWB0bmLqxezi3TMfjNpUeAWj
F3a3AAtYsinmnn9wTl8el7V9QIOugI41jLO7WZdKx+v8PbOv1sLa5ENLGdRrPrUzE+OuuFbbp+Z1
LtpPUU8be348rPuMOcGhqGRZAPHbcAvZ6CZkTmYvIGO+HkMgJdEXvF0li7buowHn2eNjbjn3heOL
VN1gQM4vlPmSBn6DjH24uk2yNCPARcKl0DbpRh3r+dmq6JVNajpbnrWdyeJVcNiPuX1w2Ufbpp9L
E13L0j74SvVaAsYf4mKo1C7DA4GN1hqVQpzidKLnvnf/zsuAi5dZqt1BlueETl47+ncB1S162OnN
nbSFZih5SAXAD11Q+iOvrrUOYJi4UjpTlDwTxrQbcu7X0Q9ELvkL2cmc0F9fXVfrYXEaqOVx1KBH
B6gsh4cmleN4B5nEzkX9uHo5T7xWSUd0BWmcsDoQlvp8r0JQDTUPhHpRg/6FxLbWlwc7NXnVcTi3
pTo9944frgB+UQCI8ok0w/CGYVSsifDvfCe7PYlSI94ifnPMXchkX/J72do2lKmdM3rzH1KZIEj9
MQS3zoJ6Sh2FzgsNu4jjxJq0e9TZU+0Dz8owErblSWIM6t54f2HPRqGjJfWFoSfr+iBptqPgVIde
IzvFb72b0+3M93heHk1J3zBr5izXHwKlFuT1M7/+xDE8GZO7FOXpWLpMGzhsU+loGy5vMnnPhsLz
yYGxNzHCGRMgix8pxdU32g2Z8ydRuRFEtTUg8owEWbKLLMdmgpgP13yZWP2gDr5Jtlcrm99ZHtdF
GBrMPT/4chsBIwsQhfA9EK/I/VE1ChsjjudlL3PTPEcsyelv0A/TO5uPUaqL7L1+HSxD3dAy7+8y
2XqBv7ZvMlmN9WotRUJYSHXXTXybMOdxL3bA8bI9OEVzIYGbhdgfLs5ng5hyuZAcj7sQMYitHL2W
exjkhXKJl1oEEOm8dCjRBc0YMD6acSmJbbTS44Spgq1vgu0uzVuaigE+FCABZJ91YwLKSWIs9GxE
v1NdQ7+i1HEGhDgtN10a9LJ7OJRA5E+AAZDJIVmYk4W6CtRM33QI89KoegQUCHWrF5/o2vg0Axfo
7+D6hCoXCBno51y81rG/BpkXTyFFxW/M3nrOcCtXY6QnsBTAfGgZwsqQkAnLjprA9urYRc+O3w8P
vBLt20p6EAFL4O3R18Xja8L7+fkpUZdYlhujr2xtrPuBySUHFFix9aHGIvuX+TuyAfCsdInSufUA
yxEEVXHa4uyEklLe57tRvN8XWoDq7CmsCUAiocNDQIlpHU7EZqrXxm7zo92A0uTValEBopMb9KYu
NLvZ8Bbo0B/jXVbpJEyFmh9zPdm5N+S+vdLx9KsgUbZuFCu0R94D/y/Qw/XfUsaLSrQHSXu9jDHi
T2pOkriCTByNgpRP+ju2KP0YMSTzdtgyLXZsInzeb7/WIfX1J0rHdAuEv+21plESB0iBIRwpGaVX
Luk0EWX7rRrqoZPRy2LZaq4q8VC/qBNuOyx72LRCH9zEIJTGNXnpry6+rYasQ3pE2HAS65IzWxOR
xO4lSddo2S5GxuAsqYRuVY8Ar/uvnzjJDQo14EAgvPRet8qifzj5HvC14Nmb0vMd4tfZnfnV2w4V
TmOJiwtpqibC18X4s+hHvensq7HrHiTURt9oVUum9ep7m319oplyoo9sRFO9eaMxXGkJH+XSLRdX
3RnqoGVIFPUY8I9Xk0aJrDRaXS0PG99HlpacgPBGaONKZbAkSwCRRL/w4kIty5uhALJEonxXt1yT
hDFzHZIXLl5XxR65ZrudqsfodlBHLuv5td5zcSPTK3RIFsxqNiAfmlcqj6NBVAEBbXEta4cjW4gA
uOj2nOWCZdActx/DdNTZZjWeVSQ3CFRvpMe1OsuWXeUwh34RALdplAp9hi+A4/wWrArcc3fWK71n
8izmWPxBoyzgLxL2s8mzGryrwUVeJMzpGI2FqfEb0Q0sewHloiSgdoNt6Hk29ZUdOVsEzc2w3ApQ
UHC+qyodX7j9vZVaPQ/8fwwGMtCD+yo+Mkwbxb0EKn4dquyx5yi/KSo5tr41pK2aJNiFcDm+f0lM
5INj8+sXURBhlokvO8TtWLiYgerTsntXH7Zuw1oqf0Dc3kCnheQrpy0x2PUmgzAIGCdWXSpHJ977
n8ouF6y41zAmSa9aZXO1CRNgVv/BRiEKsYqAeKdczkeaQiuLxC6iTwNqlYtrHL+DTBWMp1QQNjzC
dv0NT4+746RzIAmCUgD5D0nyJtVBJQCW1KG0bxx7RoL0Veyb3Tac+2mzuomNIdjDGe5lDoen3fbN
tdOWDnqjtHoinpKlThfepuKjYkyk9X8ifK+C10dz6Mjq7xGoR/C5wOT9w8r0rzD56oc3atSKIAsB
haeMWDEoB+g40z/AzfIHe1s6LEKxzbYzzWYHQ/ce8DwWlc3+aBZuhIBRFv528hiZfKGydDorZmBy
euLeTysTgY0ObmSnsmItStE73l+q9VIzzt/RhypS3E1t7RFB2SRwtr/lZ/YDrVkF/lGfGpNcUF5i
kKaVZSQdhElBDd+p7zpRYhQHVxVmKI/Z7ztM9WTxTca6bycBW+B44SC4U9p1msd274XBCzddGMJ+
EbITI+aDXztrYQb8dHtJ+Y23aarGa1ZmjqVh8GCS85Mxcx//09EDNt8jf31BN4HBHA4P13nkpae8
DJQrXgsmJySg3j4mWxXbrnxgZTt5tDJ2sIxRZtlDewoKuAOMNLiHV8OrhQQ+gqgYVDByQdeOfEmQ
A+6goO/gdMkN7AGtc6RLJOYDjEDWM7blSXhdQg8Bodi5hbQVcaSmsjAhQkMWIdKXsO9m1Ws9Ps+e
ExmWOg21fUKVBjo1bFxBRHGbtb2FnPFNnuh0IXe5jQZyYCJgRureH4ztYYUPrF1vkGvVHTgTy4ja
9+0884WHPa4vXotry2fe0hHd1wsUl8baCXM3SnN6x7ULxFRnnhhb+NdJWfP2IOGGbotXBmdW6jJU
+EqXQJUs3HjGiWQaBzVoWKLFP3rRRjB00LeJalCcUPsiQ7lORf9kH0dx6oaEEsdIgD1n4nOZ6psQ
NxnTRznwPpddbmJATffWfnCa/bAxjxYNO1cTxmr1J9hZdArD7V/lKCDMwDS7usaFKru0OZ9315IL
6C4fF0l6atOiMXKDt9uflINXuekg8AURFSv79QO33M3Lsrsqyiy++tGaHlqiEmrWUunt/eoDY5mq
URY0QHurXPKUAJnPgvW6/ghh0S7oGeyllBg1n+hcDGOAsaC3aBgcqsIybXoYRQQSDJ+55ePgymhA
kwKaKY9elr4waw8ugnW+2/tNQc/AOnpYiP+wcwWr1tewH1xaNMkFKgxuxKsaKm6vPtbBCVFuYcbw
7RyFXL2KI2BQwO6tNKvOZQD6rgSj/ymVHKpAKWIxtVuHW2vTpnYtylhikBml3nenqw==
`pragma protect end_protected
