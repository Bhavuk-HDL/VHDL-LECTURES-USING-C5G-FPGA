// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:25:36 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
ka5YxfzL7YSvhozkOgG4IFj4yzu86yKSoh8QPIzZTLtNOvn/MiW+e900JV+thg0r
M6jZ9Ur7A5f9emimHVJ6p2ONvDK1t0mwgk0EC3sjFcNYoZ3m6+aUJhxVmMG+WZt9
dgRJfIgoX7nglaeMEw2zcuLIs0ZN7GDsH0oKW8mQzss=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 37216)
oGpX72uKRi5AMVFk9B1a22QujfxD+Z9CLwQdykSl+d/wn98iYSlP/O3HPUsdR1w8
xcVihYc6C4LchpK1twB/2OcNe/mP1q+wVr8udKfQnvqnzgH4VNozvOQM46N4zGah
8LSLqzPsIirsuChaz8xZZjRF2ZIGyCLME2vt9Qn9wXPUSSaxjvrBKmXFIB9l8iRD
gF+f8GMZxJ2gyFxTce5sP/i0Iy8Mstcih9RPyB0SF2LRZ6TguTfflmwTDuNsqdBS
5f4oDAh9aVpZnRoyLmZvv5J9rWHNSexm6NaLLUFgCxb+3oyWlVq2Toa9sTnu0zg1
2/407vT06bE+nFsPfaq6Yn07NmscloZfFig3m5aLQ1RfDqDfn6cKNnnmxfe3dRTX
sLweGdfkjfOsCbqu3YI4qMlhrAOTEdxhAgMF6OXOiNqWxMHXq0jdvgLVKgtHHMjm
lc+dkU227wpUM6gF5nuCsf0gVUUjTkWJ2Cmn9HrNEHuv/18YkW0gruOP/TBLBKPs
GnWYBSnDDD2yGjqHkEz1+x2KBdcsiovOsfILEYz5hTHugNniHkJXKSHIyLnHETEq
vibtParlKAL0A+KTC/O8N0NiXkHlOTPtm9Qp5WE3PqS32WmnVGr9nD5YFKhnE8nC
2dh4hdD8NzJmcpaC/hDbFIK3G7L5AXMRlHX/SFYA8J1wWN5nj9mZbs5lZMMWhlpy
XVYhZ2/I6rnrdu5xvhI7Dk8iWzXVz8wlBnf0GY864GgUjajJc9A5qE0zUKI3qJof
Uol8W2YgVCzRPzGbuvH7zg16siXxLzlfUUmtti/TjkKgJHnYZWbQ8TTtfYxJli0B
A8OyK/m//miPIEdKpyIBEHvSUqCBJRrIA5rj0nPk1JJWiT73MTVc50ioxNqWWZlV
DSHcT8RJAWj/MRGZSMULJ5V2rYgSCIZDAm9iEXsCGJS3ywsj6MlfgUDkeM+0qfr4
EIVwQbejGa5ok+LgaLgMbRCBlo/9Zj7PBjWxZWt6l4m1Hf834zTpF8o4eH8yA0es
Qm+8tsH7J+Hgpmf2S85Yz1I2kPuD/sAtaIjoC7tTFttdnu2dE56Ys4CsyIfKrZRe
2crxo8CcKLXpEsWN9pYqszp4pcnpxKgfHE/woCMLutTf+4BZbZGDhz6FuqaO2j8W
oOd7YHphny2xyzVXt5Mxc8HHf7wwdnv7Y3ZFqn9fZxMGXQ9b7bfATRfCHi2Wx97X
MIKLp6UWVQbt4/FtnYQ4nBAquQPtrgOmXc3g4EcSQ2/hmJTuBHoRDsuuKv+rXiPi
0CluPd0a1PorJvZEYtHwk/GCCvBg88lt7B18FB6gYXlwWZFymvbXrRxcUj+UCvpC
7A6LPFZHIPcGHtymDqQEpKeqI4CR0L1jR2pZ7/k732J5ZWPkx+mrtfO/xe4V5sd7
hJec96j/jnfif7MAhB28M5uumwBraxSjhOGr7NsoSrnfmHfApSPyZ5ENerlAiqjv
hC1yLfdh86A0P+omqEgt9MClI9G0eAx1QlSc0NVaBpl5qJnpCnbV+UR8vw7W4myi
W2UI8GUlbo9Z/FFR+liTwDvlGxNlxPWk1MLIVAVpTxble0v27yJ7kEqCxUOVcxCI
Ian0e/VfuAlnV81K3s1DHrCWtDZ5rjM4fX+eurFzh+d1jcuxGxzpfPR6B96Lws+K
xa223Ag83m2Eda3IKaUoZ45XDawzOilpN9ragu+Sg1LrUyQw71pLMNVB3LSEOekG
x0F4uFCpGSb2V2LkRX0D/1nxVyTjsmql+/ei324dkAA064wj3v3OFnmHSYdNfgPw
rNrjEofPVJ/csMNKWo66oE9jPU8+NXzvg68QdqIEhKc62g0j20j2wTm/7F1weasg
BhKu1OnXu6mzDvNX/w3oyZHheJJlFdoEiY59XbPqnwS93xQvD2L4X9SXbGEnE+ii
UzFfUINYb5gHO3rQzSN+Jz4f2oDpZi4inbwuU/HSh/MuTGgq02NlBd67aoB3byYh
yCAxnrVeoXwqPjXbJvN98LjTvKRReSUwTh3TXzs0KWgY07/fcsim2yZ+XlSahGQj
R3wO7qmScev1Y6CRDKioXfGYWKKxOs38UVGaaDOikZ/GdKZvkznMZpiPmtQ7a5yR
MquG3xFF8u+IHuZ8XPaZEyQ/wiwQ8wRf2j7WUee6Cs15cpoDTu4NCynbJa7kZOTw
6S+nPfyWXp6dA0mFcqg6SIQVu2cW/yjTmKOsGcqGbgDZFhCmSCa50azCcUhipdgO
73hgIiSUi9feVb2zIyo0CGpblvz8yS6BHrZAl0DdLZ620C8QxaHuFDcjS+GC8ag6
ApSE2POJkvifQe1y/6jm73I4WU3Rvv3iD37wj+VX3meTF8gvuLy+tX9HikdZbLUw
STeYnn9XYqtV1xVFnfQlnXc4QPrat8WZsnyoQoithfwwc1l2g63OGsRGZo+jOwjn
CH9mm4OtNKbAgB+D3JhIThZX+zkG0z4HoxD9JsfI08gMz4lWwEeE0Sh+bPTswkYJ
wbYqn2VyiYq89Jgm/OA46Y0sdRq8+HMGUbFHpdQz4QCe85/0MIaWQIKWPiEM8RMm
3BgRI1Kub+NlMDTbL+L3T+u/DwGNSXVPAdyb/hoMxf9v85DsjE1YvQgf8jr498Ni
EJN0qoC8Mv/wjr7BeTKQME74uanIuZGp61a2By/3QsyIRfRiW4xBhMQO67hKkUx3
Hi6ExDiN4AdezaSOdQ+/YiK/79pmkkFyHKAP7SZamw9CBJ2C5/TBeSeMb3Pwf1J/
ri/OEsJZmRv4rgeb51L9hQawDEuXvyd8vL1RvdkTlFzWlYkeOIO5s1b+oYwQam1F
y9SJ+jGUAsa9rYPkSkdzUbqftO/emAek4ZDBjy3jkKhmaerwwBUiDstNtEqOfXKV
dppcNMHeDoHw3BspUg2XGXwYDILo5oxqSVIeG2SgdQaozuZQEypsMOUooUu10l6v
ySSrGCB5SaqYpUzU2KYKBxyZOTpngzdCqIAA168NDrGcgd2FCnyjwDeKSYMjU0ht
VjZ1xThwPBlPMCKz+FqTbUlja6TZU89awfBmSTgS3rVVxMiTqaoxTwZ+uJjRasfj
ksMK3eaXRcaQbO/ZwRL+pAVxxA2Vtm1pVpry0EkxIUJk4o5G5C13xjmdJg7A+wtx
TrEvfpVMcqzt2B1QXgH+yGJpDPw4PZar9lPVw1CmQ1SlRUrq/xp7FgeORHqj5ghk
N2mUFgI3rzDjzdMR2TQCMA15LQErOPL2BIFfENbrRKcfpRS0SChbikxAAEYCYvQX
RSWEouVrWZnWz+FbPlVyMDE15Ds7BvfolEkvyF4j2rG3HZW5NJd+0EyHRRgXxjaY
Mp/IjvWPWb3Nr3KAwsL5K30i0YV4aqPH/oIsTOVfmP+rrJg5bb3N887tpfhUUQx0
C80aO5ni0y/GZq/GnOZZvqQL8eV0y8meu0inI24Q7jDiMswjgGvw2yaO9LkDEucf
IfNpPZl3rbFXTjuvxx5hg6LQ0+5ulp70lqIBVZUfUwLXHwbYh/bI3GGKHG1UghEw
JXXthy5PMx4/KWKg/q+dsw6IngvR5pgN+gycX7wAJJ6SzA/n/t/Ymp+NHgtrnAIT
8t3WljxvSyVtBPWXU/jspJTdSKjDQnHbDkxe+6HpaLrn4Tyv0V4xFQA80N0KLaCU
ZJXheMBAMghM4tnUBLhVEeWmhXjwJs/azAmL8M74OnxNGjHQ3GjS6nAxw2tsWalz
mvaV9zAJuJDkHk58JL70LQTlDEq6Gdj6HkbhT8MSHoUAacY58hv6P0C+LbFb4VOt
gQXVP0Bmw4sraDP6pQEsoPp8wXVUqnyhbQlU3AftJUHrxXl9Pcg6tnBw07ujo9Jl
1w4vn8TDqLjiLE6nHzyQ44HTUrBXTeVq/+4zLHar7f96XmB6Oklc26YBisxgBy7p
AGb+rTkZq7/1pY0kVwcmpqnfm9lbvyeu4ojJPZpXOhyem5jvPYuKyVOUwdUMST5r
QWHCebp0sR6eGzZgTmMwPZwKxVZDGu3VbfkI7wVVyKaX8KfHHvN0jeVqMvDiTelW
weSontbg27afdPlEok+Sr8k4I4eZYusvhwgN98JvJor+LJh0bul8Q1k1x7Fu6bL1
EqPYomvwxWpkBT1i1M+fWKPQmFH5NSzHR3Bbn23u8ASMYJQWu5SQMa09PD2PhqIj
GKEIpv9JKXjorpjb6ieqAPsLsxjMlo9JEMR/kUMrly1GP/UnhOlDQL+roW8HC3rM
ef5IiytHyG7LL81fWEqB6xuQyS155Vs0O1szBpKdQyE292gwNYGqUHKuW7Hg4KWp
uMlCFRMMY+M6R4+zkCf9D5QH5Osl8GhmwCWOJ2V+MIuosycBx7JVVrsmnpWLcPEz
CPNZDOVFgQHuz8zLNGSuBcpyDY0KOWegqMPLulqmFgHaKiDICJ688U10tk3NKiig
d8ANqetaQQ9NYRspRVl9Fn1JaUwFR25+u0oY6EyixzA8hVhOsJsaT+aDoLV6D6/z
5RIB5PMP9B7uN2TdqY1OrHxn+0m2ZVdTOkOQ58umLDH41fWKLhqHslH4ZLlo9eS0
1IowtKsaFO1LAlwJhj2gVkHVTYxsUBOOxzmBnTQ7OrmEyFk5FSgLMygf0ZD5cGXO
1Rj1NKIz8gLDBlze7v9zEPpeTWmSkUWPD6MQHH4ooGVdqcL4cjgZ8CpCNSUC/Bvb
+AZpSiILVLh73ashOa+6N7hkl0ZJ4cGz3e6uMdJkzgGgdaIe49dxiB83Qa4740g+
QNmO8wapDDFoLSDaschvnVMf4A1ml+ypcBhEa2UR+eqiPIfuPGSKbY7C0oG4T/HQ
hEqi5LB3gOodJ9je/VFT0pDbORQBBoo4sq99ExPeMEEM2ulKMdjsehR0BNp/Hf6g
9a4HAGl/zN9AYMaVhxornPYayoQetxQ+b9xCPbYQaJqM83I+E800s9yjROEzL1iY
gl8/2qiwQI0IzUtBTqnpCKrtJabHuQtKiAmKIPTvnkZGDpM9bR19ERsaBhPR82rX
IMyBqhJAg1HE3O5vnGzWRYzY4sFm8K/3xmMFjT52WolnijAQwkXjlM2vy21QdE2/
NyUpG5qJaWl944/unkhUQ6xP3epRBPvomRlwELqz4B60O9so4xZM2ChGUe6G535z
/0CDzadJJRYY/MQGNAx3iOJnp+uJuDO2wYKGSeCVKL60X0EedwPJq7vLO3xmcrf3
w5pUrDC6/BJwG2zJRrF7u1tWGBDlQK5zaatIonWpW0jj06Tiu4QYzfUvSNGZeoNT
AKJVY+QxQm2hPLu2/KWAmdt2BBI67Cfertf8bd6AC1OxKqgIfTzuZQFh+IXrTPKL
ZRnwo+B9VpxAAS2XxMvFQJL+L/5TH1/tzdStrjfTv62VD6k1lYFg1QZ2hJ658bvI
Z6EIXJdOLEHewUmn7uzb2XY8uX3QtJ/ton8JRI1jAXhl3dSosnKjk1y6lC5ABbrC
t442GR7RWax7ApnRyrPBurIHHWYBB6oRHjuC1Lh+qxvDqPb6fbJXWwvJu4cBWZx7
5CvwcnPRaFA6grndXMfe7kAPxvk8vEt1Qb7kKf2AZYWVR9DQUk8k0VvRBaH4mRss
Yb7ZHf3kmF/TapboivzLmdNo942WXdbty3iKFGbvgeSb3jly12ACVEmZg6eIle94
s8HK8HRSFPUgRPjEbKEfvZ1LnnIs/0zQZteeLls9kITykClBgoanK4Fbn6L6T99H
zQ1jQfjVKtQfU6Xw0wpOIFjJiMtgr5MKL/VNjCT5srLucoi5WZj1GaKZOaghg7q2
lv3/xHBKDVz3BU9FDMVg5gihRGFUS8/tcPQCHgcIMFxiNNaULK23nD77MkT/vErb
sVuNUNL8thoKeQl2cCzwNv46nlGSazb+po2XmtoKaZRaMbAae1O1/p2jGlAt78+E
qiOX9N5hXEM3gzN4sxWf9H0Y8ErK5qPN3TIEea7ibOICLk842yKhT7uMVf29lTYv
g7RDutInxrrMxR3I+BQnrexhQd50xvpSdyUS8/4HKZQ/9UrkK22G5MwH6Py/aS6s
dznixxhhmFmtsEtJfZMWIPNOwKXwUvC8Vhhl0rAncytFR2OPpLrKE2hPpcHjTOup
xfj+KJnGZbAsmzaE37VA786NTcw5ZGmrbL5JO06Om/vAiR+ZMRzLO4J4AmZdw4b+
mJbeg/o22DJ0qUA+WONE6Ufmg7MUQ+tP7IL2GAvNOXXYGt9RHLyGOmS78eEH697u
QE1H//rXO/DDG5GKzc9Jy8LHFLiFiVKBItT5Lw/9+/SzGSPE4QZXQe5Im3z60/f6
POQzBzN6gCI0JDjnRTFf/9OMmdf8UI8xYP0UiVA+nvvYwUWjNO4n7VMqhiS2fhD2
OIai2lhob23aE0n7L0UWGFN2y+ANzbTXhBHD52JJNBjRmJ2wetj8xugj+rBm6JH9
p4N0XIYxF4WKEq7bsyPpE59c9v/RzRywZNI3ytBpvPgtGCsRO3aofglEBTcbeLsD
sVT+Rk7vsIGJCU4AZQ9wMLfqE3AVqnhkwlfJP58tS4ey6jg58aWhhJqhOm6p0TmU
kN6cvexpcDZhmJ5trUFp5DXM9R/hviMipgJJAEhdW498lo2fsFE85YVBXob5dvAt
lmWsxJKi1N2YGi4LUCGPFB8HODfr8DNbZWuvWhHjDiVTg9yaUFE0xfY88U03HmX1
dh7sOvlI3FQ3HQfTQuvzDKCgLI/rNALHOKH08sfX2I3cHMKrBbsyqW/KuDI5icEp
K4Hfg3h9WL/8znqXf5waXZcgvcFhO1EnyK6510GMES2dFTcTKu50vJazS/Tgy2X2
3JIazdp6hlJP7TWnwmNiYZLpc3C0D1yEY4eYxcuY+FE9shiqEktanIrHB8O5DWYA
Fq3QWwkX/2eWy6H8UxtqcuWmXCu8XWf5YeanmRHtt8pn647bYFxbPP7Tt9gmFj8r
sJn5QO8qu/O4tjpNwh2fY2B9YzyZZibwoA5NBbEJZExCzPWMhQ0DLHHMW1hoh6Dp
uUPBaN/GdOJpZOpgzPB48Ew6ZPf3FcSsLHyfhOLzeCxIKtZvvKFRLLyBNCEChXAU
e1Nh7WhF9jPqYVjImp0OGP//ub31khkPmqYubYvlmu7VGd8wM+l1Ei2ZudGJt1XO
Hspp2ZqEmtebX8oDvOWdGCTqWa8Tw2O9anHYlPPGCYUdb/4qNpymGiWpJ1S54W3n
fc7hJFjNj+pFsDAyjPghWeljhO1+xFecC2O9tBj1nk8vDLXpQ7zSzwS8Lhfs8ssV
JR+mYCEKzkWIIwWsNuxAAKFbY7Z//ynrx4FrEC2Wzx6zq7CcNHnKF+dtO7tbgSOv
KQZNLpjFAQwMhsGzJI+r5RrvV00kSIn2IVTvtRdgG1F0yYhQJouh7iNcolTdvIzV
r98wXG0KJ24JryLkKvay6knxX0B/GrbEmbMtvsBJfWlHbiFjEWcKLAiv8dxBHUST
uexkMD7ivzomtdhNJiHZnBplovmtihpFt9CLyldplhQAz6+5vZsQImBd3iL9VbST
qhvXUjkxfEWI0BghMz1M+iSGG1tGc2XbVm+X4lUwGitvBMzBYVNqyN3gKY55QtJe
Ip+XUq9j+SlhRKle/RF10Scln3ybsk31q30wlMIpJtctqaCJUf4mSLwTUB+MbXDh
mbASFrYZH1RCznhbJmmVlocfd5/1tlnWK8WLoG4/BMkLl3UWfjnGPiu/20SlPDwi
eIQVO5gFZ2hq1cvPJsbeJuR4fI5HglX34cvh+lhAaYeBzZNHURBr36zOfhfB/apW
zC+pDnNDEsZ0InEPJ+y/jfw3UdYfKNYF1VHgdOxzrj1tBRUMITpeXAkxlhVoQySF
iy0x0Zrrf7zdT0N2Je3jPOapNtVB+Pz0ZZlWVtRttXx3Fnf5qoLDpW11574M+m0J
1Z30vCDgRFkFjgXg0Qjz29iUACiHzdEMUcZGgUxV9PLtfvY4foQpkEPn38ljbelY
bWEhZ1QU9PGgvMAic2eGj/cVm9x8jfrTXRXSoK+h1uCxJL+VTOJ+zmJx18qu95Hm
nTpUPUWMf0BXVb4HqEsT17rZiUld8axJRrY5mFvLwXJKLkgqWn9xHvhornBbXv77
TWhybPa+rW67USSoJIlX3lahcDp02Z9evOFHQkfIMuZ0ViQtQttKe6TK7Vckd9kA
LPEy4jjLgbaOoprScnCvVx2hFWnwk1lnbDqOOdzqw7/v2e/NEdQTwh+FGXrY66hU
MdCbeNHrtzfvHnsPDIGRe6afyeTbsSPoPpf+x8cxJBbwqhO50ryGKD5JZ3vr3E26
L9HEtWn9Nf90g3cizfIUMYVYgLs/DtdBgYi/gdESewHCn2C1Xo6QgPQT35BwP8XM
8e0c677rojAioHbpPvIZne1rrptuzx4Jjn+mF17rELLjQKyGc+uP7yWMFbT9SJEf
DYQaCPY10DPDM035EVXwLDFvxt7nqIDYuEzKPjdIUZ2cHRRCkjBDddyLUR8kKTro
0Ghg5fTZe3s/72F8XU3GPDh/W+qk1EfuBZnZame5ldIZXHLENNjzN5vFyP1uo/WY
aRUta/t3tTV2zrUaFkjvWpgG2kv42+ER+sUOLFreuCQ7qgPNQ+t7Ud2QFTKhWBCo
p1INa25/WEjy+sYqLcs9Eli6sSsWP/4jL3dit4VIS+iEUc5qCSgKhTSryweAv5bK
qfcm9L4wOWbvC4C+AIBxji6N31OEKNXF3CgEQNMX4MDCEMDnPmYv+QH6vc0JwhFG
fKDgdNWYNTl79aHwMAeoCYD/uQ48VqS9kJMyI7vpAmyTkR1MGWzKb9KIkuPkciTw
1i8U46VWXQKKMQlEoOX2+i94K8afThcd2zX1J/mRcSazhF1so7Z3R4I9dgYZzIsO
eQ6nXvWdC36IRM3t9bYMMnh4guNpqckgVRVUT7ipVIXzm7ixJHsQ82aHDz5hKvws
oIUwuldVeKlMmtjwiMC0MymVNYJ1XLHM+l83+R9naaD9TV2qt4jtt8WTizPvRf8+
9ARe0IJFkx+SDDTpvWTx1uqK5C9L4L99NScCSKc40H1XtygF4TfazwqZsKe/ip/4
j+7w4bhvU2o70FVW1PwW6fAntPdM6klI4FzKHcV0d+xFydb/t6EuuYDeNAVHNW1H
YcS8pVr5RkvjSIF1ZLToI05AOuK3JYhj1dR//6tygrWrkumi65jMCJQ28+AGKhMK
tChCaUV7L/yDg554gwJipuBv8sPC96BL1t40pAOukKf8UZ2oVuQRhbgmgOie+TeD
tm0YgvqQQWKehhxdo2Z9sQjBKhE/AA5+CVSVYwmVSWO7JLC4bzvfoPNDDFS3Prl3
5VjwZ2gzROWoac4UNAOTMKGsgMcbaM19Whvp23celFDmNW4DrvCGrStvPnA39FG6
bYX2XDhu629LbZhi5V4FeU1EwqtyAAw9ChE4YPhlOpClafq6vc3mtiw+YvvrRQSl
Zr1F5JVCBFqAneoNHOBKHOq0pEPF3f3GtR9GOY5ejHCiAATiTyx1Lje+EdgB5Taa
tB272uv9JYl9FL1ZIgpxU8co6le8pfbA+wB44pPdMvJwhRiMG/RibwgdTJRXNqB+
wbHv4WtUM3hWP/pNtJ2uaC3FIpvlJBeaekZa446nJ9PJUDlZqdRPXPkOnJVc728T
6Ta13gPW47m7OfLGfbDMLdyAO9loGZ0R8wXk2vPHMJcxrfff5J8YLXo2iFKjjLk2
VOePvmdLM8HMxT4zg0Hjs3uvr1CzCadKfTeUHrYYvnr95d7wATQ17ySzgFHCo5el
ovnRiEFRJVCIQqf8BB9MpzB1Vf4ioirFmHzfHAQkcPOY49GyDJ4brxGe8AXfADTw
HmnjTBMk50+tK3b8rgFEDWiEOPQ1h/JrBstu0TGd/fvjAwcEXeH2UEiwsWFg0V24
tfBYVR6yawsqMBepPTba0+1AqH/pdIXDp/vSNO/4PXuxKfOzCVI+QHkXY9Wso3XB
C4i4RMeozXv1OeC8sIGxDcgUFkEeA0r4cYWcKnZqKomRX+3E9RUfhTSsOFyGwoFV
PtmCi2J9bs+E4GaZu4krFcLujidva8KABqp0anaK1eku0fixrmGXehGS9WzHiS3M
SlpPMw/5b1RO3JpudCHSvx3SoxCCEhallKThvJI961IcdTVhMrcXyMNfNLe2xSGz
1Frbu9JOhLcIvwj7aCpPtjwYRJOPiB2e9V3d+d/mQQAIoiVz03S8Tb0k1JN482iJ
G19eaoKgfubyEL6WJD3eVZVKX1mLZVvPPjSq1PWHXPi0ZvEmU59g2Q2tSBVzQ8S9
rvF0tex+f6rbC83eVprQeX9pNJIhK6dJ6KdPoq1p9hmLMES82I/ooSOxNcxo7Fg2
j5U4YnXQ0l22/DXwPqZXww2jTXweb2jIxglcJ7YcmlJ5/SQno0Lq7EQuCESWJ8l/
j8Kov7GF/f1MvN8fAXBpuBP/NXBx9QbvCBrufHCPKbdhbptSvVZKHmS3uJzk5vOj
3xNVfuLM9yCXXFYpvLUR+lvtBrXxlR6fdIAlwruxXHo147519pOpIe5b+FHIvsu/
4/d40WKSVJmpw8F7ReBwWD00fABTFH9Z27fpcdN0H+iq5I3Ia/6jqTjqemMpmSsh
JYw0+CfCBJyidgeL5LBCsoqmjIeXxbD46wqCKokU4OKH+y5QWvZg3HbYcyjU7FCa
UG8G7aimI2m7yO6pNji3oc3fPa8dOzJxq8usGLmvS+zu6sAsCL1pj70g0ztt40Re
Jx2QOvDcRHHk+xq0P+00F8ipq1Ap7bP7lTXG+uZdFjFXxHcx/WrxPsIhTDPqKCxj
vOPPJZQIybs4Vwj4p8WRDkp18rQYUyRUTJeR+f5ByYr5CH+1kFjRUEunXMohJdiv
SL93X3ymcdatWmrINTV1OU0xydCILCFljvbC7dxePee2FTR3Uax3wuo3BHqurRUw
KpLCgNEXkekLSokWLtI5SMAki5bOZU/NBu2U5eT1bODtPAxJgkoC2GOlEDoxrLvX
mlS1S7YiIxIskQRZ6fqj9kk/q81Jn6cghIolZQpdXyVm9n/Fg6ABGKJoPUgfJeY/
WBgVC2uvBa1OZiAoRACRuFsbpW7LfUucQvKsEeKPd9IiUiTPdfI/Qg1IbAuzr8x+
y7Jep1zXRebT8UPYXYkCG9fzGigWFw/W21LgXv9UA8g9wRYedLRww3zD6ZNZkoqq
FPANphuOZkZESPsMq+PFNM4Ko8+76TLdWny4JZEx1KLnpsTBkNRuGrHB6xSgmLMH
aVtBKU6lQOVjJtoCzGlIHzVy3Ir/fktrNGM8roJEOuXRsBmtWpCHoq2kCp6EKY+H
qTXVfb1VRL+StFvSFk7uxxJYZclNfUWXjQ8hpy6a+lURpyRiXlklbQAGn+UixXqk
z8dbhKiqzKUN+OxmX1Rt2IvGlSG87cQg/xXtbXmDirM96JZfT3o0RybsMRGXb2HW
XvQWoXzNz2EJLHfEBCP0jXrh0mW9Uv4g5QKBfj+XcoiKVffzfCu5zVjlchGsK+QK
8yV5hQkJdUMp5WPkm0I6f4sqypoNWA2ddJvI67ZxS0Xg9CD7+VLjy4qBYNZOFcpk
X+5kblWSSHTR9u2/O6iIoNfVglWpIJ4RmtJ3+ZWYVhQvkTmdSO0W0WR6ADUVu80U
LTeMHW0aZ2agcQcECaKca38rXoKfLGVdZUnPB42GMP3h0Khilm4JKcFNz4lrTN9o
aKTTo8PXkE/dsrPG4rnmooj5vhH7z8v6oY2vdqGgkNvGAjVl4WxjuyGyNAkHRSgA
TplVDfpKn//JJoxlLHEH4xBEO4eWwtx13zHoFdZ5YyUjxwT4u5SHOpffJv4fgsr/
ssm5sfy5Qyb/PtBSNJuyFeLNaSasNpV2j5UojRPxGp25vZa4oh2+zWAI+Ln2GEFk
NFAm3pTEQo4bEu3KxANf8skbn55vEliqmc98XIFnZpMyX8Hqp9m/60N4h0mhEuJn
8zK+2mZcUjLTGk7IAjcatGGJgyz3QE7sW2Kge7r1H+XruAHGUURxZAdAMpPs7hFh
ns4+/XLcw74fpl4xlANEjDk/4tFAme1mzooraBU3I2Xmef/r5z02KS8I8H0a36m9
vNePsZ2fBXeMOiXNJHeehPd7hz+/dV22ifaLg5uh84t7gXW6PvIUoThXCl3rjaO3
k5SVL/Dsh8+fe3HvUp6cox9V33aKLd36+S6vQx1AUP0DO4kRCxnswXotBgC082fJ
7sG6ocTDSU01dnBJYYynJnMQ89h7mr5n6GOGJfsrOM+n7fPqF2WT1BV6kYfcS3JH
CmjI7vyiR4VcklRJzC+oub8UI37O2pwnGKxbYIfXnsD1jhMcZfZjTm4LoqVE/srr
BsrHC0GuMq6TpA2lA7da34LUvkbspHzHkuzPuyQx2itQ8rbgNUykJAcmn5ckUntj
4SDSdFP1g89uiFwYlVAKXIaMcy4aOKZDn9RRgLHML3NRr7WR893yzI2zFVv1k4On
GRdEotcX5UKpL3ucZh/lcypT/qniKCEsUSKYJb4RSKfzt8mPJEncyTing2jIjn9u
oEFm3Q0sdXuof/+JL1vCk4cIuvjpretT371KYOdg/YmRIerJfBBdUHuhTH+76q5I
EdYZ6LAmC/6aY7aSXmavyGOg3vu+dX5SkSJPbBrFfNYMTNRyo4aP3YBg3vu+Fgsn
JR7E963k60q+hPhNPo3oJga2u9xHBpIzUwYaEbeWE+RlxVZSvnP2NJacxNEEw3sY
IOJUcUpwR6OWwntHCOCZmGATmZ4hywESutzrYr9lKqTiXkFbCP/jijGbjMkvH81p
dY7HiNedrX2D9J9mjh0rE9ozu4IrfI+fdruL0BCEp7nnV4ZqvL/v/CtVIIdOdH+B
2z2PkE+uBqzsMyGun3cuFIPsiFcEUOyux5Ms/KQZZubddxuxmjfwRzLH3RWuodLD
LbLkilJhG5GxB1MT8dUQCTVmi9JZmQFN/ZoZAeke1WtuqNXoo9M8qFlPdvxw6CMn
9woa3+mbTttQlXrpSaQ9u6PK/Qq5j9k+2ntLp4EaTkN0sr72LQBSrx/GKhKjdj/l
L7wZNUETl5Vs9waM6CdB09XOHVvbWF8x/cRY4IrfosmT2SH/PCZ5yu5KrC47GUd4
zQ8tUAbI3zQ5dq+MPrpPgFdVEIPJhYZQAfZUkCGTIN3DrJT2LTQslasXQ9pPzfpY
XKx6DnH8vN4rcxTtvef9yigwBXvqS+/9rE+mp1+1JzFBDVezVhfOdMdSgOzPfh9h
o22e+gme7Ah9sTb2XgzOotnP8zAna4YPcblcHXTMjDfvvWWtYhxaXDWvjZELOCzq
to7TgtSkI97KfDApZSjAT2cQ0ytzXj2OBzNSZOjNKu5caVyPfelJidH/Y6IxLOxf
xCGUlQSRYffW/NH6tfsOrbeCh/8G42fdc4o5frtNjoJtmE9c9h0otLdYNB39bYDp
zCvfoLSbAa/B26q3Jl65ZgeiVNE6Ay7PY6ydNlb4iwR2Gwer0lC3rFFBAe8uOTY/
Ih1KYqkh43AebTZmo51PE2CXqbWNtwBSYI7K9sDY0QPcKLbE0QFBKieKl8eGXCAr
zGAnC0SzCXEicqOoqw9HVmNIMYhrPcKCGS8Lmv/50vi4Af43zKW1zSiQr8CO9yKE
D9QOndOrDtoMGQHCltQyUPaCsATlklznI9QhvwwBigYb1ht9PCINE5ymJkNGKlRo
7YZv1Gps46PASjVIRAUHovUQO3TtFSgL3RPxWXP4aT3CJB1rKR0+V0w4Md/BCCzA
jaPO243Z8Zsv7KV8CO0dzBequTNM5NL/ltQ5/B/foDB/FCiyIXevBfchvhtooKGo
qQbx1S30kiGS+QKCARb4yupKybbmxpkSmW4C/H+iG8Ydc0IBcReW7I++mfePBAfn
tjRgCgMh2kZQvnef02OBz3/hubnRTSL+idyIF7NnxZHA+jTVHlxM+qoJ8C6eQw/i
eyEZjXle5Hf3yOp+NH1+DDWQsjuF2bC85vbCk8vQpCuEenMzfrHgfX9mvTcv2+3s
0FEgG4wP0Hn1pluy2ZgAyQfTA2cKSR1qOfv0f2VK07vDdLzn4SPFEmUVNFNd+T1d
g9+Xb2JUb78yZjfI5TAS+d4wBUD+Kxdklwnmq1rpEZkidfFtMnPWwLAyPaFua2tv
e9BESIzjNAOpQS8d9XeqSez5S+APfZgXsxG9SxjOKr3ebnbllunKd8L/eXjROLac
E4DiSEsFVHCtQVdI4UFnymFr8JGBUgnnjaAbJB2rd2xvrF2tcpT8otdF8ryBScg+
/a62p5KeLPnkSa9nxVUqheIPZsTbCo+Plf6OmLSO7EQ5CO3Tlu67yEUK/VuBk7Nr
Y5nzw5ozfWasLQUhNBKVBUm0/EsjyvwnubvV6Bz4+MQXS8yT3i2XVWn9l8a0nhZ/
RxJF0YMUaUid9thVhlgo8NyGBkIPpBV4PAIMr/R6NOU8cJIqtSyonXO8Q0xWjH98
pSOEBSdm1joCN2Upk9QnQSXJN5Dh/YTHIr+NvcZzjVeeQ5rUWCNloym/chio7hEX
r3ccv9nQcoWP8TRT8jS0PHcObgXglrH4NNS/nH5oulgwkuhGZfBwkBCRh8Gn0BOp
nl9OHxr/GRTjMsoBNX4b+JkEhSMNcKEhkQ+fTj9WnNwgjiVnMdqQv71+1/jxU46n
35Cm+QElz5d4nf+GygVPQvBLn196bVXugdIP2Z48Whg1SCVPnJASMOmPqAB1zPy1
KK2OHi3yvZThXJYR4hBpccORI2ETFBtDPqHl9nSt+JZf1jmvEMqxPOvLJdZQuuik
ZhyuHF7HNSiyz7nbqJ6pJNtTJLUZ1W+C9I+Wq09pqx4k2vV/2uJlQSvGisMV57iI
LezoOTreNT8+0TBGFNvGNKePP/QEpmJImhbcPvFZxQnihnoDpaLKscwaTUoXGEZc
uZyzwAmzd/+65Pv7IIhyRcVg+JmXDQ5qFXJch7+Y9hN/3JX84X+cWOCwDfL1K0Go
a9oovsNU2EYndWsDMsdHD2hUQhVDQ3zuhD7mz4E5eEZM6Qnjf6EXxj+d6YWLdp5L
NVjqR8/7AGmUxVj8vbDH5Yba2GOIeoGaKkDww1GS7wf3WgKnI5RpRImIoyGB6YRU
Y0j8tk3EDu4wwLFn33isla0AkQIpvAFde90e/EmqzrG0IGdkDUJ3C9DLOBicZWjT
VitXrZ++YxraHIlJOtSuTMOLA+sc1BrUvVLJsFsqry9BRwq2PTSTfJI0/lFq/nEm
zPKccBBnDzZURvQcWDuEk3I3Y2NciaIsJv9VYWqpFxGb+NiAsXkPFmYtXe09eVBR
EFGPVEpreLGaU/Xi2wp6lXFdi7aTGJb/VEjyf2LpW61WB1LNg31LeF5Mtv5m1iQU
v7i7EK68dQiCyemq4pXxr51pW8vzRN/ljhs1TKA0r/SwAM3Qjoeq+U9mLo+4Wak0
Tn7M5GaLwh1KDR1i05QflNCBD1Z083DHDkBtu1c3bf18VX/GJwQV/LleSMvYuLT2
AVlGjqOTQGR0VFQQYVw5p2iJ2YFkIKfbUIXa4y9hyc1AJfNORwSgkJ320QQxukUE
qHYwpm+wEEsWT3Gye1/tFosSQb//znsAZ/o5u2c/cRT+yDjmk+32lyr+ZZQmnmvG
nP3kFsHfgyYvNjOlu436g6xbHiPKfo739NzDDzeXMf0XRnVYSzBfDkXVNpN5TXvw
C5HpUKnK3eLklTO+/kcud1B3mKZta3KV9kUYmAmKbOuZ9rHs2SamLvyF5Xa7tAC/
th0jLkpRGECfbvW9HjeZnP+tyJdOdYfgqgZBDgVD1caqPpRtI61PmVbIc1yiT4Ln
JgsX32rGvenBTWJb/yKj/GJF+7k/AlEaR3dgCpGLH3jMGmIzhB0EBLNaNfEaaBr5
9EaE6EuMdNQRbnowY/4RBMnzae+QDlX7qcwopVcotKyTey5/0nU3UHExvx+8hHak
vNNZqFbY3oAfM03xnjMtxe2zqpsdti/qFEr+f3pYJxDtJ+Vw/DAXhNfBqW+WM8i+
NV5m1rnec6Sy7dzQb2Oe7HUqd2DiMnkOYpTZIitgWFINphXY9a2OkTXrZ5sTnui/
iD/ZmxFsr90BQYAiMmaQjUy85SRXWiP7QI9qk14bWU8HiJs/90czg+uMDRBH7XsZ
ABM/DMHE8Sj3t7C/g+UcdHDkr8dZjRl2nuhCui6pGjQdrExXr47GPsCXLEoMD+v2
jje2PM6qk5gCkcaCcT/7sZ1UB1Id0BAHeztwmLs51CStrfZD25RoxQfa6qhCUVW+
t5WZFgCafP7mOdvLO6fYMsO3+GeCG+v6iTiHti95M/dwinLSKCOUcwHZrCALvyoj
Q1qu+Hj9V1F9NQ3zxXu2hpwGNpByNkQiwUyTObdlEnhmSHOinck623e4RvuOLR+A
opjN7Gjx2RUfJm1v1J24gIcoijwjJNjb2brbWrNslX/xBZrYBTrJvS3t73ZjzMCT
krDlDA8NUt0fGhzuxGDA1Ok4/DnISPB4EXD3foRBNLb6iW/7Kx07cqWAdTFKohZO
agjUNbwoL834lqqCBY16FZWKaxzRX1MDIc2F+UTVh6Uz2McGPmnG3dlB7PcSZp+m
DIEzsjxadhenYrQ1fhOb3NuZwx96pt0jNlX3gkY+7sA8nR/WSnhNViv6aIpu4f9O
kWvcvKGxPdcUM7x2K24z1HoVVYDSkJ+hlvJ49jdPhvoaiuZQoa54nhsqsHESPM72
sT7Xq1BDtA7B7vFkmr1AGyLd3PW31KqE+En9io+UGND6kIYfvuKnbwp2+x66EltV
76CYa50Mkda0s1vdkOseTC64vTuCRhqH/0zZ3h9qCvwNJL+WFb+UmBYpuOGUvykY
j/HafqtGQ5Z73lnZE2M6GJ17g5wZ9CUIs8hcCtdIWi64UQXdbvMHnRQbtvfHP9lb
CCv3N5VFNNQfFUBIP8Mv6rVsMxqe6hBEKOCMqsiokT7XGOG03rcJV/q6YriReG4P
FIc/NsfIOXpec2dIDYZRDWDPYO9RAmCv3hpPYSnuLT+AixTRV5bVR6B8fAjQ3T7A
ZkPVGmowOBTQiDszb1L2Spd+JgmKIDe2kvyk7ChQz6Pdcpmd5WZdSaIe4A19Pmv+
MTeIkStiblynHghMT0t8W99MdX+z4fgEmWKDrPp6fA+D3DLbWqPsJkZiyccAvPHt
fJqV9Dhgz33fq/ZnBhCANAL6dJSmr6DX1vHb08ya0g8XX/15Q+uJqSWap4U9IaOw
lfNyr2QKiSufDL6+HBQXnJTHhCD5m+nqWCUlfjs/HXTBEmu+xqIhl+bv0qCygg7M
U1Rjt9cLKrABClbvg0Y62/zqAMGEqU9LHBgZNR9l53mtQNpNQ23emvvxn99kMUsN
oKf37vpcPzkrhmjJW1ybDrMxAQNd+/1hdgNE0MRoHpaeFCrnxW8UNGa62lxvH3vc
0Z5biYCNiZx5io8zw1Vrfwwg9IsZBuhTq4eb7tjW1T8/91AdF0+bf9KEpj/4bhuY
zG/8UKczxiT6GrwVOzKiOjx2uqAW4TZ+L+mh62kfZQUjGXya3QlxsHle3Q0FqUvf
qJbxG2/9NWzHviF+waZ7cFqZP1xvNms6sJ2qXU/PlvnMP+0K6/qpwEOao+GneUDu
bMUtleYY4afzwmM0bB3MvPLPhoxjCytO8ycI9Vnont6jnCvcgPgE7Vus2UMeHsgq
HTJuZIrYFNBwxvpmg0F4a4vVeYFHL8+0Kv0P49cl/L6MBxKGTZNTPJfpdeOlzvDu
3OIrmEXvlVEX0DJFPCqIH4m3o8GtUCPN75Xbn/lqDwi3HgGox5NpywQCXXLEjkEZ
POtq2WDGQ3JDXWvzrsRSFpmO+Gu7GmB0RLC6GPva0qxkz5zEsCTBm5HuJf/0f6Zl
1NrLPc1C3FzXqHbtYnJz8l1jj4hJTT5hVRfTT1bfBxGtWe2brcsXT8siwB2UZFS2
sr7+0w29Rxz1JstB74dJlPdJwxNHCt6R6B36SJDn44DaedwLkD2YszRzI4T7gD6l
4rvn9CChd5ttVUKlhowpvQ+DJvstWieoKvHhYrfTUjdCIhaoMRw2sIGOT0McjeQ6
WWemCTllxxUR+g1ImmupOt3KRcm0hZqJpLcUkhhsJTBIvAqz+U6rKUB4KM0n/86N
QgrbOAoPqRdkMm7Rkn30LT00XETZY3yJpoxdqXRtuw68ksFkzhdey4PHbo7fmBc/
5XU9jbgiknOjorLUGNocI6b+z2j96sdYcm96+/16Xo8Ff9DVYJ6cTKqNOCl3FWR0
MgpKtPBqjnrP1xqERBaeL+eZ2rtU9nE1wdbBx9ncXYc018fUnyXsPrdeXU3XuK5y
Xxw6qeybj3XGDDz60rD8Jwk6lPhYxNftc91WhN2mAYV/yEDM1e40n9Ej9vef6sCn
+WNZUdrXlVHQXjenmM3qEVMy8bGJv9OYGl4otZZa2yRdaBxTE3DFWPi7jaW0gKkG
sdRWOrK54KVze5P2HHapboBudgvgPiSGI1bFzm2X5Ig3xXFcBKKjI5lB7cSlJxGQ
9nnLUhi7iPTAsCNwNMTCrMqRTBDT20/VolSCldCxMNwmLKaj9iVU868mQ867ejZu
UxayYbdbvMEXlP6sdHbcUh5JdCSkbUkgJz5egBC+3e+aG3oOOnlyqgWkYeQpAsqU
BnYJSM1Nxc2puZKf6ThBImWEHxb2ZXmkpFaP3nJ6163GTiri60pTZrp2RsY9E/1Y
s6J/mocRY87Hf624kvwS2xz/t1Z17g7yudMju5lgWIQgCoEMildzx/s46c3j5Iub
bXnXxNNjAqV8Wg+Kr3vC8xV46nvezNvr+mAiuuam9icl91idpezP5Ni/RQyUt4Ii
PHVf6rSzvUWKltXERJ2VsZRz7ZBPVPinbFCXxb4+DKy93/WVq1VPYjHXbDjnuKGD
ceYaebrbyulVdo0Qm5U3anUTv/HAmmKqTUhllTxTih2ApwWXNMIbmELYb5Tim/nz
ojZepPtHCeZ3FDG+LJDVW1n3mE4OYNrq04yldVyJ2xUMd1ZAiWaiD7iDIX7vjWNy
5tw8BbZPB0HMIgDsjAEJlcOBKrz+PZRzQ3fKWL4JyUPMHCMlvgdQpcunSCVybpoG
WHwk/LebkFW8v7Qat4VAp4krDF61/qkUcbwsg8rZs1rbTpRJ2KHiAIm9lZvF+4n3
Kmi5bYfyog14sUA6Zk8vbulk0drP8phlZFEjpmLEoOLVBOMsSKCqiZFD3xdzKR9F
RfQl0Us8HBPvLJA+WnTSdYZNO+/fuL1KbBEjscN/s6C/10U4FvKGN1AdpNjInI2v
vcTpotMBxde83gSFtfV4go18lH/ODEPG8EgrjZf+/iC1Viwhx8b/hn9cLFmybQnr
CpX2G7BdYsQ6OPgi1bXzXnmPNhWxwMzyEd8iRLt7f3VOLrLNKLvAWj06o7JO0+qc
y3Fi2F/y7ylHHrQbUNJtUFGk/z4k+2Nx2NVqcuOmZz/oeAyavVxC/Bmx518b4EJ0
50mopXJg/zISx3QvMYjEA6jsw3ys8kRNvFXDOXhHEmRfuQeEYm1oZQHRsSrfzi7l
UGwbErfUJzie5ydbXsaujtDGDPPKFXMM62ell4qWseEhPoAlBZhf0AV/PLS9qTWs
RL8tn8G37AxiUUh+hJaLdZYK6grAQHKLyvixqklY8MiRhHE02Mh333+BPWp7w5es
D9Qv4rhE3KjuRG5XzBDnidgh+eFzvO+2kEQTFJMrk31N2/AkmOb3+FQ4331Bj6H0
rtc/cj7b57hdJ2OCFWulCa72k7MfV6E6EnsWV7zo9oo5Lae0Oi5/dvQmEpQLciYz
iqvdCI6d4oK2rWLSq3FdbDh3kpX3ZrVXqrNHF0IeZk+4PmZvWUl7tl8uCI6Zecvg
9r33z4UygqoFGfig+DRxq+FOCehrB+jceI6xi/m74rTahDOd+RgAjFs2BdvAk22X
AASixY5S60I7HF5Xx1urbvtefZAJb66oQVz1UhIHqV00geqowjuFQ4oUE9GVKq+D
QrVdwZ1g1NnqXVcq61JxIcQvdkPvRDzUtka6TVBk8TlZ0pgZOT22QqnUxiX8Ljut
BlNCwAtLHokr2ZU2PORQmPTphLmXUxYcJfVRghLQz3P6IA2/oFV2NTmJzJ8FRcEP
IH8qUsamJPc4UAz57qxLrgADxFg7IBwx5Lfuxkh29xkaikmspgR8AeIZKyxOlCYO
3jfqyhAYJRz9jaoW50bwR39zHblPvpJaPB2XsXpONWR2BZ4CkHEQKJWonOuOHWmY
F12y47vRApzqxG4D4CfWSlma2Enm1B+nZ3RNudenTbhIy1MioYUxx5o7OKRyRQTa
GHXiYS0tnwR7v7CoHeNv1Chok0nZupLhZsNL/4MMhQnPab5Yf51ec4f1IFE7oMlK
58cRG0ZsUW4K3W86E+VoFhLhPKpQrqZN2YhHnN0wadW+OEkppBO+1PZzqQoQEg8V
wlPyN7NNdQAqkaGBT1dpJz7rXLsC/xSe7Lhi9b7qtcoWNbpTibSDMB0XCMQdeJOi
U2rkqMbaCk9pxKoUBJaVCrP2c0NKndwsrRuqoBC326hqz0hZIKpMQLHJDAkPg1zv
j0RueW9ak+ClhhptDZ87518LTV7RhhOChl3RuHW95TBVppPBUGfcqn/ct2wgw48M
wL0KLDlZTJppXiToLr9evJhUAH8mZ7BpcESnRU7mCxt4pCUIJQWAWNIljX2Pi+Ca
ILYd6vX8K8ycyIkkXocZb0ZSIAs0F7mhTJ/nObTV9PjxuaQnkDn6U4NMT1vbkJyR
m1hPjEzi0fPJpeOeDl4FdMaOvtk10UJrnA89sbIo2X0nHCoxWcI3IqrrKfxFbo4j
dhbPfxTs0QzR1z0NWkynMEIdLXaxfZATkeHK3QglAKc/lsE8/7oxAZZFsW/XBIgM
hDxftDWN9RHZ4si5MKutWTIZueAjyJFuhtEgFvqJBmv9ohvnsYzbbxYN1xJBb8DE
rlAOBpQ2bjMtQFlih005EhUF3vtz4p5JQfzQrwuJ65TLRap+XWIVpL/SbT8v5Mpo
GPFWwJYEP5rqysxkdQ7dUZUn4B1kR5+jZwFHbD8moFds4sa8/uzMWKfoKrTmTqvi
S868lIJ3JCdiBg7Eiu7Me6bqvLTjHE5bE37msoZKzX6J4CKBH+ebahwlaPWfb8eD
TfV3SWu1lBsVzw6MY9NaHVdQsGXgyoCeg1rmJ4A+eoMf2xfbyLW6pUdfKOrCA5lw
RVhutyJLmsJ/JpuYaE4OAzy3Sm9RzD+JzDtxw0ScL/+kkOLgKpp5S9M8KgsTtR4n
WimwDSLf5iElDbSWCqvCGYowKhHBMmcQg2tSBLGEQZ074sSE1f1xNjIMg5wylIUn
KS5ABOLs2S3uoX0xerFQY+ou/CiASrhoKO6ewr6qAwGJPBUmRyz2FzwxMtJGRdpx
FTSK74y8RWXTw+fWhRZGVnODrm0UKQh2OP7HfjX5ilD3VHC6VYQUIORWj8Bh+nLi
cUBWikAaAZWcy6umRE3Fc4Rzmv5P02gSd6nnV50lJ0eKBLM4Fjskfxzo0ycej6yx
fDbc4PNeM9G+FEoZtKx0qklWm4OwgG7P2YhrbS41bus1plno7jfAgc9aPmun0G6L
bm2LB/6uutgX5ZkA9VsBUF8c5fZO2E4ByghzXzgir+dyodhlfAzjKbj9u1QiQ4wD
8GC/L78Zls8zMQSYyRn1Mu/+aW92XrNVcFeYTKbfAG/8mYNl8KvEhvCNTarOKwWV
WfiLgNnlFdKnZKhjL3ox0NrgJF+j70eZ+FnOlTbgKClKKaopDvYz1vXF/ZxBvnc1
ng79oL0UzbfM5Heny5GrX35aCxgXh8axGxm5Axyitg6ORSoMtswS9IdLrxeNp3z3
o3vOZ8cFdpH959a97vS1fhcc5g35y87GQmYAFQhdhe77dhrIx7t7iTMaEchqZH5V
S8alpk1FAaVBwtm21EDlgH9FSR/egBT/Gp5uiz6C5dYzu42XO0kSPS4qN0kENjxA
L5HRI5IZWY/wnpP6TJUlzMWdPjRylRIU6p9n6DpEXh9UIg3/LC5Kos57a85RnDOp
+2WSgXcas3S+Z1MY5uQitGHeGd3Eupvg0EAqnd/6KYXDY3IbiW2qG+E+shIXqTHc
YV0QjDRbGwPSPDMxvuaeWoxcfPddI6wPppq00yYyzLtBl1HcSZWcHVpKo1U7NUTX
qhpJ7HxA72vEsYXWsS5umgnptDTJK6GYl8osF/Qa4uKb4m0ifhg+2yTtjMNEnXKa
tOwsg2y8jwNZIuVMCx3NdszcKoDVX2bj0tPVWXSwq15uKXh254LX1A/WG2T5+Y3o
KNKQWiIoCAXvrd5yp72KfvPUYBSoQOkkgZf9xuoBCUuKrIR2q418G5Ii4qh3AEUj
t0TuumppxOm7ay+xK76IiTX2puYf6Qyw3V7wNOnDgNovthH+6u6dQYTP2minrKnh
jgfR3zyLsginqJjlkBoJVKs+TTJEgiPSez2QLqD5o6d9ySt4ZYzavNZn1nau0oYj
ylCU0p3kRFVdHxuYJzaxZGWqdqE8reIeKErXVsbwGwCWaIXt3M6oMffPlofBRYy0
sm225Entg4HM/ArAJdrgz6ZuJdJ6M+IFbR7hNdcPaKpDss3Cu9hQTHJDU8drNZAo
KLJKikuEXK40QpElhJEAT5LRmwsAlqBXJYQGgy8RERTahLkUrZN7lwFLCBXHpgh6
cNig3qiWdZ9+xHOuyXAdBEp1A5qEn9dsJ1PQkceYzkU27vMIJ7QOQvPDSkIvNXHy
u3qkezRaMsd3VaxUSisLZLLQCBFjU4+GOv8aklzmE1kkBIgBPPQjzKyrTidhYSr3
+3jaVs1K6KUEGFCGs5IvFKvSixsjR8LiZbBOtEC9LBCPpD48nwXZ2p48ZNwFNpAO
7eQxNNZc/BLivuu7G3HcNVLujy67Zx55EGw7nGehJSOjYi6S2BqauUsDBWOh80OK
1Sdz8S3lLgT0oIq4/E1bF0dgJdLBFFYc3+N6IEfAeRuB4WgW7avFbmjd1/UXF3pA
/D5WeY78LB7McooL237bQJNMmT0XevF3jqYcNy9VPUFUjOscx5Wd3vPpimrN2YfR
7MsnGl061c3+U7lnjb/SKYB5XPy+HQ+2EtjERn6cU/dl3ZuHB7f6/O7w6f9Vw59F
ZotCy4Ws4hndBfa+xVT3WVAJ/aIaDE+Nu1gngFhrkzy7I/myyRHn8OCq3OpxgIcQ
FjYNOuOAr+DfmtSmGCzW/jLaNCwqUB4JHIRDvDCxN/ljjxEMTk8+DFpzcUyTPp8J
tYeE4AtJohFesXNincFNC5FZz85rRumtL+ud2TaO+nsBrbG/gn0wHDKsnF4WL0uH
2vJA9ccrfknpEiE4uGRlo3z0iLnar6JkT7G+0g5+4TWPa9WT1TDStSUm8JOWG6AB
6GBB6ARazFoMedMgKdz3yAwJBdVfGCFY4HHrkzpcCZgUFYXKNaZqul0lUf4zcjBr
EZ8hrJglxL5Z2QEcBYYe+d67P6bgKApWXRQNYoJ4kET+IDZTj74xj2YvxcBBp/ll
ucfM0ETRGwY8Qx0C5I+1ziWh617cq8Zy1Bc6LN3wLzKV9xP1PzNYxqvXh70yDV/Z
/Zy+UuRhPTBFhzG682foSP6CV7SjPK/V5+dNE6lYdR4UFXIZpyqVRwa/2M1gttjp
YLAlvlkWA0myJIoBIxu+Zzh1DXXRL7Xgu41KAl6KroQwCLiC1yCT3ojN3khfpaPL
+P/5XeMn4ylL16zj+Q5x250Sp5SaMS0WFRgOvBQYfrbDxag7hjxO2KANDfX0mU5H
Z0zA3bBp1WgdIcYCo8PQnD9K7QjnBfKS4h3haGBVghr8D/HH1ThsTkY8HIpRvHfa
JQfSkCoEi2YRHWlbA2gFbMMEYX3GpOzE64+ry8nX34n2qkGVcdSTBO2qZ0dtlggU
d1AlSVlaGnw1nI44cyJoNHmds9MO5vBCr6QoGJ2gK2cvdnyzFDp/mVwBNcV8TMOf
A0XksDZyVErb3yGcf1Rb+zA/2TELOC2EA9ZrUQw13IR45+lMgmb8Cg2CgysDmN3p
Jxi+uG40YbxqegUd0WI5CdeFLrhV5Z4TNAuvupPMGKleH4xgj2MgWJnxf8CpGmZd
ijgtkhCIfLCZsNxNj9RZHIUSYy3hulr84vkhsIsJSEYPtytSWtRFUKDdbYF3gdHK
8+/CH18tqUkhhMnXalKgVGovheasdEmu9Ws7f6ObN70tBxFV6jEGlNTAqVVwtJ3p
utjyk/AgDBLORnganx1gJkYIwM2Ia15JTeSM5YihkX7MahZbS3Gd5ZazBXgI803h
p8EpVuz4h92wmantivN9b4gOT20E6e9f/uh7JLIC1YGKXXJew3rmJanKpRKjcfxk
bllieawHFdOJc8Xr/2hggQfdUI0ruW0TtVdkWiaKfegU6IjSgUyTK+ZTnbPrr7sb
GTlO+tvK+wk2L+tXybpdh08NR+nMRMJt6rupJaaDt0OVxOf/L2JdA6cBcIS8i6uP
8zF5+WJYgL0tM0T6iHBe2kd0teQO5WoCBu2BQA/GvEOvixOKlJisRSqB40g8AQba
94WgKktdCkLVwNPvYSGhYnwhhWvhZ8L42LLZa85ObYCJzL1PIfAduG1Q3o8PtTqB
6mJAnubp2cBUJ0HP1nuZpOtm6Mk5kMIboA3nh2Ya0HdTHqB6L8IBbiH81aGwby+I
UWMX6SBO6AAAdx+7qeY23AmitU0gzhFx7jOwtMiYXlNO+JhiNFGfycjfO08arHYI
sqV2h8JlJ9HNvTHWnHU1JCKcSdxGdVI0yJHiHvo4jdo7tgC7iM0+1Pweea1SQ5Uy
rDLUns3yCMMtTW4BvJ4Ks7EaNYZZWO0Bh+ub68p6dVigCT30AmmiFcwqY5fgHXSe
4FK9qatUGHgU4iD7y7torOnaRS60MBxtMMBYAzKjNi/roi1gtd6RnFsvROsswI5J
An3Nzgvk10Gvx4d5SpysIGu+02uJ7Z/gMpy+c4RlxPfESR+baK/8Zt/Ve2GwaocC
mhQig8n0JgmnwXGfr4FTSvLKCDpmkaYl8hgx3kNbWc6ZW8bckd5F2x9EzFMWvYYh
Usr8K6nJcp3rlaL5e3zTTkht0v8EFzLtexN6L3fOWxtm78RDR4A0oItom95vgpmG
EcPj6XM21/xiNXNR5/GppD2A+3sR73t2LBJj2TgV5SnmSgKbF3AjBwHuEjpdV4Ea
QOmiaK4TPzzFndjQvzKeBGEwMRk+IMnkSo8xpgUKAtVsgc839DHIMs/vjXOf6aZg
sUa4IH4Rb5f8W2Kpo6yKuY5XaOQB1u20jeVUvwyBSp/CN8FU+TAAUjv/9g9nQiDQ
ibctUJZXMEBr8DBLoeZMSIRBXu1+wgWN+ThnThDVENptoh8hBqK+FJduh96rmI72
OJw4iSpIGvJWO1+5U+AT/14k/lsx8oT1uPvn3UwdzxMtBhxTe5OS4QtsrvyxNrDh
6WVBSA7XXt0f5+APzMxE+qBa5jcevXVDvA+IokCI5PUlPH6jdAz1g6y2dfSfbJSv
pJwhiNj3U6o+y8oO4By5WoEYZ/7Ed7z4oTCsToh+Dt2qQYWEnSxYS21hV8cRV0XM
GgELCW7L2eBb3FBECqDdeoFZ9XP73gToflR5joaB9MgGro/amY5OeHa06k+6gK2Y
JGhkN9P+Jiwl81hgAyD4G5UpY1HPRcekejFNFFIHXxalxZraWt6yZ7h4kCsa+7J6
mH1tifAqiVqp355QE9f+L6myPqOB+0UOkzxkteJ6Zk2AHrAuAIdhtRuc3ITIXxux
FGBQqDV1YovEfct6jGqDsurzpmFGgzoSlfscXpVqLnXYWuwEIw75oz3fzMfL43FA
QIuuUkLllvXBVKBMf1NH97Mf2DvIzgnC8/JQTrbwxLwUu0g42MTumLeaM6M0iBj2
LsNIqHspc0BZksmjqUfXlRl8lavvKZSEOHSq6D+soTK7YTTfkZg5BP/LfbukRhb3
LorYw9OK+WHnamPdazL626WISZ/Y6sE7izfh2kpyrGmaHHp7fEj8y0p7xSjP67Nw
NVawqIZJtyfDwE/eo//N94pK8aeajaaayav3M3fTDUeOvF0z6vi3P7ZfxJ2C4TwJ
YYqf5+R7wsIMunijPv9BG9pzlZMiPlkURUyu2T431bnBCPw1eUi2r16n7xUnkWRZ
bH4WDAqZGKc6qzRRxuvMnzh26B3PxJB9ViALqq2LZcnJm3MY9a0Y50BubgpI1D+q
N+7f86IV0GAN49rmLArwHlpAncDY+97c0Qf7zl74PlpXvkPLEp+KQE8DsXQr6cA/
ZLK7iJor6mjSNOxy/Ij06292u2UhcNvxOo+OxHimzAPYCpWLMtOEEZ5+9k56ppGc
6WXXPD2DN5LF79Jz5NooJFx3cuaBgzkORi53bKdqv7Jw7Lj6qRK26b2p6RuDTC47
R5+r+wfsTXH5N0SYEGp5hwZuSoqTUfzvak/UvkhluX6dZcB0Xphj/Az9SuqxGZ1O
KXNXdDY65jUNi5ZxuKsApi3bmMBf8yyenPTdqVDm4etX6fG73tcjqD2BU3731lv4
gHtZCtekaPTcTvJc+k2dyO6fgp2A1F2YG/wyVWqbsT4n6sVq7tdkulOVyCvayRdU
x8S06aAoc3iBmKiwiinFv7Z55qKPwQjGThw3s4MCvnsm7pAwK4elXxikXmywLPSR
OXAQFtIW3NZDYSFNBhCVWVV0QaHLTuyIVtPgI46x1TLytqRxvKeA6k0gxRr/mfJC
OAPWYJHVFwl/gVKUtUQimXPI0LG43QGWYSUM39VSde/KSb+rg5gSGRyq0OMad22p
ANL/4Dc49RF6wojcW8cVGFpMxRObdVTbLvHN0fMKOKBNAdWlLsQaGatrbwKq9UY/
PMjaUiU1TYhSYsqVrzpyI4UdXp7M32rIjEkSHHEStCEwVXU9xqhKbk8N55vA2qAL
hBeZBvt2YocSEJneNRbWyLzQKfuJ7/VgcvtydxClpzdt4rslctzNooOgywwjuQDG
y2ItABPXnpu4QqyBtyM7Nddm1slBWt3f+KsrEpQ5Z6q0LBvcwo3fjAUwjmKQyokz
ZO0MKxH8Qyc9LkgY5yb6mRU1djoKGRMMcc5FjjdtxxVO8NIoOFWuBTsTOwrEOo34
tPgFD+zybqWt8fwRGViCFRT3586dNAqm/FtsJS3yhb9oB3iF7rRItU9gtHsGhDYD
/T30V9OO4QdK7A7iu0viHbE5ZHKfu5Dd1xv/3brXdEQT+Pqhiy/gZdGNrm8bFnf7
RhV8V62X8DPOM+fobLwtIdgvvDxB3ZLfjitbqI27+PDODWNMSiZf3bD6AO5EBw3S
SgWmJRyw5mi0q5c+55eepGoWXSdyHr93OBXtgeFDmnm3WhQInoegUJG73m5Z7SO8
cxjUY9F4RYAlcXlBnaaUOYD5Xm0Mc0XU63kttJ1rg3/+9DnJ/RD1xWOTw6M6sbJ7
uinYXYPeOMhduPObECNs+emrRB3+vKT5lheb7fN7iUL/0JF0T/aS0e78CttjEw1N
aWEgYm2nprVeqdZelgkw0kNfcrpEHPSaSB0EcWyyQypYtG2OKp6efSeDFH13DzQw
AE4o8jTNjBJc2iX0awaAwb5+YeEJhX2xX9DVIq0n8TPxGbef765LnHyykHaIoIti
q3hhitp4LSAMm6vpL8Subo3SC2l2HGig7PJaomcRU5lIXmJCop/de7UtU8b4Zbkp
wYomtEmQOmW35MJIuBeC4a/18nzFuYRxe6h5UBIa4//VRPsMohSRbOuXkSJHTo7y
l/amDck9PH2TTJBfxuxk86HJEKcuAMK+8P+O1fQXuG8KlajIqXpWmcI3/AU8fSi3
CmbQJAp396eS5tdigOar7WrCEb01466r9M/zNU3hNPys8t73ReEO8FQsj3vowz/K
9bVlZ4ankFbGnqcJDrLR7Bhl7yuFOkaB6zG+uiJGROdAaKvPjVyZFhQycJH51b5m
rsl9QaFqIQgOYDEJgIS6ffhn7/NzePPwJm9IxRDW5rmh05blnS/hxoe0niBGr+7j
CwvKmF45T22CXhS5RTBER/QYS0SmUAUNWKucrN4jAxPyjMWtfQFiY1FOPaDGpysd
6xVMr/O5SCfJLjjivCZACn1xaZqbdgPVnBxLSNyfuyNq/6x50xHAHdKAwzAnqjrD
1XHd4Pxb+lNiMmlVamNCex6xX5NeNfhSEsVdf/doLhEmTJMs5AZQo6MspmnpxM7R
VO41vmtc3rmeHw7FzLBZTgg/DfPY81BtYllJISb4iSVDHRtjTp85lkDzUIZK464+
ta9Zz5V7wD/GS9mjTHYO9oBXh3JXXPZzGTFV4ldy0t7FgOUgR+0BhKrvYukB81T7
wxx8yS/zsWKSoBHujoXUxnmrRx9g8UE+iz/vJFLkuHYLQbySCteLBIY5ZxlbqJGN
c1b6Mqp4jy4zu2M3cokhp130eSfpVjEp18QMJbYxKhR7pEpo2Df1/f9vfRduzJ+4
lsecvDKrzAw0ZkFJNxxIzLnhbZjfxmrstpHimrO7YtLyoEXLO3eZ3mFRUbkmGBvp
M+kbE26ey74ysFQxroU/IGEbKUDZ7/XcaW2Bz/Vqe7rckZbZhbeTfZ45tyF5KwM2
u+s1tqCGSTOWHpsKtvsYF4z7ippRlUmKn8Pdag2OPM7mKLpabFgCq+JRBtgYZQ/j
b/xkdeswrCn8NEA1jdTk1u6z4Db3sALsm18x3/i+CNq0rA2bpvLUC6KTmYubHOCM
cb8heQLlTGxEoGN93eErtymxI//ogq0+c6CCfnQiPLt17OEKgjrq416KQdp5kQZw
+VGUlJ4Yjyg0p0qhyOYG25hgGK+CV9MVdjWI4o5ZtuHQaNTgsQdacBetDPPWPjsy
3SWNkc9tXB1CGBMESkR7Hf7CGOR6Zvvrdbzy1i++Wxn4Ds1jra1s9VcqtWp3vgMG
XrmdZzvcB0RiSlpij9zscbFECaiN9z1hF7hvcsm4Tl8lAGw+N3eRhBeBTo7SwLbQ
a0NftzQG5u4gZ9c91fUH31aEiGnS/PU1LmCtMai9O5Abq7HJLeN8k2hK02PJorP0
tABuWGzxIPOiLS3NurgWfvSmFmrvVQUi84hsS93t1CY0ucRxCPd9OleAjHdfRRpL
2eryo9A3xxVzeaBV65j/rg6AtjWEBteBwgbxiIOAnvXqrsbPSdhdL7XVpr2QbUxd
VZdwq/Ka8/LxbTajj5U68FF9qr8chpuLtUhhmwy2YyQISxAdp5E3v/1mEGp5+zh/
nwugAAcroWJdNJ3214hkEa8+EIZGuX7pXUjako6Wvizn06MkT8znF4Xr8d/TVhiv
6oFz6jZhrIUgo8iAE3bxnXUPmz/ed/oo0ffKfYQqOHZiIvupvDi08H0upTJQRSse
Uh6DpG4yYaurNP7LTt74+UV1bQuq71XjanBbRP6zYrjvVk+Nccci6aQJsfC0jI7V
pbdOERX0hXA7w3aO6FWCm77QOtaevRQ7usXZSF672yVHM10F68/4n8TBxaCauVvs
FXFV7VtPIJ9Csevi6/yMvfPf9+35pNsc6Bmz/Dby/lhZKHJovT2ZoIu/kP4OPuaa
SMXSmbylIqF376a57vX4kHtztxtKTLr4ZoqtZhCLXyA86SDbFBgTxhkERqJxaQV9
eTubV8ZJA1hq1WybRTh/oonllwFVgViZqQSHzLLGFRS2czAaL31iCnHjlmbUwnpK
/srSBcQ6zQ+W0uIPx7BLbHBfeGqrvjiSDQ0Z+rgRllosLp7OTz9Xt2sqMXkr/99O
BmHabjdcBwBGlLYIGJqwV4uFoK1diXU+5cHIEncQA2KjkxyniHWsk5iRp0QQGsOP
FqtGeqM+J/EqbT4GwbUMOw1qaAbvUyg8m0BmI8v/gBvxRWBFtjlHog8B+RTPeoEk
X1F6tTLexVpnajhedos4aDE5z+DQNjtCkOaMMEvF0Pojl4LQIcvftIEGtfoU3XLD
b5gJUu/yZxSVyXDZ53vJr9Xau0x6LD4k8aTXaxOXFV3PI0ESYiX22VapHe03kHHy
FSo2ZHu4JS4qGmjiXDG3xzGNtgriVaczmYr/cbp+1vxozT0FDB9Dhd0ThOVtHSw2
cvjYiZ4XmAJolSa7dkx4yiuwa2vUo9RdeyfwT8H3EQwDouGfvmEi6RPNRRDJ9arE
J6IQpW8T+CP4LhLbyTHt8n4OcgG3xyLzFz33LOEvr32ebvxI/yWw8MA7c64O0Ilz
80dcynrOJqqCnjDY8d09fvp0npDSPuslZoz0KhbEwozZs7psWuR2x++sv6eCFFkB
W7rt46gmLP7poJOHgNWlhQFC3tf862aY5FzyOT8c6vv+IZeIJ5by4HFM+mRQrwzt
a/B6C6eqS4Vv4PcA3Xl4XImkch8vjs4o9kt7xj4nUlm52MDZ7vX5FEbLL99Jvmu5
AHlJlOw9dBdPaXA9r3K6rVvekzybUZcNalWUSQrr7W0fML4iM3IjcfHapzOd71wV
MpbqeBe5bLntjuRlXxeeLxoJY+06qtDbZsaUDyYPy1k58O/KD9yjtx0qR+JhI+et
iKPH5sJbJ2k+sMN/9k9qw/kQSZVwwwUvoBC1QrwE1wnmVlQuUdMEcFDuItc2YX2c
KXE2jTIcTjqrsTxOYPvqcgzrawflSvIPG54RHzSWmFqhDS0qhQDXXPsS5eLiGdNw
mns2Copd0f8H7qUa4A8nufFhbamG1jCe27C2nMi+AkhDy4DMMayjXhNmu3gSmRC9
hjqFRGvTbsElLHGMkWfu/BtJtmwRmLmHwc/MV1hLU9LmS+JfLvqkUjzzl+2+Mx04
ZUND5i0BFt4XCLEoPtyAGDh/28IXIdieYG6ENc1Y4VpsCL2WQABs7GG5YsBe6ydC
otKezFggbWW+EJHGyue5Mz/m9OnXFNRfXtTLepuad8JoYP4kJHbCquG4N1vbVnOI
XnH8T9s8oN6j6F5BlfG7H1dSWm3ewKrlGKO3htmyqn+yW9RiTlcKePfzxVYFvK6V
O7ytCNF1Ct15cdVlorZRWMut/3agfqHlbNU+s7c46sHfnyDXMSNXZgbLNuahTghw
JldQy6VUgV/VEUDK6NXMW8TqrN4BuVqJwgv+r6SzK79Ja6vnzqva8SlM+2A478nq
WZ/BUA8Hew9N21iZh6mjun52VBGaDuCp1elNR7MRZ2RmVtcUX24eUX2jg/AGa/br
yoqAFT4lgIDtAn+T5M9wWKDeS/wrugqf0GXF231EVk78BOM1+fAIAsOaRvFE3f7f
NcqiMM7A0C35ZGsEDamqARW9XTGRjxYZYEK5waHLnTM1BMc9qU8ptre3wIP57IiW
MRxIq6FFrvL1rCLy2SqlJ/SkBCZs/7hEnOmtPI9e+LEcoNsp0vYR8C1en4DMy5g+
oT8Wqy/l7vBeOpsmedNJ14ckgwE5txJgPAu7CRqznBNviZcWl+fU8wL6sfpc25yw
YZnplfTSeV+8ruOxOL7MYlgceLBYOM85jgo78IrPL2yHfOZpbhDT6sdRpMtCWq3g
nuhK+1C/cYPMJCl4yUTJ9IbYJuEO/VrMJruexigG2NyRBe8Syma9OLNbKprV3/3I
/Z2wnsdgofWDJunZrqKJ4rhJEfNz6C8evSykOjCN7nhKARoJbat4U8m+SYCks76m
AfssTaETIETKfv0PI3sqEpuWN/6hc8y0eprx7wVRM8UalyEhb3knovzzU+GxcMn3
gXTXzXqp3530AsVjc0fUnC5WK//TjhOY6/fTN4YdByBJCvMdmhU1Ac6DbXE8RAbD
WoyJCuVgoQh187AWVg5lMr5NmLcRSgbM4vTqLBdexR7RxiceOK17+bIhUmkJGfQX
xFPfqRxoGdZ9xy8FexTCmHio7zguz81B/9MLvdNI6sJtSJncgCB61FD5lvDhJYoz
myvn+jqf5lEwm3FAzmul4BXBLC9pW5onU308uF4i7km/fwDFoVDOC9LaIr9opOoe
bTnH4SWSfqrAs4BO5D9c5dvRcL1uKKb+0KT0KS4QlEmH8YgQUa2UpkuFeVZcqM61
4czwfR+Rvfaxh6Q01oAKmDeYWERFnTViYCx8YiQGz81T4ntE7p1emrxh/NIEUITx
wYOM0WAFxvzy8jiKQ2qhodhTUogmLKiOgmD2QziVikwYzmz9Sz5ilau9qPZomIuu
N4rscIhbAIUBB1sCBSyXz+ub6dXec49POqZfQYhtu82TjyAxHEYA6fL/wzzNVDx5
pYDBIxhhAZ3VRduDAC29UQrnLBkL3oKDr3JnmxC0tnfJrvPxqwtiBrkQWuFwMzVX
k9gEahtFo2kUAyqn5RcmOLZiqSMHfkoOdrW1EQVlCIJf5IeeZr6wkSArdmNRVFD4
r58JRTu+vZEOw9533Dtjpxo22ci4AvU6C6gGHw17sX24vn3yf3QZ47oFGdu4gjpk
XtAIp4QiGjOzzk8v1yckPUxvt7hgNm74wBmsBsRXc7JyCSJRdK6Qcr5XHpL3oquc
FWEh8nu5phLkqxAC+LAfuU0TAJikIG9VxBL2/BihztzQQqaEy+0LHmwLoXwPmXth
qJca2+p3kdNNscT5JExkrcQRSkYIGT6owzUxMZ/c1Gz3Seicx6xyp6RkNoEnvTw2
/y8xnLZLsI7L1Ax4q5559+Ane5Tmv/1nMWwxvImYL8kfjc5xbC9YjwHtxM5RXaXd
+wBHTrqH6n14f40sYWMx1CMpKiLma87ugh6bHo2NkEBr5ayTUkOlZMqz3qqw14XO
Mm0lV80vFljT4MhLC55SR7fw9UkHhsXcsQMlPzlgrDR9+UUGB8nlXuKygjNMSeDd
1Mkh3hTYyNevLfuWp4gqB8vbUI3ZjWNnnGbU/c/lEOlApl4DYe1heRsBaueULLGW
J8QPjmFLnc2aMDoo20H/Z0+UKprxrAfB23CcLX1HSP46FrJDy4wJKa0C7UkEj4HW
/RHfqn95O6Q5VFSYYM8PVEuAUv8BFtls3Pq8W35dAoQ5C1RJi92ISYgUNMYqiKSt
FKEtSz9Jk0NuUm5uVAZvowTjNi2j77U+/Ld4tsu9Fja0sLsuCWDu6Jcydq03lgLC
1AUBtAETz6q9yi0EVXh9xVOZWJ3UGjIGyA5J84HMPrLhaiqDUCoXKhOr2hLi3goE
HE/zPuYip1iGW7kZu1iBe8RKDoGHoW+No6isccj8VzolfkJPYfDQPIJ0GiuduQsN
C05RgNStIrxZmKoyqnvG/3XFRWazCH7R4bt9wgkjsEZ61lRTB8pKEMAamp8to43/
MLxgw5U2jGXW8S0vD9zs9guywqEZGj0Tkj8pSuP9bug5HD/8thlBr4oCkBFJxO90
tjDO1z1o7+aaJmj2grDkp0CBluBNKhsUPMJ8TmD9T8eD7s1h6KTv6BR1JgGP/03k
ZaDI3/dapK7OZtfZnl69p/k8XODy9lXSf9xuWMYSYKZk7gRIs3xlTIPhZ9XisjTv
J2L81EcRQ4uLDThgx6iYRYyCc4d3+U9idgVRGdnSh+SqJwf/jhFJKd/ydov5Te00
CZthK9Ox0RbjN58zsJ+QpnH/sFZ2Zb2LaJdG4WuaOSryTOPplKNQr6k1LjgG0e6L
zRjjK45ZsmpGJGIGLFLd7dEDGo0eqFSPHN55chcD40b8jZxbxk6/do+eEczgwLnN
H51y58fVv3T1iMPdIYbWulp4pfA/L/J5EWzI7gJkl6RqE5H03qzUh5t30xa8yrmV
kJ9x047ha7vKHOt7GnnJNrIRRO4EJiQk7HQ7RoT9Hu/9XrpbU2l5G1z4QVUdMtyv
TdFfV8+MtidY/hD1y+ZCKNlUM+nHtTa/i1YhJXC3ul8Fht17+Eyy1WpePuloCorP
t93OiefCT/gZY5a5S4AUacS4ejS6BBIKvtzqO7+3AinmaIzhL3gKVwEu+H4sbzTe
Nd+9+8T6v5N2OuwIZ+p6MbFqTwbVvBSWttiv6JMErWT61/cX4l+queo3xMYatys4
77IQ9ZbxJjwd+rZ7vGM98hMG5J4yA3XZ5FcNYIz3JjJCOLmdNVMMcDgmt5tpWmpt
aHaumHx64itwJcCHk8HHdjMkHtH3nPLbGUVY+Wftr6FET3LXmEZTXkL5Q6UQtbI2
oroYiPDyaBMO1UqmTxJFv+h9tIUjw+rTO4e8mpVRWjYD/lV1gPlTXabNRXlipMgY
fPh4YUEkDzNMaHgwD863OFIRb1AlKfOcxXh9aAIwspmWNAVMq4/CC9cvvbJdH2cT
tdjyTiP8Dvtw8DJTzsO5Ve9P2qIkvgXN5Ff0AnAfk471wzg/MZ3rUiJ0r8RLTYzE
d8Q6ejHZbMUUojDEzxiINkJ4MD1m+lYqGq3SQ5oTqVj/j8S4+/n0Ix3Ygtf6PBsB
1IrKGAT1Qo8cm6m/gEGE34xw4icwNwChXbqfwBekCsTAZoIIIDmNu+DTpgLkI00B
IuNaYsNxsTBcICJvTQJwrZHbCRrFhvXcNIrCReH5wLQu8oEJHsu5mZ+jMUSqR9PK
fnhoRXYzlNnx5z58rvtoxn8KuMu/jJAux5pzyKX2aSvGB1OxAmA3Lywk7MYNaJzX
Y/1GEDqt4TsQTXvVGbKw5dVVQu3FhOodql9zmTDWXLn2RmVeAgslN0qpkjHmon/z
0TFlkpqMXQF7cBeCgyoZdLPdmKxS31pjMWgcIOTes5rB9DsRs+1PaMr4Dm552hIo
9z5uw578A03hW6CHAnM5UIe7N+KTB+H4/FO6/PzSRjaqEnVs6kwBUE8XEp/3lUvX
am1pKM4T5yg07ZyyH0k/E7DoHtt7cijqGhGQT5D/oy8/6wSI2QbWzOes5MLJ/hN2
0ZWrKFpeNPjX6RZ8ugRuI+Yile277iskEqxBhi3IhsbgYb29ZUXI3ZaSBaaVZZhD
p6ou1OCVyGUe4oBd995eh9Kf564K/HRxryL3PrO4sL4IKEfLCGbRQ4YkYn5JZ0/V
TgrVgeYr7m1ug+BRosEyFWKA421dK2eVfecUaObboOeYKaVO0U6rCzVAXdsHZFtN
tyH3lVXPdAiZt1hf96l0powYWCZaPi5kVPV/65sUfXaxdqzA0QOGd4S7eEbE/V/r
kXJGPbzU+OrmFG9s89VGUkv+GTTK3TeoZnp2KksUtRqfIAxvvd9qhCPlSiSdYmxs
Xx9tx1RZ8yNYKHrFNUq8yWzzL17SSQFcnOYhWUG8+GQKc2l09oEZjHzhWR9rzxXu
yIY0F4uxIr9Pq7QgYdm0bQmB84YIrtr4+gibrdGm7gFMZkHcoLV8+WDJgPuux2eT
EQ2MswVnLgvw+WdfOtQRHWfiPulGGY44KrX4FhiZi+g2BQoQVelgpG6kQgl935Pv
9B2YAarwYDooOuXkGbAeRKWm/R4+uaELS7S5mf0WceGAaUaSaDnf9cvHYfMHblfM
m6Ehq/yfFMguoqjGyJzOK0CPjxBYoUg4Zwgcu0hoWngAa3pcoFMwjs2i/rZt9tre
vBLeiR3tUjyqq2V55vDeqw0oENqFbKbzkH9wVRWvoVo8EJUxfDtjXWx1Lt5bJ8i9
VNdJQ8itk90e5XSaJ7id4YpmRV4L98RaxsK0PMV1AdTVNKYWf4osJBVlnnViflbC
e3zvud2BEP8nUOCa/G1WSKXxT3wJHjf5/oVeyWyp3WlL9Pi7bTRr5nO7akrc5HhQ
v5jZSIaE8sXrio5vSLBhUWboWDf0m3lwiTCYInDs7ytWhpSaolOV2c93cDXh+S3P
QUq0cGwRApdojS/XxaRpNbARCicyU/KcDzkiT/3e+3uxNWYTOMjAubno703+B6zT
D6PaZh/fYR6lPDbmH4nBoZaDnC0CYfy7CZBQDRMcgWs/PlDVtGtciddfpXoE89Vb
XIWuDLsrZCuu51OcFGlCQu74LQqVzkfVELEUelVn8P/trVMulqin2/P681n0Xzty
gSMbG6EoMea8NIddOV9XCITK28rxuNqEwO7Zzacg4wx+Ob6v+Sl8hNr4kUG5f/W8
cxQ9Zay1JG81hBcDLOx6aPFVYXIsp1ybwUcm7b01elAVCuMs/QIRFgCeh8uRRxsX
f8oT+0tuYKzBM0Lm1OwTPaMJwIYJsTdKFjMzO+sXNOVjb8lLSPDhBAzGssUy7DkT
QsS7OO1yRkgCwzUFFg8UwQQQ9BV3PBpFUCudKEflGHI1wMl4zqGtlQMv1yAHJLg8
jBCuZ/NPp/K6jzfTaDQmvRb7Vo6xXOwRExYXL4gqyhwNoNeJdVnt6zol8wFKqZI2
QPYLMg6H9Qu4x1ky62nOhyRWbEcsqxzZvrDyCxdW4anl6L+OI56DwPgvYT2A+tP5
EzZ9/GSl97ScKwSqBIom7NIYwY0Q/32MuJ7LyiJ7msmjlLRmh8WydDTjE/o789V5
wxCQ5156Nqg45WTw/AeQNB0WTcJDTiofNEIiqorsVsAa1sniqvTTf5+qIseLDrYn
WwJyKn/sNp3mpRy7C/elUcSyW8f8Z5I+fO84OyRIOWgARwFQ20lnFX+lTowWDuAL
xhJhESfYWjQCUg8y5lsBXhxyB5xqlzAekGxpqp42ICObHRzP+OPGDPKXsxns3y3W
oWqPXDc5c9JnxADCZXdC38KmJGDrSK3TnPSXHjCJu70iab9O5iy2q5Pf6yzqCwa4
DSgU+iSCZ6LcHWGqfDPmwYuYmn0I6urvKg5oqdevELgUENk2GxhIEJbppVv/ew4H
ANV7zzDnKr1VVLOuf8TXDlDQoSHNSqudD2QE6OZKL4eASSQ4FAQRR3z7c6QEr8O3
3W9wlL/i8230B90SS1nte8y7C2zKYjbKDPbi3Re36if9/vDqnh+nCFoM+ytU71rE
sD0y+rqNOJb7twHkZkDIElCYoMNYuesYzyCPeCpIE6ijCy3RntoWvOA3+OzWJBgt
M8pxwsIz5BC8Nsmi2SR1HGBk+QWTlJQ+LbSDAc9oin8dsSX4YutxtloSoE+UhTGa
Z3KbOYFN+9q/r/kHHbqek9g+qoF4svTAQBOoQnfUiC0jIrazdlcJCiAR+mnfoOQo
Vuq3iSb3Qz+ifUwQz1TyP73cAGNhagUIVpNPHY2cYyrW/MMTF3X7gED4LWVdc/NB
DUz431byktruP2rfl2t2lQQkOzlUq26zgOi1royzAY21sttxbCI4toWhd/RungjC
5fZlz9YDcPbWrU0YYSEPGa2kAi/64+GFSnyOK7NmLa7vo3R7pQewqKWqjtjs1/Qo
XZjnoCNMyNrVur8WHTROHsL6XmrQWUIt5eDId7M3MiuDa8pVbub6kDWOZOSC5nrV
Oh5j4QhwpXLw6+B7iFD0kCQH6Mdz8JvaBPCAW7friOlr+Ptw97YKK0ajzL3nMl2S
WEJiFx54S2XB8CII39SBegWQUlSUXZzZOXXtggcAbep+QqemxL+2KY0yu2nNefPx
JPoWhgG7qvtRRJUA3GLs9frEu0aO7V7jZiPLAVXFaE4AKaw/hLi51U+gbSLFTrIJ
6ObCQe+J4aEAGdsbAEjdVtEFGufJgH3CGqqw5P/tAaaEYh6PpvQj3BBOVqZEkmWw
R1tVRV7VQfDgacjirnH1JRMCbL0SHxxTwqY+Hnh5TreRNIZjnIwmFmjC14OU/bCX
gnEfjGZJlWGQv7AZ7T9hjT0Cc1htwdaDyO5/ze9K8YFvuk4ElFC0RQ1kPkacAXLF
KqeVtdGxf4anJfssm41/N5hYxngCc82OnV37Xme45zlmyb3V0GKuPmMRXZJdYdKg
4NnDgYMyTOmSa0KYh1+esbn4Aex6M5fU5OjIGX0oli8ubQDknhbc6U0IAMDMrD4o
N9iyE7cKGE48Nkzeboo7rcbDs9UOPW6WOrVxaLTs+XDb5uKeKvWKRjrirItU21EC
7hmDKGRA7FbE8bbVKEu2/ip5DKmVB+jgebAtzQMo0ujmLLrZdCdITBYlCsBfDu2p
svrVd4hzkOuxz5rs0pWS2HKrTwefk+bFr9ZKYmZPVsH8hsRW/yLPMch5puGElLP6
El+N+KuUTzJPEEIcoQaxWy5/f8FDXrqsTvmmEW+k8/jAt1QVmdETPs4xDVVCd8zc
tivfSk1kAeH0lZzOZ8eylrcdZKG5Qmx9S3Th5eHkc8pozk2wTdkMl+OD6N+ihVcC
mB14TH2h9dk8IJdwJeHJ/mdagdc9ceGna8d7BqyS9TzgyMDEWpdBLtTPKxP1Htfo
3TcJ9sqspzIXZcBOUhJljYWIV2luC6mmBeGEAtdK1ViIV6R1USbfjdYXL0Aa3jzF
tPLl9lXjhFZwwGFsJjBIfyJaeaPb2hBtaf4u/9oTUxAGNTuk+hj6BAjogSQv83A5
qkigH8Qi+USsvQrKIgorcFmkuaxKXfmFzafBSJDRE4orFYxwBJvdVQfVEphnl7s8
Cu9ZUkgbdCHGr8dTcf6oa8yT5YO138UlLXJaLsLjITcKwjJP6Cn+AvTtdspn8sTL
dnYS7MfgeqM8zR6rs3XSAlIP42JVgUIdcNdLvfj7hi5SatDPD59itu8T71x7I0Ju
oFknBkle8pO+vEPx5dVfJ8PIZ77lF9MHWexN9NAdVqN8gZGlW93jFLsLtQXT3kX/
ICyWWNmdeWsHFO7Mx/5L8znY5EUcfNGQElPbHqbfku1EwXiJ1LKThdJvQk2IZp4p
MrW4t05rDSxDGgkv1s5rj/Amh+jX04Bq6zWOYMTm4T1O7r1tl7Radu76RBhnqlry
NU3ZMEafoac5tMWxpBAWOZZ1t/bTeheSngW2VGvbT7fDkhgVRAXIK5l03v/590s1
ZbZ3IGEd6tQWwVm0JYbbnaXZU46p2YcuDekr63sPov9n55HQDFTgkzvJ8H2DFuuF
03T7CRhMLe4BCtF2EyYCk+l3eZM57t9f4XLn4iW4Z71t7z4pmdPeF9vdh+BA4yWB
rRjWNTGmjR4Tcqu96nu5ida2jg94EIXnZDGxGv7/BOsrnbshuBB4zNUM0iQ2o3bp
mxkyTyJBeR1XSGwfJdUp+/87aM4rYUWxLGvO96evKUZUDTQawcflbFjhqWruPGKG
io3Gx2osZPsiQzARB/O5cbJSmTb3rOrLhyJgFv5/xHtcmJiUhjj+X5wVaLwL9klk
80pJkduJl0uKERv34CNBup7Cpxr8gwANEYXA3vOUdr6CD6CfXDGtCawfEfOj9u2A
68WDZKdxx0wvIeu8rwkn0NdlLseRDjlZRQ7VPA8Yomy2KELeQkbp4yets8cg6RlI
DrrZxzVyjxp31zlH/TOoGsG03oYCLUTH2UwocUnSAVM11rhVvAN/PabP7aO3n3UR
gyECqNkdAhbpbJylCr7N0EYniDoEXKTnfjE3OTL7bDbAYATdOyFQNvLr/TRXYdJt
ee9YXuV4CHln4FA9zvyFyPCQgOkVhSNV7bDG4j1PV/shugboonJTylzwqrU9rN0x
83tb8p6x3sOGQOg99UYfWFY6tNIe8gSj6USdPsAMwsD5WtQ/cYI6gys0qYSkpcUo
lvZca59SUNo0P2Dl8hK+ZS/6FYUmcdUjrEpT3FGFzzejUtdgrUeMaa4IOMEvDcyh
y72g6Vj3HGR3/gfOdYgZ304Lbi3XVMEexhnbmK65iH/zno3kIBPhd3r8B6uWrRzA
Ld4T+vcJd+a6cPQYoTTTl4KqqWm1gDh8xOFY4VDYCIZEVi+vLnEbv3dswTpXho0T
W9Sv7bndIFupMvV6MtkX/cGhVjfOL8d914onLe+iKES92nTCqEuw72YJBdtKEy9z
wmn46qDSfDguJammIfUlbtAeYUtphrqkTROBYo03PJhjmGdaMMbyhnrSFa3Z8jmx
8umjVtFEh0NSUqm5IM4s5pwwod+j8qIuVfiwQDiaHaBpL+fKVgIzkNncLwAqcmrl
10SWJYRetAFcTLxiiy6/u2+4BOkbg+DBjlagPvTzJ8hVAE5+4aQHTQYX282/70BT
aE80M2ULQ/uVzPLzPY38gB/o1UIZK8aEeqx39KE49oJCfmCfilvtM8J9FwGO5PGy
hZdgHIDGa+FOxvsYZKCrMPeNMxwgtOJ6HIpS9NA9G9cPBEybvmhwdNuD1HaZVBGT
Avp9W+Xf6hTzVDYKxvY9+o+ImVJW6+wDsTJlQymvIwoN1ZbSUAq/dSS1ib1zFSpV
U/T8q1tyCkUEHpVdWdsbdHQBeSIAxvS15gE4BdbMbXHEa3SbIX9gek3009fyYM1V
ZhVkmihJ1WqA3padpCypjg9NmEIjORUZLY/NjkvcG7FckSf2NCYMEPXWpLDhEVhw
emDgJc7/kRt1u13G4AtFE6VrYBRd0MP8PvCkeA8Gml98ZwFO8JpVV77yGN81GhOO
bCakLDynRSC6BFnK5hI126QiM+Fu7L0lLGx5YdwPrr6V+r0h8EaPr9c8JBn8N1UU
rJJW7kSkHGkHMVata9gsbItHQePDacurolCSmrWkcVn3Ay2M46Jwns7k3Z+dgYKl
YIx2ewcBT6ISyimsxAt7heqmSx0TVcEUWSvcKvkVPNpExp2pbZPAqWCN0rPLjcTl
xJwRFmJ5o5FlCRrp0imXZ4aC635zLfmyTLZfX7EZKNL2mSOm01Se33fdMaPFXdFI
WzgL5kyMZtVzo9wq0sjbPQ2sCMA6DZ2Ek4JFIWClvLOUwhOzOhPb/1gjujXMQuLL
Dh+L6AanVDncaesUeYQbRPwBT4L9IX+ppGNcC2Qj/wRGVPojFMBvUHBWRen572L4
y78FSoaDrmqrS3gQ9yceFaMtv4ZaIsUBU9VoUFTckcrspum+1XGe2Vcg7Tv06+nC
wfTt7xbX7vRwOLLjarYbYRbD2iaYyf+LfwmZOJrYmFDMK4Vm/9cNX3FkBcGolJnf
eZjsD6b8/p8v+/U7OH1ekVxIvvdr077IjvRNwQu8Izr1p1J2wfqEvJBEoeHMHo4L
0QRyTuIARmv7wDmA4tVCmtjwrl4hwndbLZLT7Jo5WIpbyiXiRYJ4s+lVCpRDZUun
9bvj9a45zvmGhd5UhrEujdvh8fUi40jDxlKKYLNx0OJlgG2mpzi1f5h4ASrlpC9c
xVDvRlaUbJf2d8CeFikNS8pSlE6Q/gTiZ0acXL0Asc7yC7JUHqxgqHqHUxehl5Vv
n5S5x+2jMvEE5ZI0P6fIY+0Sh8ktQGaXb4scZjXjzEngzR2Nil1Ot/DVS76Hn3/n
q3BHYKqmLLYmivAEdBY3cw513ZlqZueYehpYmoohN9lWeARJ2dVTTcHATmhr1Iav
lyBAvKMJeGW7DCXnLDR+QaRu407F5EPNhOEpJOSXkxmXd6Z4PwPHlpyhGRDka4o3
co7oYhlh/tVIGkGyjnuxKzRXLEAShODbvC4gGqj5w57T5M5XwNS2CSnQFn4A+Ksi
iXS4CW/H2n9X8ekcDvhZrivUioQMZXR1XIvyXHxT/tdMp/wrdFQTED7syaIGVz+V
HkBk82TnYpb+Nr7TTTxirA6JqpQ+lcGQKwPVGYjcomqZED1XU53zP/O/X3m1R2Tw
wil05VCVkFQXykKsxGRV5UOCzyfAPX6XhGLgKsHFIOCp95ZSCx1sERcGzBkw6ZJW
/w2VTQJEEbVzbHaNTZs0IdBZk3FVop/81z+oErJImOXf1uHE19SmeG4zj7ueSkVq
WZHaEb4h6CmUTKAm23xZCbD0pZWO1oi7bFumpwN91SyXXA1ziyVlqVJ+qA6Cqkyq
00EyDwzXuy4WA2YHhzAJLNwT/bsoWLb3WaotJKsDalJ02P3pTYQsyR3zwmxFgPR4
FQY0h2O2ER91NDL68/+CW3DiD63XqstuYRXipGhLXtd/aZdVHWsrtcIJRloObMtt
6gqY1vh6xQtOp+l4vZQFDeNNIYquQJRZIQMhmiXVR7Ags69t9CicX/zwSF6KuT8P
rXfIE4MAhnLQ905DSy9PMZCR/L5wYskoxe3vFLF/id90s3ZXQHH9r+sPRiElOYr+
GUhzX7zzEB/ttxCuoCbEVy1ugLRe/lEZ4WGWRxs9z6F0HVDlpMCM5FBdbhKws0hy
sfsfi6td+iUBz/61W1RqpW1myqumCAxQM5M+a3TwzVnO7yXydFPZBVRpUxGD0Byd
FkqdlyqFZHalEX6crSrh25vTbnUAzArteY+98dvGVGKoRMiAF+VU8eEhmqR1H3Oh
Pu8u8FVeOMvFRHs1wG/Aon7Ykc91O7cieDwYRg3kSjOaV1tI4z/JA4BrhtwedgQ8
59kt5pECuDr2Pdfn/pLzSK74eT4zZC6/YbGdg/mJpzdtHHSIdKlloYSfx81ZFpDu
629VfwjPHUU9FuvXreScqxbp220id344OgpByQxRlRbfx4cdDeY97Ai97sgT9WmW
MbVdmsLsTS4Mdm2Yl/3IsmOdmr/dYbbhAs1LXYNY1jOJHHptt+zAaO0fKFaISg4N
Dyr4J1xoZ4upBacfhN1390DVsZINhatxF2fb1iC8ZeHKnG0/w74VRw294KetyUyj
Xo8SZTjsmAadFwORNNM5QBX+VJbyk8+ahk6ZnW56qAsy51HTrQJVPRDgF8J06EDg
N9wH2n//JqVC2jKrrTGBeTV1emQZ7OngWM8PnoVN2scb8uXotDV+U7vALBfvfNv0
AsaQ8u0v054GB14b/1+B/unaiCTJV+zbIzg/2+9K0H+6Ptu+LXNSbHXNyV8GxuL7
fu5IMoT3SvqbTINI01c12ON/nOD0l4Bs2LTdbZeJ08hlHdihuif+hP3ZhhOgPlrp
7wS05z1c21JR9U/uB5cHM2Pog2vISpAkNWcMYvvATYcEoczclPleexIe+EfejZT1
l+7DUkf7bDHZZcIeeboG/EU6ivSFwIiY9jlhUakAbpKiwSCfJOneXtLkBaXfAdYn
AqZKmoqHgfj6xBdEvo+iQC3xec5gZ4PuRuqExpYGj7Huc8ZLirTE5Clu853v6ac2
D4daTwZ9WFhZQOWU4uzo2yyFQqip+KNWPOmdvwpAHe/7NLcEmA/XO2eQWpn3WXB7
lT/6RA63ueZuio25lAdYIdtfwo4FBFUsNvRo94AcO3IKQOoXmjJtPrTYaofK4ESJ
RBynShn3+Me5zRtQCwkOqfqdN2/5PNKi9LJIM36X04q0BgXK6mmURFXXlPofxztD
vmeyghsmO7MWLRtIQ5YgPvFo843xArH//0fCMbvuxnLmvSCMwRsvPX2yugxiAkkO
wij0QVEMzMqQIXVdOq9LCh0KkfSzg+CM2dkb2+Q8kxYd0wE9O5GyYtA7+ZTbRb+v
ZSkfzzDImqDKGFrND40dC/Ez8mbk9OAXvh/5FnxBCILV737fF93jWdL7TSHNDq1F
5SWNDs+XbvN7mj8zHKA7B8+9BkrMJ7xiIdiBZluDShE6Quqwb10GK+q+h4a+ZUVW
Gwp/93/2PAfAx2vyETFFYLM+GB7PbtjplagsiJJJvi8p1hIbVabtT3QNpctlcX/R
aLVIUfpX73zrFFF4m8CM2UtMkEqmbHF3ZQQGO902Uwq5dCi+ZNEoggRILRqhyJxK
ZLDtshqLVUkbquI6u3wlMoeiII3NagoXDxvEH6BLfsDnWDPrDz1SqoBSWvQukxsB
6Z+Ja5Q2QNxFkzWzW7BiMV1Yoj83hqUs8JStewDGOir6T3lZm1lu7ug/2P2YLhjq
kAZPJCVTZ1P84EUg8oQXRQ6IY8AFIh6gNt+b3yaepMPhFiu7vOpyBechXl6+E+im
1+5fTTp8jJrq43A6VXajC8v4CDNplapt6Qrl3WBlwT8ZS52LI6meKeV17LtOMgiw
4yUcHXqi+t6HH+05wQeIqCyia5JCFDqf8gtuDqLQ+i70NGQYxJBhvdxHKlpf1QHP
8Wxhl9teW7eCa7Y8iyJmlo8wtRTHyPDPtnTp/TOnOfE/kE5Fs6EgxA2/rFGIbQ5K
qLBhZMPAOYMfVFzsCIeJAEEZCpTRZW/HYK+k/y8uF0GTAIDcQq29iVHgb/ENFSgg
JkUUbhbUEAjSKsNx8JXWXeggLfestRqm0mEwIK8EJwGmclPkPkzF2ZTuxTJsEm0f
HtJJ/SblOTF7RzNbDVVt2iTVgmTP/aehGW/ojpR1xo1Ji4HJuh2XnhcHTWnjyZyw
GIfEALLsa3x2+NuI/VmMnFFMXfwyq0WpJ546BKM2gJF+xZPPmcD8UaTsMxtCNn4s
GpdMj7/yQfIH2Fq5CsyoWQv4TbD+Bx7xaLy8fIa+z10A2SiW0hLv1LF9UWnf24v8
mGpa1Bgr2IZ+pZscu6ORxjTsYX4b0sDiKRh09auwVFMQgsBZVeokH1DGDhSwdWRV
HsDjqRPP15O2x3xxyWmCOvLgSWXLgl5it1AGWbwpghDvNusaRrsU4NoxFqJfEJcu
rrfUa7bM46PeLUWwLCr/6oHAkmP/GW9u+RFEHcoCEmtk5E6u6LFxQl2+ao5UWgA5
THUV7grxQRS8R5Pw3CEHiRF0vrYNqEQ38lafNYJXmUIFHFh9kRgbGkn90Y09aKnn
FDMQlcpueSfcp4Q7sUjwdBVA7zIHJU0oJQk7AYMxX66Sh1meMKUMeavuxcHO57bK
0+36OY+b2a87UmlL80/F3OsiqS+5BufikEsmbWz02C6MWOqi6+y69a7uA83MyRzJ
0ZTRGAbSAjwBZ73ngM645kEIWkT0mu0TpKhsgSxW1LChaLTjvtfYcL2fwjYRn1C4
AqtlFZT9faqpxyu8tZ7Luoau7HQKCMEjkSHWlZLYw36xKTBMnu0IGUUJjnS9PDBX
CwquszDw8gBu1HP3tf6+YXKy8nTzlYqe7+iFT3d/npz3eokGWcVwBRuv4nZfkHq8
5V9F0Y7Avn95KW3HyPuwxKRGXZs+ZsvWzz6XzuCpm2P2U4fesaPypOuJTdw6TwFb
NZ/Io3QQESBBmjPyhK2oALAdF34EqA4KkSwC+7S06MsWB4TeTKJAkc8MyaXmDy85
1AWSeIbMNmqxe/zjtZWVwCkBjGCDul2oH7NxU7g5Vh6cxOhbrJUIGVPI3UvIMBXz
gkZAQcxqQbPurAqicp5Le8K4AO5mDo67Ed6vtUR5ehMojwpjRlvsmxpH4uuUm0At
QP+9a+q0LMpnJVcBxddHZzycVL14jCA2OukDeLItUGbMXEgdcGNIDSyb0urbs+ld
VFJI/tzMtrqbuNaIQFn3sTYAXOe2j8gN2KC45ChUfNvRitIFubgiG7+5QJw9EVmT
C0AvDecgGpzp4k8lCYSV5KN1dkZ7ScSCKvl7PnzNdtruIoZkDBsthozTJ6cCuxAv
vAOGL57vS2qkSXqvYzvdqnen6dtgNBX6ymOMCFTEh4JI4cxjTc72dX5Gw5E6YwBS
InpzN2Xm/B6KHFd61TvdN9f1sREIW41AJ9toIECQb2iKsbbIbpOyfT+vXVRZ2BtC
7mB7hkux6K7JKhtJ2qJA5dCpQuKseEf+4xtTZAD9A2Iqi8SZQ6u3a6kpPERdOHTq
yJpxEVQtTrOpfmFRpYMZpXHKCVwYizqLf/rtoHoP7OaJxgYlxbrU1XFOO8XERGcO
WTDP+2C9Q57qEdMjFeP6MeR+7ymZhSSvB55Z5MTibcrfa4HVLdC4cO7YOhWLFXAv
FzIZjnm6xje1u5pocP03mq0bwd795JV4xqC7D4fN9+Uw9Q9o3E72lmOUKJxDdK2m
7ELA/ufzavCPiWxLfqvo67vQr2Tmf/cY2YnshLE/b1rnRsZQnf6Ub6PYRaTbKGhs
QnaGaIxm7Su9kXqgyRZEW8rpwf0qn7a0b1dxuR4qVEoL1WRea8WZ8nG7p7HUoTiK
1xcK2mjdZbDnnq7ll1fQGCyCKnCTRkQGi2kDhQP2UQVVqmvrWYDvbXhdKM4ELljM
p/ruL6w/oyWqPWPDSLyL4W3rGz7m6v8uq69PhiX+NrN1rmmGRn6vFFIRtVpbaKLJ
juFEYJKy01TJ1HqQFBd1zg1q5GtrZqP211gZQHoOMeCyP5W6sxzAGzEAZfVGEeOZ
Mb2LL2f3Az4ysS11gFNYyBKmIYOdq4zzb/WdmhZ8M7Go5ePG2y3TqXuWlxRfLUZf
ys/eqSYC+YRT3eql2uMmMq1BrBWUxA4DyIFpNzhyFSz5wKG7WRGIgP/HjKEmNios
bhraiWy/DOg9Cwe1S98ouTC5DaazyHdlh5SQNh6NmJl8CIRutUrvoiqmd9yJPSYQ
7C5NBR2OOxIoxij/x8GchkBrJhZkJbtsZ3FKkwQ0iRIxUiV5wOWFFr7fQPunh09d
+7Z7Mi+Azr++feuT7dOsIBJ/Tl6yTU6/7qY6+m/V+sErJ4cuz6reflHR/tOT817S
IS4Liobxk9FpnXTBBx52KHehs4W9UbEW8QcNd9zFTJR2bJ7hwmNwdi62gFBgiNCd
D0RNfG/Am8OA8tM8ZIakepcUMCPqScVCIndb6XMa6WA+9TkQfm8Cq+KzRhdNOLq+
gtF2ZQXXZWnBZ3d2AGZJypH0AOqdMMs0qDxkhYYEBXvDiEyZhAQPzO3BrLtsVvk/
/rIdbZHitUiA4+Oj4pwSMJ8CxzUiYa1qGt08QMM7AdZTSVYGHkLm27tgWxhkYuBv
wrs45kI8aIe2ScYrUa5WBcBxvXHj/mFQL1cCAeWPw2IZh/nWHUo6lbUe4r2IdB12
1wr8JYCSQrKWx4TOIWteiVHrvOYsZygxxX8G+mBZIglB8zsJMMFUgVcaBiElQOUK
S4HBVtdKNWym13l58Ym+i6mtJxOzncV6JiNe8XcV6NVP7FypC8V+6croVQ0mIjuJ
d7VtH3SWhzWloBmGm4aEaOIQg4Z2NTZzcGDamwGykL1uk8Gd8LvI2TyZtpfzHn8v
0QMIgFEBksA+io+3OPUkLxe43y0GtACc/MNNW0mZu5ZkZbo2PXYLvIvsdRGFYXC+
sjq7Lj0Bp2ECjO1Ylts3OmXngrABX20JjzynZrwLMCm0YoIU4k85Ic6zTsbLckxx
LIwUNuqNUcAIZIiw+HJk/DoQwfcQ2tQ81mPSeH/yJM6+t6WPKKOCnO8l6weFvKQU
gd661kLBQpnHwh+jzoy6XMQQHHQvGZP1C9wCEAc36modyRhg9fhyeL2yydBO7dxk
Jy07Peh7CTbSEtXAs72eIcNcjz0BfVcFEyE16XGW7EemDiwzQfEXGfBzrdy8ayV6
AzU+wljwyl4tYy1u6ZlPtQ9bWumgfuZSSGOoQAA7JIu64IxJ2lAuPvZZDD++1yMG
MZTFxcKL/eztzibPWzEVZtVT2LHLCUqh6IAdmSODynz8Ymaje81bAVP50IJamwnT
HkT7DS9AoMHUlTOt+e7tFU82ZibT11MNZvG40zHk8cqI+kDHVPNE5780cMNjucoJ
w2Trf1MtNsonHtX96+NSQ8JQgmA9g/jxOYrningKxjCmyA9LB7/h0VlWxGn46FI/
8+dbx9LZFH7NKcsdpdR1fik1FQmE8+FmSz/36/jFDMMHVDSa810WBfG2/nxj6/9J
/MdrRZEyFLV594oOQwsdIRyXsDWuLTyH/Tm/SXT97eopMR4lLpJZ+mT6/yatNM9R
aN1IzRIR6mgzduFTBfpnGcQNEEhzEAIZ1PturT8v+FXCJ+6JUQXUWpGwUQzZ/iL9
Qqfa3zmRnXOgtrCktDG1EAm2jd1gEplIr6NQw8xlSzYhcCx3HnztY9JUJvcLOIlM
IzY4Bf9uIuhYa8cCcEaIuyeGDPN0SSzBwRkjhYHK/J617db62GEG4mTjNvIiC1sM
aUVK/ixNRJbL0xBh1B1CQrmNZV8y/ZkMsOl5GSFUl4JblV+O0RNmDOUlG3ohjoxu
FcwZL81YBrsEKjOzRleJeThtTMTZlAH0yap9RwTYxLOzc4quUGuAlFLim20jvni4
Yt5yJ2rryO9SKzyQumEGrs7b+5opUpXnaisjYI0o3wSx0zykaeRgJ1xPmrBHR5bi
HeKQbjaciexa0vwL3j75iTjU/PVB+xeeJNs0sbmWyL7lcqdmOoeGbHPz7sWwsMXL
cwVPrmok+fVU57YqzTh6jG/XHDU2EzitEU+qT3/i1mzMI1QuqsDz0kzbN73CX6tk
u08hcj9VrkpYxEmoSrBTSr9Zke3/O28iVoJIXucjg1fCPgiz3CTwQuw2/o3oMNhw
iWPooKpUTetr9m8VAIxDXrWHp73cOkTwtLGH8AnK/YjLPK13wXbLrNS/YASuZ003
PBM2unmjOHsvD7VCPZW6yhg1DvGVknpri8Ek6LgDb58bhQvm0NUqCCjL2zYl7J8e
9ahtnQPmsvoHG/IQinsTUDHB7kfqvFNPohdduOCh3jIr000Wp6FIqfafKkmtKIOn
rIEfvLHPYNbZvNfum13yCaeR1rJiTkRzDHdr376W2cqIMTh/orj01RbPLqfi2mEv
ZgUoUF7K0QZl31GV3q44ln6j2r1WSSHL8ZGnFU9rLQ3RZvdRfJTipXYZD7p7851t
HJtshV8GY9PU2Bysg3ZnbWOlP0Je8T820cgdhOf24d2n7mwq93TwHvYSQElHBahT
a4uvr4bDcMvqPW9xuRJBR//bIE/wP6tcGIzJj+eYbNl5OvibziJmReN09kqQNM9a
kJ02hiy0Si/2nn6fiMPsRz9lRo5jncVyFsIJYpzQJohb5EUs+IC8FI0zoRaeHBj6
6v1e+Lm7ocOnBrnn1eRHWDteNX2M6P7r8qvjm1IQNEpl2PgjrJbCX2MU3fx4Nk7T
QyFyAsNlccTJsPauEa9ZFB0Pyym48JcAocX5AQyx1xQPYHmDOVT2PXrqQvYg29Rf
eDWBTIMf6bMJiv0XfMy/N8uoXajRg94qyOFmetJ/a9uxIlN5vo6P5zmoMxDWjcGJ
30a3EXZCk5/rHXGYFMSgb2aHtRxlWOuGtKuH24jHlVcEmxZBjoP/K3rEV0Cp9Mo1
9E9iO9kVbCT7D1bBp8OEbojBZ97wQUdbwQ+vt/mFi3b1xU1c+GeOIaANvJcN7JYD
53Ty35GDSf2P1531GqkruziU1T5G8CmFq4fzaQNGEZaULvhcYJcIsqViTr/iACbZ
ge4QvzPyqUx+meYd8LCV6wb8vAkeow9IxclpL5AxUtkNUPntagyBr/YAP0kQwAKX
IAZfqcDAQaPvdxn/+S+YGQUDYvmUHz0Pl8NH0L9SygRR/7TuMzfupdltRh2T0WzQ
Hr+2fiezVR+HUy8mf8mcPjp9/estZYIzmrBqUYfG7VqCu9KzWzKzn6cZbIpgg2qx
F4/06DccSLESPXUlPdlqzr5yza1HxGR9vyVpoyN27l4lgFkTGPBOe1jTwFP+hPpd
7/mUP7NMqN2da/FWBAOh7r6yYMmpEVvMUsDmu1wa75uJ3NPLULwaTTt2hYnOjNGr
vcdu0uqLZR2U4uYyQI1FSIba9scnfr30h1DU9oBYMY2xBUBmqbdbU/ZUrw8u1ohq
xwpo9iTBvm4x2jw/R/j5VvH3zKBcC03dToF+kqG/wtTSrk3pDagERAakpBVmrTD3
7wHcLLpKwZFGY/100dAUxhrt+UlVXUt+Dffv7qzu13Ig+WJG4kcdcWQSA9RJM89K
cJeOIscAQYacF6m4ntxsRYH8AXekqV5gVHUTXOVlu42ZudzJNJ7Ojk0RcyRomKMD
1+/56rYreX4trEOhTPXfMz3E9nqEWOh3UL6XSLVCO1RQbuMSo1GexGxMjCBf+8iT
nvWSraBeFKZjLVRa3o8R0PxFLnhH1JeTsM42If8QMXhfHyqWNg3fF4R7RVef2UVM
Trd8v7e/kgoMGV5woR6lFRbmS5cJHjz4xO/PTp3YTl5o30iZIagT7dB8DvzerLZQ
RGCCvZfRJC/4vjAgsqw+H0osa14VHg3PgjCtWjuGyc0b3slrEQNwGVBdJnoNPBhl
GAaXzQ516yw5ItRq1UuJwTRvJMUPBJtTD7SXTfNTj0m448R0sZbWOom5/CiXl27x
QNZNAWrrBbNbTJ67bNrZejwr2qImHXQVLR5epa3DyVnQBSueTawNXct+aVxgFBzJ
QQasG3a+gaZ7ip9IHAyqHA==
`pragma protect end_protected
