// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:34:55 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
BCi9Sg6TpI0RmBkwCFpUJ3RPTcEfK/2pXKuKPLEYL570m3nPVgOMeKNBt0zOFHQ2
HNp8eHcdAbtH9S7iXjiMPvv9NpCpGqweO+2XClP8Xs6ThMMGKDQM+XTR+px67ZvF
OKa0wdfHhQPd6cvSLIG6DPO9Q+tZYD4KygpD+8NMFxs=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 62448)
PZXd5t0BUf414AQ90g6hXLA0iLkvjMHK+/7nwVlXeCnv1ZVzkDB2wM0u8mxf7U9I
CUlpb3D5gfE3fnG+/a6p1axhqrvbUKO6q13dIqu2uN1WUswFCNDShwJkN0KVIIf5
S5m5Y3UhZXspWylX4tMIaBHgLkyzvnBLnHtr8eFgQm1CaxwR99ST94y1nCBSeSSC
hIsGtnOlrqs8Zu6kayZL3huu0OjnmQle43Bs86yISdspZGrk7StdltkiSweY7eZq
R8ZFXOSm2sSaC7iq3aj4vjQNpVIV4kWF1O8E4U3U3oE30Bch/DEBsjLqbFqAipCc
w6HjfTTO3PflICo4AqEU42oRk7q7u6fYcP5R/G32tCrMf5r24QsMv2O9+UccCX08
qp5K6O5K7GN/ZZA59icYMGVhyfoeZ9J15ZQLV0QwuFgjf5gIOnf1caQ79i6B2Bv4
z7A/qrajC27g3DsEp2qrSyybiIuPz7jlqF+a4CB75FbMno86YCLu7cn/8lAW3B4x
6Tk06zdSxHkKFogKCJZ6WEtajpoloHPxn6Z0KEo1ZHY9qqVPd8452Txk565GfG37
C9PETZ7ntyIpePSM1kb1vV2YjklVs8IbqUqJTQRN7VKycWCtqZiRxIxNOUeUNXAs
VDBnZ5nZanvH+I9fQcQycw5RqBK+zquQHRBbjceJS4O0JEx55hhCvyzv1VhA2v8S
KehjnbdGzEgqOP68UPJxz6JvNg2y7pqlOVnpG1sP38afC/BK/VgP0v9GTvKbzjHD
MBaZCxz1pKe0ufpmVy9MzKq9DhB+Cr4jrjP9vVtSaF5zCwtSPDek1fbLdFqQvCC2
G2kbQlrcYzQVKuCMm2IeqN6Hj9XxWmm4zcx8YKk6qkuQ+No3YbAb7wuSOcDHOfhr
wN3J/6yjbgEfHEveamqrKcME8xyIaXGRobYpydEWQoV0GpdoraBoBNAm4NNNH/HS
UFyLITQtyeI9oiKAxnEwgzjeo1o7jG/ngPClBiRvD9n49ML8fSTc8qzioTEcCB/t
MUrFtb5rO7cdeRh0D+X5suXsG7RBsAJn/ErxgXGY+Hl8DXCGND4fVzncMzOMOBxZ
4ItQ7lAhGGUx9qAouPrvX+EU64Q5Cduinxdl6YO2k/P9OrQfEX59nPw6IVPJ3mp+
PtEZ33s+YhQkf0BTZTIY43qDXVQ4XzxrDS3enzx0ueXzhmXH5lL2b95jjiC8dcSj
938c+rhWgzSykQQbEgXdn4p2+LJZECt/VNo8HESK+LPGjP0w99fDOXalhTKD3yd/
+mLNUiZ2Q7szVrnvkG440R48dPAbuBQ1KKW/4bP8awr0KNg07hlhZM8gSm/uUdgX
fr351ygrRJTbl86Q2h2oDaY9+b0luY3nDZpgM6mJ3WtL1l/hsRyeeERHLPiImIfH
xOliqNggLUR/Ji5Fkh6J6MVEjp0N2SyTKuxg3f4Du4/izVPUKDIXWakWAzfMv9iR
Rsf+Nf4XMxMCgzkO6yu27TH3McROKz7q1vIlXhBngKHKxTqklptX0SaB21v89jWc
KfYXhpqA+ppTUUew1oNiKc3lfJtuJJrYsuRJqNbRbJTNYeHR8+SmprNNRlZ5TZhH
dFCKs+Slp4IgdSxNzGvEIo5iP/SkQMQKHeM1OVg2pquy5+LVif2uYpnvr3evjnKB
BtPNpWwcHMAUSugbcCUCv7PT0N+nulFNg3gVOJn0pFUlsjxujZ5TvOwjWFxlSI/i
H7ClDRoxEanO/ZndlCYWivCB/2/BgzBzFGwZTugPn1P8Brir7DJj6pzYCo1zMYTd
IiQn+9LskxFxOHAL3Jcu6/hT7zKLP3AGP8D1KrHPuFojrn/P7yEaHnxI7niA5hc2
CoTLDIDtYt2Yl18sjsfAaBz/N93S2rjrB5MsoCDWmcGqZbOvQ8vGuzZ+51jdiNHs
z8tjfK29nOAUDJGHbEfumgmmpIbzA0l7gH27VkK4O03ZwKLGKqXrvrHxsW/z0KVq
Jfgxu0oFmYgxaL1e3BsfUn3KhruH4qKCG9TUj4fTBRyWEffpnRUql9lt0Ifo/Ll4
CCvl7t01qosM4WFpfNoo6KIjrsAjSloW/d8s3/MLZVVh4JgTz1cHWOztrHNFGaTZ
CXTe89JgRLbSNBLtLzlkdyIaghpHmtYFf2Dq94mJJjAI5T3sPW7Ndk3wcTY9xoQZ
iapYEoUvocWXAPEQuBdUBlDDd4boRYngo1EYZ6oWXPjuium21KWJ3EeFsj8NJxcD
S9qDuMu+UXIyKvGYaKVFBahxYmTMNXynpSDW74FxAGe00qPCT6G89we4Jz2ySCO8
XYjZ8E+DoC66anHxvbVpTO5ppP2zJHPhSM3wdewNoOAoz2veshA17yTHPTLQpbCY
/CgFl022oGM0HghtO3lMoYxO2cwGeLvMu+yjuVP5FNq8LVJhVGO9OOnd5pBCpDR5
vygwxladoqIMGF0bUtpCJ9P6gPYfMrZlU64FN+AGznVb3w4W4o7waTz+YKgXanu/
Tvs172h0y2SgkrvsNOqKSdgqRHXs8oJzKAVrMXyaIQbK1NVYXjarVdG706YDGQdz
BgyEhgDrhLcbnD5AGmcZeyhrtF9hYkAbiwPgT2KRzfNhVjsYGbVMi08na/b50Bgh
2ujfxlb1ggjQnfYeQPaSGzBY2pY4qaG1X4pzfY6wVsypN2fMnp7M0IK8TKQZxAo8
d0sJmVCAxm6yLUNRgQ7eeFRokSxYNW7vr+cfa2OxFE+NoWpxTTh+vjLX2OSVASwR
Io/y/FTc6O6WtQa0ihw4p8rSgsJamOPUrRoZnyy7h0sw+7v+HIafhaTbvnLF55/a
cTZSOWhGKKnpPEeXptXGMbvoruZMs4WabxH8i75RxPDLvJaZ4qyYvEikWWzOE0Wj
RkNzAmIVt1T6TEneQ/kUTvbPAaXsk9GMnSm4ZEzhTl4ktNPdw1Fvd4wcHQ8XzTDd
vKXdtT9Pke0fjo8prwC16NWUxEqqJ6Ba4FZs6zSbB77UDLJnzP7JRxWoE6yKTFmH
baB6V9u90fu3d/+hMeYeppM76xmPZ+rqEhjOBpXomWNUUZMPMADmWUJfQ+w/Qkfr
lIFHL1+/8Ao5XnneU6d4J55FswrxCOQydaFvCeTsu+WTMuI7nwa9kOwOcrasMd1S
06NhoqPrG0ylhVSn1b+tL/FLiPD0uRFu+l4ZqoNeNHOOiaRx0ErYccELiVZ2wnqP
9fyo+Dm6u/QpgCpXyXAjU+TD2W21/7+BEHteRYKlBawTix3m9dpP/Lh5Y98Tl2BT
NSgIHrHeHvZkEwlqAiJk4jQ8tyvyhdMX8bmk/sRiahfeyeKGnJywszZioIh8olKC
6bRwH7qkzVEzLeHRv3+mSqovsJ+Ub7oEsfsBw1bRKkQsWipZ1jst73bcCLV+xEt7
LMXWj8hkY/hi3RUIE2glSmls/uJ+eEHmaW+lNs8CFwW7Z8EtG6M8f+sKV2AU6lrE
zAN0obWFznHpGP4OiOBqA5fFmP1mtVIYeB9h3gnhgMrIvGJZQV8HQeI43CYxPsVd
Up51/dWJGHENnySJzY6UdpaV9bJp1aXqM29q1g1fr7tkKF4E1amtKqgnmy2QKCK0
5qQlliAYcWVwOzVLB3EJKBzryALsF4rHuFS8G06nn29n9JlCePm/u9VNBxOHx9Tu
oyv1O2/xWuGZywiWlpsq2QGFGrY/OWoF63dj3HwQ8AwDc5wCbm0vwdB0XkXZDL7l
417sgkMey/uOBFikaYuORwMmhAxuvoLTWJH0mB+I2kcTPN2fzxvL3RXdIn5aIH6K
PLJWVyHEVthhckj8rc55BYrRGCV7NZT10Ti04ehFmqDrxvo42C4zwiIZdXG/GXw7
OQu/cBhocoOuNdx8RZRfl1Zl8lMvyix6HWYhDVR+PY3zg8siqjIQeDvmhTVORTPc
/0BFImhbE6D/OZ1qRMwrNIt/x05876f6vWTdmDaJOAbiuNoZOmP7VS8laO+cX1J3
W3KGEUYBaSfce++u5bO+YCNy6tuh6XBfTKmeF/hSgbcmvgdQPKsL9mS2hiZZV6ZJ
gTrBB8+/N7Mtff6FBorFvdx6eywjrctNi6GC6uICVqWsLVXfNrASJOqbg+7ebLHj
FDN3qCTqbGCtEI1AtZMTFjYG6MzqEowpiQ3BfeqaFS76DxTJH/6HOL3UeAx4pb6j
gqFbEoJVRO2kQS9LA+2f9HzRGCuv9HSVneq4+x3FPxiqscHclpmUVWCuCCRhnscj
JL+jKKPC1cUb1/4nHRQ25Yc/wzRwnX+fqFINvHC0DMB5qByVYWPHgCdC/9ZHQns6
eyfIjqEsA963I35wuufGrd9fHKx84Thw+t2IyAUfnsBxpmksF9UkzOS+NzwgM+c0
luOgipn9JfHApjY8TmYhShqpxh27MYGqSK2npqniS5AOgM7D6gSPw/8rtH2nyIQS
orISpDPvCiBJPnIeeUTcS1fDtWEKPXj+j8DM8Vc43HihgHPJrkjALyznlYnYVDtd
jyzLTz9wPwjKlqmITqM6B47wNVfwl8tY7xWupSgzaKgvE4Z+BjZzDAbHt3p/UxYG
qvn2wSU6xriDn3CJ76zFTLe1ihpvwEVpISxLOGA5NxmVGKJ69AfokcMZFdpixOLK
bcZ50AGpVADbfZgQdLVv2R5uoNiq1ecMxHM5oUnNWjIx8FdeOOozAh45c5i3cH2E
VRrimgyDvmP/AYaTM5u4Su2/pWfqOrZCpAGsJOEA1Kjx5RNHaSun1li+rcUu3p1c
xLD4AR70jncfps0vS9jo/83A8Ofu+IkHR3IbWcqGMDvcY0S83jeVvv5ObEGWxEwP
MMoXTjdgOVAPEOWiPDxqylIWimSiEMFMklUmlhghLLFRNGSc6oe30Oq0/RtpQLx9
dnIVZgUyqhiHSykciExJ40SOMDvKtK/zIrbB+IonK/Hh5J8wtlp0WzKiTZxMNxIa
HLZcTQ4f1/Is2ft+tX97ngPTLPOfpc5zfzZm9XycVhCCO0HlVC9odCx8xwp49QLZ
W2O4xFktyJ0u24qVYtu0RKfsm4OCpF/uG8S4XQRxsPGQz64MILw9ScOqjm6m0NY/
Ddd1xMO6ta8cHINMcikjtcKlq+HYMCkBTq7jeCqcmftOHNn9aWIOvbWcxrfqemb1
Be0O65d1zY9MnTqKIo7YxP4tbW7xGJyXbEhDNUgJe7OAx7tLIZz7cUSebE0E+Fl3
RBxfLHkAv1/7SrPUQJXAWs0sMIkTHqxcGpMWZHJORNac8nYm8D6v7i7/72AhqrSm
91bfAE6PBH9u7QY37ddxoZwx0m/0Z9zHM+uZgEE9+MqIOYu+Lybkkl0Zv2fJm1yc
IvPWBQcy3HotvEZ3vZu9d3pKZaPblUn1kdw454mR/R7INGVLSgaoHkEELYpAl124
ge2EObOKI+wH14lqf/7+2qE2/bQOK0wLIJnI6mJaIKuHyFkkNimCkcs1NkYa9TWu
HSKgCThUKCx1sj2mI4esAmh4qXiFW5bm36WriYRQsIfeBeB6zijExDoZnQy+MROH
OuPM470h9teomRHUADGnIoHmM8eEvpJCbxN2jn796R0AEqltgcqu79rxRbTe8aqd
1UFgFl+JS2LuPxJ2fgkWLALZsE2EbiD0ujQO61kryG6nvjNNt/9ifCyJ0mgdSlLk
GnS8etHStLeu1lSXbN5p8+jaBgC0QtSseaXRjCH8P8EKCW4NiqqDCOXMw8AgHTe5
h9UFSZiwsR3gbRnhqKYBeia0ez21xnoH3TjJ19660CwJHSr5eMeBxN8TJnZYgkkh
2CTktqnJCayMfY/Dv7rJFB1aFgMxMJ1dKCqxQG5U3l14E41Q4nRo/7wzdquqk0gV
X7SUJhbRgtQ2Spd6tx7hx2H9JamlseAxHwoI+t7NUyRzRRJVXwVDX5VmJIcg495j
NhVVTD4j5xjF7Kb35D21G/4oXL+zLjs72nI7/yN0NcQNPN4fPZMs5eHEKzatVeB3
tmbfMdUChJc2dRQV6Gam2FGB3VjeNYC2q0XNj1+ih5eDHQgKRMpZIpkFd2DZ66vi
8wS/Qs0r7N3fuyVZgNf54CMSn60NYGKuXm+NLHsJ5+Z+U4GHbo63RNjbM4Am8FVF
pIUBIG/g1BH5JGd5ItKAreNrhJh6ZEE0+TbUoGmCdOzI4ox/LssGA6BG2f0f1yBk
eyYFgq7GOyb5NRC8o42dxyL1zv3Sb/ssHEgF+MOIjFjR4GYCH74TVYjAymLJf8yx
z1obomTcajiUa8cp894xw01ccZBaxZgXmqoQ1DFQwyYV6yiGHvUc38Uvrb4fW1qp
a2Q5ZEO89x59OAWE2AiVxLx0KYEBehfypE5uM/45uA4XfWq1KffHC3dF1/ye7WZg
8ra3jtXI0i24bN/lb2bMlaBGi7Vxs/JcA7I6UpZjHhVe2QvaOHy6+MXmcG72t0a6
+NqScp64XlwPMPPYEQEoizcd39rfeZ4z75IkII8G8p0OclRiyBzN2Jvnb61uoh7R
pcqyVEO6xwXy/i4umvG0nglvp1SHN+kCpHu4TSTvmNsEWymQMOijiXdDF7hnbd6F
QIBLozOsTOar7SZpq/JpqN38l5bloh4zS5hi3vplUhpsUtwLKTMbWOBSgWGMe5zD
4ePDsJcPXtlsTBTPj7olwNiw81Vd3uvZUfAwuw9UWPDC3FgyQXNzrxl5qqwUIZnZ
uG5OSUkzF5gCWBwDlxEa5YpaH/EHjn1/qOeksSUVus2Gjh3jW2fESUV1MbNcsqD0
3Cv0sxQIUeNG1qzt6UP1B40TBvbgrQs0IQGoUQuiXbJwfMOscO47xUCd3GlMkras
Z6PW8ZDfP8ixhGOzUb/tf8X8A6HvjIi+qHtanTEDw1pzwXaGbq29S/rTR4LT253x
DoGAFWa6qQ5ZioxbjZ+eU3D9Hrd9+BGw2ZbnTPBFb548TOFsxx1r9H2PbixEr9+f
NayLq4S7AUIFEVYypMm+k9zzUCOy1jKImnIbn1qeibtza91dOJb3cHxJwMg+91pU
CITeHiAFHAIax1QvI7S1LJcmzFjXt1kGB7kwFcgNMNG6bfp+AJ8JFYrxts94uaTq
blM6QRzRVa2ZilyGlpvP1aIthyG4MUxgDUurBiaOJ1ZL6UaVITX0/6ut7hIis5cj
5UDBU8HazvhGJlvx0vmAlvEcyPx/paItBEZKzROF3+Av8RIOSs4ze6zQAMa/V4p/
I9fE5GSXlQa2JZUEhvRddlHyxeIohbDz4d6J5phr4mLK18tjXOFvoCnkKxIMmkAC
4F6yjDw11gxyKhPOc+J0jdn5ImdrctRhyeWms+j73MGOYpJT/gXY6uUGAHSD4Azm
ydX7+QaAQVN570FCEDzOnrKo7Vqdf2MefLinhdgr/vwt5nmgpAxkZdM222AjzufZ
Nc6eFDjTGYORyfCbQaq5JWKdMi/ade2ewBC54/VvvTnLt/LSn2/66M4DbmGzL4LD
CcIZa/n1yix3y5qySR8WwVHPr9zRFSXUi4faA5LpNYV+o/+NUA/HS6rjpnHeu5pe
A/t3zO98UBTTBsQglIqrIs+8V9ew4i1RhWRbT7W0+H16lXvwErzwRlZ1FckVlkq3
S1hS59ygTLsLHG+RO486S26Vnwky3JRW/Fnmc00jb87JLUqROWoq7qLbVdDWjVh4
/dADJY+FAElSZZFc83Rp7cvJ85FaN3D6HWegW/ePJd9lzSHQVUkQXK5pMJKdCvcN
/TPfx3Ml7a5SsmBY4xbeQJMBb40QCWoeqvIYYSucVDSXCANDf8zvwOJiaAoJeyMf
4rWR17KrEYBKJhwfd3zPLYgqP7L0UmZHb2sMhQYNdQ3iok/h4xUrWnVUwtDx2h7X
MUxAcHsJIHxSQtoqVrOZ61TPjhuT3RNH9E5seDdaC/11P4u2uB+LgEkdQl0tZi9/
bUVdxYIa8QVperNQo2wZX8Qs4kfbCCxIT6WEm+V9qJJ1z1MloH7jlj3QOLYSz5se
fjV3pM+VRRTfu+WcRYWijU0PD3DAyNIAXTslFMdkNMSxHoTTGo/ixuv1rGTR4ynm
9BmO0Z5FyyHY4FskHIWIsPyDPGMgVZFgV0CdkDzFKyumwxXXn2HK308LpdaIgiYw
rL+81OgRcSF1KpNxfNSpUpm4+xaBgJOgedw7swNxF/pcN3BFyF9lzVvgD/MLS1VB
nYK2M5v5eTU3TeWihg3IEvkrnloa0C+96NwdkvLDPe3JS/lKPUSeoRRSfjeby8sO
vofq86XruiLGxPEAS8jHq7SqFzGaxuLVtTvsHJbJXBi7FUvBe5Nqk5qcBBSZkIXa
gdUkmPqlQPtK62XF/xHOG+LJtGO5BzSEhA6uVqjNxKZY1kWxNHDpKD8Sjq50lJsh
7J0/LAilouRrfpZFQUWvcowYlVvVC6x07Mno9HjCiMyjinc9LWwIWvPBCI388abI
kxYOE5yxaiPRefmNibJWUw+ZQ2pq81Bq1xErAS4IfbBJahU2CeyiTIe7oRG2PQX8
sUyBE8n1H5K1VOfl5e51MwRhgqmsIwy0qMgrfcOtzeRP5DrvWcECB75mvK5hfXLS
13Ohh8KyCyMvDN7Bw1tuBQQSv1xiA8ODIC/yGjT4dnq5oPrBPfCaMJXBaNHDrQ8e
4kNGdhwbD2/xrbn1tZsQwWiBChwRn7p/dkOfn14nIdapXJm2CxC/6TW7LxBJ4r1K
m5JQOBsshF6k6ffgTMH1vSb243avcCpfYxUHNHPFs9Uzcyrxn45Kzh2zg/IY1Yh7
pT0SwovP8rvZo0cGrpmFzcTjjdZKVmTA3LorGrpKCCG5dN5O0wjMEd+r4m78/2N0
9LHp4gEGdO79AAc4Tt38qr/ixuAcIt10+5+pvBkHv/lllFxYYAEy2lzldVvwhsXN
gKU8BD87e7YfVjJNcSQF5OT2fxxY2b01lxDRXpn3J3i2zqIeAMd1LiVNEyot3GyZ
ctsIAUmczTyxRB7+VlADiA4wgqc3m+N6il6XWdtyu2zl2QDJ8SS52d3bEJaxRXC1
ftbMGfqgNw+FAnAgoE7XtWE5hzQGJbgR77VRF8kkUpHWPXKEH9nQ4W9vdSfhqKV1
P7tSAWcJjFpuMyAWz2gHbBjNA0G/ZDnfd6IvbINWoz3WHuAm72MDw53E492LiiZh
qaOQhXCg2ToWDS25vNWUzqay+N9HlDsktqLjGKXAUXjcVu49mi+0DTIRQSZvqIHx
cJF6B+nsmVK7DReFSdD/ZKNA8CdOf79kzwoYBuRy80/SmPF0NjjXYj+WL24nbyAA
8n2hBUKYxB5m5z6AUUEl7VO6Eu/Xs6EkOjhn1x9XnLjBlyuDG7f7aJibMdoEu4VA
WVERcbIym7CIetBEDaSj6pFqyLTed/Z6Xbq40ZZVjVgAVNb05btG9T7PwuCdrOpu
e5pH1HjZRclqERvYrElf5O9iQc1A+5w7SSqkabzco2iSPryG6UquSBfFAxm8BY4j
6kFpzkvBZRL/8w4mMoytZyEQJ3hv1oFitzC/PvdD72RGxBp8C2aWVVBpq/xxiGcf
B+/LDcNcJLWMvUinZuVD+Ss7BClLUYc9Vqot25f/TwNUAbxT2cnZpjWYdFMKmFos
RsQNllDU88MfGoQk7YKpEqVn+DKOwNDWCcyP7ytdgHctgSo+f8zB5EoE4l3uaJv5
Zqi2HF5UiQpBHf3zxN3XFcR/WpgvxfBytLp9ecMTddEf+GVcQMBDzE7U855BZ5zV
wX+5ynJ2NgoKOWchIgM3gF+T+vD00c29X3cyTNhHiBdjzWJVqb6Ekr3j6GRdesyU
G+Kv1nFm9uO9uS0Wlxy4Xl6IrUuo7dW809BTCwnDlvGT8PQjZkEMl6dKA4zNu7Q1
Ll4pcR6GLPq7+0AVbRr8eesLcHROKgAt1lykAFzWfHeVsIkZgaGY4GZwUe+EFRDd
ITKX4hi2TB4wzhR3c9iUcR0Mz6uvFFWJXnNwz/lenBoGmDgClWS38TWPjiij6BAt
1YETj9cFPJokrDIBszSZthgAnz6xnAVpKqp+IEVxsHICA1mU0UpM5IPPnjQf/IBm
YtEJmkfVbQhhYluPQIvK0s6+cttF8dQ5D7t2FrRuahBFzkrAB8CE+ia/K6xiyrNC
9vtap+i+8WijwpA/XLo2pQzxWl0O3J1ghr3p2TRSeZNxqpUb4Tv3NWwYeSF/Cu3A
kKHZD0GZzuQ2OcoJbF1ezFgLOKaw4dKi8eGpugvYfgxw/E4+p+dAqUDQhS02tX3e
d9ihWrRv+/kt3fm9IIqoA4tyTXH1eFeGdxR5j5cNpzOUMAFSTVwO9TBdATBP7itf
zN9RbjPCVEmBM3VhiHsylIyPSl38mkJz+u7lsC33aGwuBPYNxpX+W9Qq0ZdRvvf3
IDHbEcDElI02s1Lcp9P11ajpHpoBm4XzBBTHeZyJ2nRgHZUGxwOPG2LGpnREdFCZ
e7eut9yzVgNrr5jU33IhF4NgvzflhEuY2RcbgybAxeFKBY0S6wRch5veAk/a6B8T
gFxIqH73NHuBAJYaUBDHD/OItzk8jviSIsg4PuNT+y5ZxH+MRQBiMmO+7kLZ4t2R
w9T45L+b1z90UKuiQNRWdEZQ9ozw6j0vX0jg4UB6cIwloih4L4BPzhu+/osHeySG
owzs3kxVe530cjpXt+bhF4QR+JDGVOZVJ2AvdWI8FQc81YZrVSXBffUwK2xvcpWA
DVhaYSRvK2d39Eo2SRnDU/F4B1cBwv0KDA66ON8v4FgJy204ddStGwY/HE6QxT2h
Gy7/RXua6OPi6p7jfU6aOvyPAA+5gugywmzFEO1LKJIOux7AfobeTV3fuoDY3ypl
2c3ajMVEiznx1Df8oH4TXR+sBiUC0TtMHs2ymwH6thVPvx1NbGFlUBnEba6nAV0L
2xcOG9Q0Ng07A/w2vJnVzxW3E6rHoraJhQt3QpYoSnR3CDiCaHuSvSha1jwRPQml
OG1lV+lODSdy9e341cyBPeQurl75WXVnMgKG31k+y1rgeDQYguxuNTIsRbxJL2G2
rA4UVLAm2NWMfuHjHGlIb7krM6c6m1yASk7HVzUcXXDUQNdujw5F02+tiyLBj/sq
jL+SkTOegv1Oi1gqR3qIskPgpF3cv31327R5U+8Rz90Na2QdcmSjlFBFQSJV6FBC
/YYLkmsjnc0ObupMAho6VCBugDCdiD5KN0f3X/oGoL1+iI3JjImLGitJfEewNJSd
Eh0S6NvJHWhoeBogpPI3AJ9Y5/mDeVRJYikmPS+CiCtUm+TuV9qMG6aKl6KDSSO/
8+2YB0eBdd3TOb7IaopckCGPq8TwPXP/RkDs9lp7XBQCMceSVwhUq0pw7lpjaPoZ
QqpBkHMJSTOP8lz0Hzu+Oa6Zm2agc37dMqYzHnqhbqlJgh6k5gsA/boFCCLDAB0f
vAd0okEsdYGjxcC/2AoK/qhZ4SN9v3gQtiKBCUGWjKqOtOW8l/EtvqIOcIBVgeEL
+dNCy8KMuFjUDiQ7T3fd/li19eMa+oZ3Cp/9weF+ND3dsZCD374pH03lj+fJelUD
8XKM+yz6g+ENaQaImkt/2X1RVdoHLSeh/CdnKFSbmHl62rvW+/JB34P3CfvFy7Ir
yD8EhMxkLQF5+FlC4f/Ka7bkGMoUEVOtXGYRcoe+gRneST9Nq2uyMzf5YEuNW74O
q7O8Hm395fct1T6wmrUjXkhp3VI7iHZnVI7qXBm5HFR0+Cu9FAG7PMjJz4iGHGX/
M913Gzpb+nsCOQ0jUo91oe4FYmfCuqbTHKJU/0oQoNLOgoEKYYGvCJ1ZeVudnz24
VsPEikAr0wXR3D6thPmX41oES5TvbKO6TCDjBR+xI6z9fxdOSBVU7y4Rq5HU4Tia
9mWJZyt0TYee4ErqgjRVw4k0rL0G3yDqu8DgsXtyTqouduOsUi3EY9+9TebFhabY
NnpnLRgLuVqzvL5wTKQ3yyU6XjuwLORmN4BD8djpkgFrnvthNlRPMO9V+1yO4i1V
JF/U9IPdB1TfU5eXaWJEQvkDPeq4O7jzHZKZPN7lf3ZOep1Bl5t1OK3of+qbFxVE
WsSkSdMgCu8vyVAgA5Qmg9mASw8crTxLXJkcxf0SGwBeTYgvYh6ltUHa2DTHqqC7
cwpLn1M65V5p1oXRn09xdD3/eyp7rGo7qBc5Sta8ftvaDNPGGKlGtsb/xOCPtq5T
O0N+Yb2qtuUAhdkv28+HKog57v9Vz+qNHdDnrrzeKLZ1ApcNqjvZ1fEpRnmsXQiG
bZAJhzbwzLjed2nuryJf/gdNi8itvmYYVrl+mDIlMYUHwPNQcQeG2rV/+S45reBr
VGGwo8rJIJHwEhnSJ4Pn99UMltnNq62VM38v8XdYarmY+e43kTqx9uJGXwVyhPAO
c+wxDyhCMUPOcc6O7sH5JDa6hx7K0d8lWXE1Ws00UxDNA4CRCGvj0uQ7z63d9ZsR
1ddwiLFS2XYa5s/A92Fs6gNZs6iTb8RAxUrPL7QLZOeHDhPkwG0bfA2cUN0Ig+/j
2+Gvms1nY9+qMsINooTpFet9yx8bXleFa/i0+hovEDLfR3dWc+PahMfzxxkRwoNM
6lApe0VdB7fd3k5Nl7t/LlBP4QL9rveFegw5XnFTWQis8PActCNM1bzcvX8CHbjp
cDFZ1qNFddbwQdx16Z41Ud1xKyKeGiV5aTZIp8zwQGl3mb06QXnfjQeWCv3uXJKV
MnOAD9oTX+NirRpzmHPCVbp8x1DU7Z+VTWEUl9HwllpQ7037R2sSjMHXsBtCvNwT
L+tspyS5BkGlb6SzT9iTNehlBiDLdHpGNDh+INfv7V8gNDwtrhBwvKLt70HwiWRY
Sfe9J8XEpawZy1rW8h42XBa3yJLQBS/YgwFIQBUvyOlyT/oWCHh4KS36VQfm+uCD
CatBAChCNgRGRcr6A3BZXtz5Rkl6pJBhrdFlQgqaOL8xFZnUJM9Ilj/JvSbjn5+3
4jNq7oUqG3+t4bSD0s7HvAD86IIf9uwV2sRWYPi0x++pppNN7j3uL9JuWiqjocYv
00Deumo+t6H5SaMflBV8+rEHmv9Z4rR/Wn4pCDypgVr94OcVZD9Jei8NjDncvt/8
r3ocfDXkMuJR1n6afuurfApnSkWJD2/M5MWhV8yDWnutJGy9amqw76+2rR0ko2XV
aASS8+XY3q19OjkLAyFBHUoRzYUvehs2puIDB2V5ueh7a8UeBR8rdvgzeJy82MTQ
irF6z6W2/AA3h51Ghxq7qBC5kWSACrMhKxykM9tE07NybCCcstz/QKH5WRqHiY1e
ZIHTJT0n6A2eaNyuEDCgbn17AmaKTkRDyrsJzwqF9crWauiqZj/WETSlPxNMjMl+
5sKh+Udi+1pHyMFKCzwgvsoPx4SViIYICyBmvzrrM13Ro6lRALDkW1hSA98JtJLO
vF3uJQzLmslNcPhlxk3RYbh0WaH+wgjorp7NP0I49xFwq5fk8oo1x8gU62CUpt05
C3/Wf9QSNogH5Bv7l8X8On8823vZfD7wmPWqVSOhFrz67fuidR8aoy16JAyFVlAt
ggMk0zrcIM8C129IrxOoLu2xtAMQVLW8/5+HdnCRzxbgBqt5md+bjrRuqt3Raznh
o/79lqCGEooJLmLm8q2ItyrEo9iTvr10i+ay/5OrQ9H8AVP6VIIxSnhq+xsODxNg
k51rPQkzu/O6pQzNKUPE8ZgCqKS8tkiQ9bP/mv5wfnDWB1hOl50ROK35I+xLisIR
QuX92rYFS4kcshmrU7u/QlIjYicQZGRUpfHn9WsTfdv6+dcE1AfdCRj3okiMCc9P
+3MJHBB+xScZJDVORg3SziQxTHIHd9xV5rMHHclZ0iR5TGoPx54+ofhaI3dBZze9
3pjLkz9ou9LZjaIUSfsQCVJsvkkzQvjt0FoWt1aYgNHM1vT7znVaQeHzp5B1LBtQ
AUa+bXE5N5tp1pRDJ/GtWwgVRJJyKabhM6fTY1RCrUtwNSsP++R47OKodAPoWpGw
OsPweKK/lx56R+I6rXMG5QUFXShOTMYA26I825Vpcrm+4v87u6SPOcODYCVDVifO
ZO32HMgZu366ax8ClxMkxPMx5sahrnddMkBpX5ILpHcDo8bO0VdVmiE0FnE74oDV
7G3lx+LcdtW9OpMIKNT+WL2IquEdkVMm2+YmBY2NeGUfut7HKh+GVZM0e+iFNvtM
obXysMPZGSMvIC6vAs40owI4hfdpd+ZwIMsqAIYXQq8/KXLGzbb/PEOsoGWxyHgB
oqXnu8slNeK2WU545KK6RYAFlWz8yIPH4GRAZIAzuwEKsR7VBDuPirnaacwLtolh
g9RGJlfCF7O1Y4H3F8jHX6FLUjvSL12M/k/2mLVri6ExwHH5q20bvtN2UXx2mEgw
CyNHByMAKGz8HdFDqF6MF6QDbECsbFQ51nPbFPIna6qDYulI+H8fAeAGbB5ujwkb
xj1pIssJ9hA8K4PVUZAh1AVnVFC2GcgCM7FMy7OxAsxxERhVcd0ADeGw4NRx/yOm
8/5d9eR+mSz6w6AfAPL3d85z1BocVncghTvhX+mj4UtqAwmOrmssZJQhUKQjives
NRpaif720DD7gKFyy3l5QCMD9aYYzwQ6DpbuxLikB1FaLo8zTjfen2FIlLYEZpkw
ez2Q9/XY3dF8UkhASnKr/LWDtBb+7t+xp+4hjX6B1oQogj6yY1Pm/9rNes+BpZkT
FD5fya8qFbtij5+yZ3PLrhwLUlnoYzn476TnF57G/or5N6djIxarOMdqqAEGT+qR
zpbQDtP2Of5fYJyOO03dciwHtPwc0YE1fqj56aOAw3/0q3OT5ErRRe2HVHfXOY7e
bB4ocOnKqMMVW06CoCFUp4d9ns7jivBCsShMc/WuAzm0Ium4qS7UPziKfc+kmt0X
fr1i0e7QC9YmdmztI/Q0zNaktby6fQ3tmIGrFryFZqf8hOgOJ0O/qqyRyxiXrTJo
U4stZ5qFpQHpWlIxnwe0z+YmtBBMTRzFQY7+Fsz3dOKtXGXRvhKH/cGSGLebrXoU
scBjdc91AgrSc4s3FSsTLzov6xk5k74KCI0sDVZhWD2nXJwZSH6Thy3W1GP/oAu6
vDEHl/79Nv+AOt3gJawLfexONCR0yb0y0fqWep3xNyoHnoHVIXm1OhIv4ZiwQP3X
1Ehu/SxtJMsnC0GPi0i8SShGUYfRgsYhBzbNTiM31lf5sAAg+pfgQiueLhty6LyY
Kre6sbkh8XXOeQ9Kqpxc2MsDmkzIlfGJ01Zj6ILqfyLoMHl4IxNVDF1wXYo04gv3
agwr8BC+7sABKfWZbdYNCVGFAYaJoNwePHPsH0JEHmrMYWc6llGAi+r9kAR82ujh
V1at+5Jlvmh+HxQeTC7p12+MZKOv/Tvsw8snNGm8AW1CiI+Sl4eMqB1PdU/Rx1AS
FpR6ulhXrsnrCzFAU+ESXdjkRL7q+OoAZF9NZ0l+elCA6xIVV2p0Mtd6rITYAPL8
pEIjYXCpUCSzl0HdZUKp94sZnOrQ+OVsuCHn9qb57G127MMc5CrLEr/ijEsCuLRN
BlLKgszqAIdn2xmoiFoeVIWQ/vaiP/wM+gBgYNSPevHlgd30dwFuUC6aGAdHtHSz
7Vuxqyoil1OssX1/2oSzCGtODT1tijEkOmTMpPtEmImY6bldlkKofJAWiMHXvSJp
7N7Ep3dPsxlRDfCai1fyTds84HjjCQgK5nOqRWsGLNnNhQ2D8jidkZuKgPydImaA
y5JBt4ef8+tyVaaV9aNLlbuTUcekET/4MU7VgG41g+4kv+KDOVxQOs7sAG0E7JKv
R2L+Z7vSiVPTUaYOka9aUy5qw5ZqlU5N/lQT9H/D0riFa5KNFvBgGGR7Mpy8m01F
hEln440uXuIRCpcgZLESYqmirCFFnDu+herTkVsG0kCuqqz3HrWT412MFlpU1BMT
6xmfG54oeicWXAM1n0Nkswvdr31+y2n/po9dG6iU6NMM0woTHjEQp+YgZfA8vP+f
1R1paoDWXhHFRNZAt2P7CtFRxebDw/54YvbN0M1xN9G7dm+gcoKRCehgi6xoNeMy
3p3bEbNxjkuiE1or//ZLjRb6YHEwtg0/wMaZ0sfOktfQ0svmIaT+9/TO1S30T35H
eSVNiRX3RNQ+BfcFe+K6+Y3HAPUi+9lRQ4F/3X8azrLylW233OG2obNavT3OaEr+
VA5uPT4v2iMpNHigL9nbv4jW2KGRfb2io1/CDto10aUeKxn9TgWt3MVioGwg4ZxO
9ZDFwY8cPZbJCiU4s8b7qJDPjnK9vEBcqFlwawxNbrE3cho+q6fcOv0e9R1lwuLf
t13xqN82FX6j2BYe0HhFuRkqh4NaTHOE9EQBF+TFySrgFK3YPmAKVgeikKYKZcda
pgzko/4R8xKMQxD2i1o9GvOueK7S1RFCr/ITG/71nFXp70jgFA1qsPChbtEz4USi
BCHEqplm4OA7QoW8NU+slfkJhd7RUnUIv31U7e/2y9IfUOCcld+eYZmpbPsQ8Gm8
JF2a9SXnI+26q6C4j/YUz+Oz1/vJsBnU4boF6Jttxsiijm/OE5TuCX8NoNvRKeAf
rcxRXEHJsMFMZqXKJcMSq2tWrEVCjh6i0YA8t8SbpIcznkCJctxIc8Xbp7JMz1FV
+odU2HRVaKwv092NENA0PatxZeugVNBKbNk3dvqmTqiwschBBHmITCB7cb44AkP2
MK5V9MTnVW1Gmq5v6HzA7j6fKBiyfiyxUeOlYk0xOUb7D0t3zwqIQc7d++IRqR16
sFSFK8vMDUQlQR/mqMODuSZWpMg7qHEZgz9LXS4VkEDioxuYd2+2hByAyRy7ostE
UfLRqAbazQEOnU2/iqMppMDnqNbcDYhrB9RAqL/xf4MSJSCpAd4uO8vo2KtItZv7
pjHr/zrpQyy7Pv2thgb8001s8jsK59z3QEk6OtESC1Pcmlsy0mKtyx24m2EUE6hD
guncuCOdPhcggKrGuYDNvbsUb3fWelgwuEb1NtjQwLvySng0UidswGd82FbV4R0S
QAetokSv8ttf+bch9w9t3D1fToBi3SrZzSmJsk88d4wo487qn2VK/o6uXkA9ateb
QClFWQVzwfE72w71QHJ1d3LJuPwa6QKZoHSWXq/PeDHHWdNyJ9IAz53ZdiDp3JOu
QbSbVADp7HHLj8/gWJYvPzNMyWQa1zV7pRcey94QxAyj0JvTRIfX9Gu0A6xfIFM7
5yhbuC++x5IxaEXQQ4fKjaYngt0ww9RoXplMYOzz915MKSxt05Qt72doxQxussHN
g0QVyGbw/zzhgwPG3cKLvmMdwRaSV9QfG/jiq61YpQ8vK4YoL8jxhOCCYnDEwU+c
194ky/oJOdNmQlB8gTex/W+c3Tn34GYqnLWl/eun5hmme4dPLtHEfDXByHwBdJvu
D0W8direP5E9sEw087JqVy8QbVZFdBjEFeqbw/ZS7cdgSJ/getf3NHKRPbPSOVd0
8DdcPyH1ansYzMa34tjE53mtaC7pYuyEm2tiuW/htsROr7LvVX56loL80BoB5JF9
NgwQPx2rplFRPrEVAqVfQkxZGc6vIxAuyh85uCuRzAcfkJJ6d18p4es5Zr+R4/b8
1h7NnHJ7T8Eeia/EeXVB1ggtBa5aF2DXFYLOfZX9DK0Ho2IeTb1f/icVaNf0m+Nc
uvW/XJQStqUo/a8lwH4UIhZMb73aXV0jFooMhRY0gSOOrGEoGuj3myBdzmw/QaBx
D5o1kYMFgq5g+y9mD9W8Q3tjBbikOuRniVK+TkAIpuS+KlrZZUlsQ5yliDXxkOMx
FFv9gmys3cSIfgtvhctE12Zf786dQ98aNaiimSxf4hWP7+vbWseYDEDCBaLwsxuF
BTKizZLGdGXS9dMlpHLK0k6X8TUFgYp+sXzTGQD6bH2Ek6MXM15q8kEppHU7xW13
r25rFWBal3/dz58o/n1jtpLLr+h9wHVEClCDSdRM/xEiuoDmd+PHHxV4QoT7YU6S
amr3cflDgUXa+VFZqzqvLdgpxU/qiwpYRxMk/N3HZ5NTAKwAWamoSWpdnOrMAv3A
FU5FCDgc8/ku0Vdv5mdksaQ1opKrXeUfd1gnPiJlI3l09RYXTcloNNMn+HSFsAQU
N3qtbTO13B7SPPt1rONsErapj4LeKtfoFPvHilUR+vrgJVGZhOp/2oEKA7cYjQKn
ws0KeJlURWAbgZWvX9wD3w4P7nZTxLgYgkYvulnP002jLORNgU1ocsronsTzHE4G
ydFKOL2iEpPuwUrr0jD+CZC2HKIzTdehpdq41X+tU97U7dw9XqfCe74dB7lt174V
SU+az2/V3aYpYosYTnqSBZQphVjn9hUW6Jc+NebLl3EZNI+ezRtk9iQQfawyyOS1
gsubjItRIu7n41F6+N8Pbo7kWEhH4DBuAMjObH/H4RydrjWS6J26V3XiPge8gOOP
2GL80uFcZNNGbF63CO0NGqM8NZv3kFrACjpn/5LEmq27b8YKyn8IpDjSB0ZSwsTz
hJIeJ1FFOQtvx7epRTeoQbw1+pDQgjeoL22BkeEKf/K8YxuPzvvhwjc0Efn6eXFF
XY6L0P5GbuKjExtTGlwHgLEIzXjWt4kRHqRalhGFdsi65Q60C0zMcnAdDOgDndL7
EldM84lrnJCS+i46ffETwb9jfa7Os8QnXu8WNXV2hJkYmXkIjF5fV9VOI4LLSOa+
s7/pseGj+WzS65v5SUv+KnuXOqOCYv0MBEhPxHGw80vkpALIAA4tGuYInBpkuL3A
M1A4sc+Dlr6bET4860V3nxDdDR776Zq2xRDGbQ+vQDgcf5bWPCJLON7FYnPjpkB0
ee8gZdEuhSVBlBbqiSAEsdqy9MFGdNR9iuqclsRyzeweKn46AkDjoc/IHKfauWQa
wZuEhW8/YYygB/4N8cHbVHfFpx2aF51e0Aj5bX/N1H0wBK4qMb0ch5JedV0eAWWi
5ZWbWuUz1HJzC2lM00KVtE+L4JWpPs5pswWPmVEdbW4hNinuNrQe2/A+vFkuBsyD
XUtzCfY7awA/rywrLEkiCPvTl8RsMgY/Ogj9M4ieoKpyvyoB3dEzfKny2G9vc/2e
A6C+tNKBQ/aVms66as54rV19sk5ve48uyDqDAvynTSRharF4FVO5SjuQX1tTsaXF
LFWWMnXlRXN17VTVD61SItQ5QhWxaq2yUIAjgBZ5lAp7omK0RgpclFWJp8bSnk82
lAHdATuxxiP5FS14tJMWK2AdzuwMEFgP6AlkwwNNv4kcmT4fLxQRsvbHnY2/MiNZ
2VrGTCRz2JcPvxQsPZo6rUPQge1DSF9OeMwURsTL92o2jOk5puA9EmkJTcoWp9aQ
/1csJoOZQe2wOK6QwFp4RnzcRGt0MM6aouk5SQ/mvxxXMoh52cfWQo2ZIU+VmN21
zWy2QfHDiq9ORUnsEfCJFpEnW8efIp/t4dmxjgJh7Lyi2dJNIwvLa86b7XjrXSwi
KA3WP1mtDavJ3EMD5C+a90+vRbnz/FdVBTxcq2EVMS9kwa7bnR7VQt+t2N3UbRHz
TwGlLgF3xyNMSSEwAn3c85Iq60RdHflw4EmmCM09MQMQmFTvIldbM4lZBBtC2YoT
g+zdIV6ol4A0e3SBdNXK66dKlXZ3j/lxKmhKvRir8pEruRe/1Ocn/hzlG5ewgX/p
BUiZ93NNRFOMsi+4gsi2Tqpx98tGLY3/bqjKSSkCjtxQZKdLZnhIsGCpee+Xlgll
vx3CUDQODtYbfYodStYHg3CvResRa+OYlOn8bkBcLDm6SZ736U5nfv/6NSVFnt6Z
5V5z/a2wgFtAdF4lnIl2mr+dKV31hpRTWhV51EilGzb6dqQi1OtKbG/Kew0LfPX4
L6aAYGqXgh7Q3BWay55kjDVHPMJN5Nd887ytxDSLtLOuTUT6Quukt/VI9+dqkdpD
E4dRBcdjsbaoC+WfXJPZT19h2d3QPmjYlx4aE3D+mPb99rBQFyfdsY0qPBOVffmg
hkA96VZbTdEeGgTDUFnlXusQOTdNZlPh9Dz2u8nTM4yf2E1zyVGKUdnIcEiRI71I
2d/0niWUjVdJ3u1Bmc5i4CuotySY9aZ7xpgaV53catXKq1qfqqHHL+hM+K9gLFIb
rzetK5yLVKsWbqdB2Q/pw1x03jsmJVzIjbziWWvG5aVGzeHqrtFt10mfmcke/pFa
0Ifuldd9PMmMKsyeEsTtV0jIIdESHZL4VtA6iHTdmByjdSPm/gebOaKBAY+bJ08z
YuCcEPnHynOOe0+xSjIRjIxYGP/x+AsZA1UxKLpXVP/xTQ9cxJOS4f0Pm3vHxzh8
1NYEBZKz6m1alraDKYB+Wac+9tzxXg7ka/Ljq6nIv/cn7n0bprANoj0sZURcgwcb
zyP13BhJhR039vH5z+MgpQx6PNKXs5/fanO6gGpKtEDb1Yr97PQeHHVb7t/hoGlw
KGII5PgctbczPUIoMvRFE3snMmo9YeQ3O2U3odwTDnhTQkwMBnMO344YAnz37tvj
c5Dp2grr2I6/MD+5CXlH+o9NGu8bosSO3Y/uIC13CEOZmM/mRsMgqk5c87cb6muQ
45q3QXCykvRNf6+/xiqwqeNJTz9XhPILrtyOmRv3BoLQNk/60XOx88jXurzQQPNy
KTX5SDwcvxJiMbrHwwXNig33vwwy7f5BsxA18WpxeUNLK5iDRyczuRlSqyud/mak
UjjtypH2MGEQUDpYf6dJDv4Gna3f1khFqKS8/hUT21RsQz1lObd6GMh0iHpud8+4
/9QajyFD0xP1Rv3snTcRBJLI+1ebsQuTscwRtQGNnL6sShzcq+aRP5d+lfFJaLqB
qq3C6DFe/dZ990t9wqroR83JfwHprr+kOMwNVJeTA9rrPMJ/CwOnNCyNmW+iZdQU
1w5n8Xqkt0xtuj9uJaGRG+Rf8YWFFEMGjtz7zpQRYK+qSvugiXkOkxZvx2MxHBey
yTSLRmIZMQ7D/1zfFAfGEz54MZdzSotWLjvPT1e6gK3D0ujlsmXWXN8s3RFzKOoS
JXVIL14GgPP7IVm8p0dV046ruIxRrQAy28+Duu7KDtMJFDINAl6kpbNkAEl7ZoIf
HQtzwqr+32V6VSQKixxxcBYl5mLGvHQ+9grSSJgTjR1G3vljVq1Y7UJ+TR2JxBvA
+fE76aD4m5qjTgJAgGmurHRtg7Snb/97EIrrf/Xy2huLOiP5S4OKSWzyvNVcr+UT
ZZIQoTvMGm/Furjb6T2rHSy7WoEawp/KI0e0/xu6vRu2vBSNmUBueWNz8Ux6EyIl
VdL7I06xcKePTipPF5R8f4bimJSak26nRg25UWBbetSLolWsjB1M8rER0vUBlc5H
GHi0xQbmyzPgkn5lm1/SDVf/o0Ck9DO8GfUK6i2WFuWq6mcSvSMCGm5YjXZozf1z
w2sE6uSOrcqZXDeKtV+1NQ74htXPJwjId8iJwIWzx/q9wBkl1QU0ZyDDvb4GXQSV
K6CDLJClfqpQ1eIGclRP2m3eVLt2c63kdh99y/Q7HAA9L2YLXgFj6ELWk1DAv2rN
KpWLoP0Does6GhQNdWC9Ps4Io8iC6bRX+4Lj6gv116h+XSTNrHvXaJ4kJU8tBaox
VOt3JwmvcgE9PueCgTfcp9N/8VDC38Bk6MdvG5ojC9tU+lhU4zTkeOyV/8TNKwh7
hVn6S8fpaA7Tok5s3mbCUq6xmk9EsqpEr+QJ8Rbc7A8uvvxba23N3cao/1jOVD0F
0YI544QzhXDFNvnmzfe0yjkhYgccERv5qqi20+sco+7MoXEg32X6LJdq38vKI0iv
YyXIYbeCNbFCzOAJ/Qw0yyMsMYeaUQIHWaqhnO6cx/b7ZnVAorAoKPN6iQurQOb4
gwZwwpvD/iQndDXFlEkiU4es1q+bSnL9wgCv9kbXsbWLbMbBLiLXwM41ruuUy664
eOujuamAVYde6nj+PFMFGPGC8vmLXx48pNzfEXLpjqDku1h4LnF4cOYckhKJcsf4
okqyiFQqzSTnwnsQESCRRYNRqRWnnMSSOZzXr/Y0akcC9bQK+XEomYhQteba+CNV
PQYXyP2paOk/AzAWK6vJ1p0QJT2y2XVUxXxypx/bENcUz1rYkySTp+WI2Z3ong05
4sIB/+NVSGMqxA4Aqw1Ew2T11Pk0A5KCHCcFumiLobffIhW4xhjjMQ6emJqVHjRx
F0FrTKtMTNSl4ZSs1Fx7wkgNSaPhDfAguz0qStv2ajkHVRbGhZogCGL1s463zzl+
alyjpu3+jYKy2pH3iDEIcPoiG0L9Tl5n8z6ZWwqYUwAp93OOzJLyBT/WqqejlXI3
1Wdwn+aomkkNrHEtGPXy6Ekb7FfG0Dvm7NDhTm6mhVr0JmejWHUpqkJH61Rcx0Uq
V4696gHnQ6/kbqdMpFG1b5UdjrMGT2flWVokDXlA+MiH/iLmL5sT2eUtcT1eCXHp
xrqlAyXp7+fxZ+X3/b58oJQOlsGPGHmOiWZVlEcMicMT+fLpS/2irq3h//FENvCw
9Ue7jPtpyk2b2e3vULpVZLElkPBe98hEpmBP7jLjdj/WeB0vZr6P9ffd5N1G6uBu
x3DY9Sefoa6J42WwzlRcNL09HEis0KcYyxZfSIMhWh5+j90cl9JgwtQLNeQI8M5c
uPARzONZGsw9s473+XwE3ulrM/swgG29bQoV9Pe4mpFH+28IXxTsM0L3FB/PLXh3
58X6qqdO2VSaCDL1Wmm6ExT6F2SmTna5qKPo75S7uENc65aNX2qddxc3W83ghLCf
gZ0BgnfRxAoDGCEhFR81c2UmgaTCAB6fRTduq7NaJvJP7t82Nhtkteni+mtJehF9
0RcLJ9cVD566tJNUYK2EpZe4AVvuYKFdaRNHle7EpiXjxzM50BppriHsIh1aXeor
nLc8MkFbxY09X44/2D4UFD/5diHNP7sgMPnc/MgQl4ROv4RV4uu59YAirUzMduq2
WpaAbeBZ9fcycPTiqJ5ZyghMegj5DZoHqrxpE0K3iRTKSwQ6LKHhqBAOcxWQyEHE
WbjbdBrogLZ4Hus3dGwmx2dpk8aiWkGyzjCQjBNIsDoSMqKrxyORpJj+1K23EkT4
uFdFTBfLBltbafkjKOMT97W0zolQLnORVIO0+zDMN6J88SD/deyZvRz2j6D635oU
/EBxTqN6mld6pEnjR9GbpijWjKPHlXGc8QQR6PdnagL6n4nUxEuIw8MRUjsr+LT3
7Cdv25f0LlZ0I9WeQLkUJgoa0FkaE0mL9zBcv9PDaKOHsum8qQ/7ndOG8XS9hx5D
D4wrFydif9gKD2sridgpxJIRC11ygnP0IUCn7jXSPJiiE6dTNl9QxSbIy2MOEnvh
Ty3AwcZ49Za/bWYAWrAjA8v/Q0LFAxbI01YvGxpa3JnoupzNjGIzm2KQNDiv3EnK
dmPQDx4CC8bQTk2wX/TY1oKfOMCT70V/uDQw2ZjH7eXETHAsNG4LnC4UfyGsY7e5
YmrxHpqq+uxGVo5hwwOFQHV+q2mKhVNS5n9kwDx/C+HbFRGti/zpDsRM653ZTbJ8
WLRje6ooEilRZYAFgRgfuniWfOxm9+qz8Jmwx0SHsI5x57UibkkNZgOsLfVJAQPe
VFoeUOFg7MRrIeF160pAMkV08NL6xml2ubJ0nl1YSfQ6fmH508u56T5we5BrBshI
8h5FG17Ew1w+KK8SOge6pPmWpBYtTXskEwaDlUcEjaUZfYrdNTptMf1rslZi7G/2
7K5VZTisZrBfOyFFQpt6CnbEPg2nFehxqftQpbDmYD8bDIWDpqYCd5324wivU4V3
s5Fh5rxie2j+ZaSzXwJvnwf7uSdtuQXADEFOtjd2lsq92l5lmB3iz4k02BgcLebf
Y3WjTGtUM9t/pRUOEhxUWCxJVc9p7aoZl3lEu9huehDBsCGRgL+lkBF2hWUo8sUd
TR0+y+Sm4Yhe27hJWaQ1cWCXH6nlLyTfuWFf34srZCXFGN6wVrRBkO5TG/AY/ZGC
EtrEtMsFfYkpSYHZpEOuG1EWA0jMwH8ETqdTdnzHYv68ydhXoDkVTb4zO6gGDQH2
HwQtK+Crzia88wopyYhmyGsayucp6MIaFXRaYJWoh4hUGj51TNtxHAQuEkIMuZIw
sonIeukP5CPRLwAJK0xp2wCLouT+o/dnfExMQ7zWI5sIe6+WacPRCfVlB92bQAeW
IMEvOSvWhJRsRk2BR4lUHamhWq4P8LrynVmdF+VXtPh8f5q1GQUGa10obSj6ccaG
hk6JXKPPGs2tyKTsyESyEJI9Dkz5E2MMN+08dfinN2NiaInEVZTaQnEVjBxQz4zu
bAZZlyMxaX/hs/g6hardBKbdiIdnuPtRkk1fpAbR6hDcAgi06GMfNCIOK72v+NHQ
rO2DMftCGDD9DZ4c/7sELrOlChEPzKOouAojWLdERAO3A7fLu0FuemOyk0PMcMTN
Nh41khkOiNaqB8Fh38kDx35GOQvgDoyNH748hJJsLNYCzCHxLFkX9j0vPLry6Byx
SQKSokB8o+OyL7TkCxVPqJIAwKgxScwr6iC2rXZ21BryWkqthub7JDXoa6GHciar
WKtae8NcErgOT7O5fGkOqLIYYoItwHDinQthXEoA/3j/qGQZHwv4yIHr2jJrWRPZ
kHQroDHSV+fenFD90eb9mgbUwZBYSMsVjMyIEKQ91jRlQ4zjd0n8eVfNQf5srl6A
HFurMgqYUZszO3b4lauwIHdKTHKaIqgCBziKrrDXplc4acK0HO852pHXBkOKNUe9
Rq6lG/X3poPv3koSRDtJ5GcwlIAJF1GqJKQFKbISQdk1wchdkfLNYs/Hmz3HuXhM
LpL7AMSAJmqCXXND0ahTta7cT4sX2SnvzchjEV2zHE2NQc0352XynyB/ORVMMBzA
eX1Gate4wtKyCFWCnCK8mW8K7SCpILjUElARY/696L4v6+VFxGXcXNIV852JzD2e
jvbbWWRAO8d9/P9+2bE+6rov28DZL/ewvOTOxeSmV+a/H5SoCsnYpm0FpNOSOsDm
tfrWgl2r8Inx4WuCr2z2Th0mv1b3q/eVL4xJ0C8p0Til7ZAN87mjbQAR1+M37D6E
c/kpTdEBzfFEpBdn1SGavLUu847p5ShqqoLHM6o3WSaohWkCth2UdSAwwdr3uMLk
iqIG3jiBjUsHiJi2kWdf8O76yo4TXPROm609l87rpwPyHcj58EWXhvjVG2TcxK1o
Xtx/emk+phpEOXltsoOMZeSWWW6cq/qbz0O9thTYfZr8zWVK5ReqMh3oMVU3Xo+N
RmZYCVtZ4LOY/aEY9POtl2oR56Bl1FTwab8qI1MO2ymaSY8rtOtw92WLFYWiYmZb
MrGJKfC7C2IFkr9pQTFJI1TVb0JddRVsjqiwNJoJ6oXsQG3GrEQGV3d2ExFOKEIT
xJGXk5wQh9M4Tdtdx4bRX1maW1yL8c85FODKYvnrtr0MUCJdsqW/XC8d42H++JpV
GZPL5QpO0Xl/r/jBbcREy0cazQblh6/I9dW7sp3GLPV36O063UxCSsYMnA6pI0JH
s2p+Q6YW/qUQ0a5/wUTFpN7aQpUTS7CMTlgefA0ZwlvvfAyDsBnDSNyPOWy6Cgol
A42ZN4JnNii/kTs8KGiefvCZLeqP9k3W1WXJ75Wq9IS1erYaAPBPgLPBAS5ks3Tj
+xrDcX4VTt0meeXFJ0gBNp9hXGaxodJ0HUDYmHQkBoAuM27/yD0SBJC2zGTUHPIK
1vJnCsgeIOl+JfWiJSVLvJ5BnKLFTIV4aEGmTvkHvC8eYP8+gZrPsmuHT/Egy9ri
nXmbHL3IbEiJAJtpldcm8UnIMMlT2JdXl9HdHQE2Gmb+OlbBdPJ4MzeYdk9bno65
nonJRFQNejAWGBllLW+SeEbRoyjbpbCHEeZp6Hh7bG2QvU9p+MLjsL5qSi5fT3KV
dDkgvy19P31n+LCjiXYceAjyUdSMhwxNdLTy2xHlaxInIwaPX7edxrOJv+ySt4a9
MTCyfkVxm0MFySuiX5EHkpNNrOzmF1eLTnAuIyDSwG+qvMH1c9Rk5ADJ8LMqRdd0
MAnogCX10VAXOFcPmknW2y0zqydF0/6/Frc3XW4XpwO/GVYrRnif0jtmJeQfgRic
wyPrnp/BPbR6hV/PRVZ1kZltK0qSF5qWWkcYfDStIOiBWVKXnmxlurWNSlR8XZHU
uJh9fZ3HcGPy9+GtFFksKGWN67LHZyxFtYcBBXvU6bus7QnEEyqN7YXSXcquMehZ
HH2PKYgosIxncDCW0jhu/A+nHoWymGBKkQkezw5l73JL2SWbM8o+owSabfSLGv32
qXZgMAu4aq+vn3lxRJ3QEf4nQ6znpOYaEZrA8nuqCrczSTzWXthmwbiM3tyfwal5
TgrE0V78lDN79rOgzy20OHW+Z4qufM8QSH/EBROe4JYPTKqSe8Pi20pj+d5pw0Jc
TPB4EuOjUjG5HoSR8cNjFtsVz04Rk7bhhrHw0gVneW+abL3QwpF6BbDRcZMFQH+u
/vQKs3Oms1FWrsaEVd5SKgxkmZ/rFv9mSBmoL7FXooIXo8RG2rpL/owK79LTOBLw
XCAZPMmmLrUGMHg5xMbLGEr1NkVEfxmMEqXg/9punRNxLHtTljcfIARF2irts5l+
N5APYkn71DymSYkPgo+DWP2OM548K9M0RKN/o6w2t6TJO3aD/gdcs/+Wn3OFbF5l
3msqxUrY3i1r2L2PTN9VF25KtteedH8sZHlrwhKQR8/FM9uhwqxdT1JBkuXzb2Kq
yzKpg2wEuMOwK9CrEl0ZZJNr9Zqc2xWPV+7baz4y9+GoJFXu10zu5o/Sarw/Fm9H
WJfVrZ6NC57c1xNHxMLbQtxV/48j+s2auQ3yA62SeUGY8J/Goef4QeBLPTmZ8ije
N/eCGfpR5fgftqvgDX8AI99oG6GirqYwrhWzqgOnUq6N2kBpfTLLPBUANXCV8GoK
OJ35SvcFko/if+13lxrY7gfYrii3kdSMQSmlbPFz/wYEzTWtDT7qUHODL7rZGw6C
4/0WMOuIAWN8V/HNH42U+INoW7R/GVpuluU+VsHRP0IuRVkL6Dc+qXCVhwjMkUgV
cS4seX3j8HMRXQ1Kp+HBN1ZnqlNJkkD/QFjazE0kQyFyA9E7lAvR2hyQ/bgEzLMb
xZdWQlc37zaZt9FHraz2NWOs7kNw3xoE4jZLvxVKK2QepAgpGAEht9m7xTY3Swck
+UjEeOhwvGbI74Gi/TkMV8eUJkRPkeQt202iTr1aD//ZtWhP7HDzduboRwTNjd6j
+NQAMpjPqjLyELK8zG2eLdPtgBRMMt8oi30oeRL2xYt6on6E8L/cAyIUK2lv8A/H
Pi2FTV0EbDnS/2IzQPZ5AeStUXlEWoLiO3gF9tMf8YHBEg966HD+Z+4FSw70aZoR
g+TyTfuEg12jaqUjKq+wJauH71wLbin0jG5+t/s7oYz44ypT17QDq5O2EohkyHt+
dLqDm2SCAoydbJXX+ZgbPl/hie5aMepSbHlBnXJWJ6JcOAyav5ItqkUpLpmOlMlX
d0F6j/DAckWRGbiCbNcsTIr5B3pdamZoZIGc+MP0A78on/r92I3BiEPmfUZzSh/a
bk6T6NTES502dHe3sx6L+T/NLMmnDJAwbDUPn98NgK9tw9+0HlSpSAZPr0sC64Z8
/szeRweBqFJjCmiv2wSz0Z7uClc4PyqA1VEDs2BAxlvI1fViEDLtg2RHyOZPLTdn
zhuGmL1Cswj5wYl28utcZ8fVSyTVuqEaTGiCH6KEct1R3krjgH1JWpiPFIfKiJQh
l/V1XMtFKNfxpgD+qV9hH/RlcfLcpZowska1tc6aYsddmebx/vv0uGIq0GohusZM
hZDFPWNEDOOpqUBOM09tXoEv8URjZDPdB8GjjSglTG6IkKmTdq2DgxchsduqiT5R
S09e/MmDo+MeUgr0+Ac9u1C6QsZGF5p3t5bQ3x7mJ10c3ReAuhmQF1wmaY0PcFEl
/xGX0d04MLvWlxaAZ8ZqVfNJTd3NuX2LaPs0uFHylgU1iiqk3vMY2k3lfgrFDjtT
KKsD0T6neWVo9csubSropHI/bs3/sCNNCnpG4OUuCyxGvSgaqLXqgUtP0Qsaaave
S1tNGodpI+iHYkMB8T6rufBWbKXoC+HOMHPONuLuMlzKhtbKc8U+2JGdbyQRJIHj
YbGtQuVzkqq7IbMNERFzbc7jc9Glq5FlfLxWLjxD5xoiYwCQPC5LHlA22hUw8BKF
vGGlPNz4U0vHKcdSRSsw1U6Md6zCyhgK6GoA1pc7DK9TTgzEwcGEhAWAQ1C+7d9p
drS/JU0+Af0FBxERVBXazXdyHiV28Cju90z/Tia27N15mCIRmMuvRglfKD+gMXcH
1sUYXeTG7VLhTtFuW3ed7UQ7Iy54UHm+XV4reNCdbj9Hwk347DBm3fJxmDqG5o7C
RL/9ItkqK7DnHrakv2xrnLyoxhC/y8q1Hmigd2iYam0svUJXXw5tP2d2wojAXYhU
mkGcqBVQI3565QbGHhVwNht7BasXT5mRgTpzwEUbip+bpOplZbXVQ5JW5YNP9TiD
fm2owluxUne7yGNNzbmbJ4il7K9jbywOlJnuu8A5FCSjlFZIp0GFpyNF0F+6c0Sr
DH9Vg0mObvMIZjeYUugZcbkIEG+uDE6h9Vj4zohUg0I9WIGKXdZFp7KIkixS0PCg
X9Zug576/w/Q1cqyibJtLsfRivfm/EnZBTgf3A1ESv5eJ5nwMdu2HxY1o8ucsGSx
B2k+pNBVu3wZivVBjAnCUescqXbIUDBjqhXjojf6VSTl6ZXmIl1hMd7MhXz0nwcw
e2kC3vVVX19iBu2wMuGtdkN2rG6TX3KojH6PsmC8x12i3RQtkjTBhzPGVXgVaHac
CNvI3jtUo9dlwQ5DhOcEUkXlgR9joVokMc3Ee8qcWRBz9+pl1XO2534gt2IGehsd
arMI4AJ6y+RsD1j1gO54HmehGiGunJkptIbGbmM8PJQ7BJ+mL3FBLELZtHw0xEOb
TMmW5j3cw6Dmjq2Z5lOhojIfVGvi6tNnCBBGpIA1EllQgsH739bE5LYZp1z7/Op8
pvg7+M5abtUzwK+DRlUdPV1GQPdguvoZqtWseUaZdgWMUvZfADlHQaCbRdAPyeh4
Q9SnwyW2EcfNRafwNaAXQdKQNVglhlYR2ZFNUXV+4UVSTFa8D5rHBfjQqiilj3tA
GXjSzU1f44a2FUiMGItQu00ox3/j2fzewfEDnBR35VcCJ2grQqnbu+rtE53TGq3R
0yIsi3w+MPhTEPPKdunOq7wXv1I0AYlPh4JpTAW9jxWFEq7XtlZkHeB5Yu4o6RT9
iVcK6KGDjPAoZJwPam0SMZSW0wdP5LrjrWZ+K7uveANSfPhixtArRsVJRY46VsrZ
1qeEtADihNqEQtL9iVTc6xJgjqV/hyirutXNLV89BIzCIgF89hTalwsT4kPgIKGW
IK77VUU1vfjngi4bknoyC3PwpCPFCC+Q93uNJyaMJI7knvl3eMsxe9QqrdBoHSUU
IVNQRHicKmkdOWa5u0WwipVMHgfrJjT99qcCVCccPRnf+09RpN3HanCph46fGllh
x0nrrdw3N8zEbDRl3R68U2aX2q//u1io25AcNx/DdxnwsjEnmO435AQJ3be70OKA
S8cyXw+cVH6bklnJ2L18dtGDKkpPDsXnbGRIhJRef//3PUzGuaEART4EWdB5aAKz
RW0ra7cInfbMYO/qmcgpwmC5n3WLMktTejHYRc9aMthZezy9w4INwQgqFLc4gRCj
pASCzRjf7u22jpPnNf3Rwm1EsK94gG7z/9z7C+X3CNHtpVDcRaF5k4HDTyg1gEoS
GXWdzjTaR3jNmWuN9OKN9V5+1rIiv/hzgEYdmaS09elICjkqatGCa4Ow2sMs6cU+
Z2yUbCn2911U3V+xe0AgTl72JndY6q8QOJESO0FuDnUKOptV2NigQocHNdjFUNaF
ld7qVaADVl6vYHx5PSgurlAIllLV3/iCiFBkAa9kI2MrnGART4ZrEOcigtm90nxf
VfDrv005sRZBIelVbh7jYlsGaG29IS1erW5N+yuEyGuT6Sfei3Ie5B10x3wRqKFy
96+1g6g8iUdFzH6iTyE4SzJkOLM3BbebsjxUsCEjcKZM8TWym12WkJ4Udzia6WdM
LngCtU7132MdYkUp2hc16nVyb9qQa4f2ZR7zZrr9V2sUcCTc85Ktms1hGKbig6XY
lPRE9SWIZhvsLicJaoZ92sjCoRu7tzL6UErXz7cRZyifVGgkc+a+rv+xJKs+6MKz
L8GrIuJs1hRTDh+UDQobFJ2e1ubWRLfuV6lyH/6Hj3ykDebFlHrePyK4vjjmyOuY
0/pUbhdorl8/XXb8XcaRh48xu6o16/60LwudnO0vjEk3wWGfSObIbPHB1+VkBgX1
9sZDfZqNJo2jAXe2GTNL5M3GA2JljPex2dRvHrkacG4wFkTMu9ieEjP4bSxpX0D0
kBzmwiJIkXh0PPW585P11YoS/94UToocK0D6ANpnpXwS4bWqxgthAF51jNyOYeXe
lnSxt/t4szN1MdeqHiZHm/HsUnOWQJmnz8vJz2UtmjcZZ2gvoL0+mhH5qSRtTi3p
+6ONyy2MUQd2omMfE1+40aF8hYYi2d39Cq7QAyj9iN5i0HtU1g6/nMy7kmZyS2Al
aU3Fn99ZrbLWg3Jzj9Rgjnro/NqrsZKrTruB8w442RL1xHeWe6BuyEzO3LbYHxxQ
bVmko+B/ey2LwH0XLzQu846uaDR9PGbeJbqc9B2hhLbjloKEFlfSuiHr+8sqTCQJ
ICV/pbWT4jtopO4DTBMkiUj+D+VZfKFYCKWtQgAJa1HyJ9FbPwl0qEta+x0lQzHt
Pgcd9wSUTLGLTQFDCdRMnnbzwlCsbgjYbnSwBWQKVlQelbBSFlYRIWGFAv9tR3Mn
q/DFoF4KJMx3USP70oQLA21yUA0QyOOEwWWABet2QrgKqCRzyCP0ISkS6T9tWBOl
cVAy3AAI9FSXEIdpVoE65xViruQ3/P63dj3hp2JgnHX8Ji1o1rmua3lCqldTVkNJ
6euMDKul94dJfX8G/fCUZ3yKWTQF5CpoXRQuZeoJK/gr94bIpJAtNkp3kZhxqtPO
fyaRsTuAbkClQAdjyiXanvCa/2nmktgmeK/PE2evbBx3hJ59clqYhlQsRB0CCM6a
EGYigR19qJ+R4klB0t6hurkyfA805IXG/VgYeuPmUncY+osct2jaEwRtd3wVK5ak
I78V5x/0n8hp5bQzKyIHkxMGK2Q91eAiKzXRHdi0UruMBm2HRBZILceIYEKomQvB
Fa742b7V9AlzI0IUDoxH6KoBvKl3moCccrgAXc/u4m6TfEpYYWxKqtTtkrzzQyCR
xvE/vkldG7hKD0BmpFT7yqY1PZeX+Hi6ICYxOACPNQZUzpLxOA+kvSbZK21sgdrC
GMOJzBFMfVbfWMpJYnrgt0X3J7wENS48dZqC83hs0jIQdjwJvh2oPHW9H8q4T5lA
9Eog+YJ7Ws9nXHnzsLIgHT/BQkGOsjDRex0q6yOce4xaO/oXiyifA+6UdQDczWTa
kvJRIJ94EDg3NjxVYp321AsrOshLJPlyAcfEYE/PZ8MtzpbINy3XJKcxvcAgvqay
B9FLVDBkvw3G4Un/c8Xhu0NgebDnQrYgVtfs8MQCCtADRSk7hm0qOhdEJQEPweXw
Rc45YyvXA1upBBRUud6laI6vSCs7MhA83KRrJhcs2ol06pueY2sEVmQpkh0R7GMt
5gK0LqcTnud7h1RxBQ3GmqAjIWfE16BuY7/nIXcuBWzkCr+AF+YcEyVUGjE09CJQ
/5BS1tf4O7+Eo+Js5m/7aIj3YzMMoklFVlN9EB4NLzYSRxG5aoPz3fZidWKPljg8
D2dKsKOJJk+ay3/bH5YHNCO5iRnwoGYnmPjPNh9FPP/u1Ncc1IhuRZeL4SwTTsfa
JXKqJ7PdjUSFP6LCn4AERbCR8B59kygYrU+BgZDlVS8fV7P9oRQZBElo3lTMqs0B
B9+YOHoowLZCIzD5f7bHp8plZa0F5vYElF9/fLf5ZB0q56L25OM8qrczq4jHQwyj
Tonmh9CrSpacWs1eZWa1oH/Q7i7aSmPbNTrmk82hLpBkhfdmMlaZpPL3waFtLctd
YDSD94yKYvsrb+d7/4waOGnQQT+y7WigZ9LIaOruv8oQnPSmt+AErzclyrTEZyY5
AY0wxhHImogQZOsB2ZzjQuyxS3Q9GpHICH/AYaUyWZNn1/ksapH9WC15ZqcAlvv2
mIibotc/xdcUPJ0+ZHfhWctnehZRigfNCzKcMz7uKGMDZxcRFoLvb5l+QFZswDR9
K3x5mAooG2i+sE9+54MkjoZ8rIkFk8ZFVr/poHTb7o9PnFkS90VqQ131lo31JvhB
dQxeZegAv5kIY3dSWcspZb6AZkC0WDeuOoN8jz3lCN1U3+bZwJcMF9v2aZFGxdn1
KJ6+SDaOYG7H5RqLKl6J3u6TVhJ0e2HLixs+ESC0sfiAd6lwWefU8mtWpTzidyn7
jZNNwBLCB+kw2e/Y1k52gN8mSFP5gMgxGnPRpjckfBXIhbEUWkNKLTuHnl0Yqov/
TyRboAW4q9YTobmgixrA7I3EXzTLdD+9GV3VKEkUD2c3ta3I8n8o/04hnN3dcSEl
GFvIk602Iy9sr/HfI7Tp/5wCFaSAxuX6gRyQv2hPaVCz4YOoem4bV3X390rcPS8s
39xpX7DPi3MwYT3qwu5e0oChjXBqp0dhmEvRB5qAYoeBkV8yE9vyKm2XlSgpSkBy
+g2eWEc/aZaixEu/bD0Tx/2aAwPR6npcOvgub6vr+Gx+8saQOsJcDw/QxpBbej4K
EB7WlLHI3iplEKGnadC0o4x+a0v008gay7cM3USj3A7aR/HQspShtOdR8O3ruXpv
WB4cX9/sySSOgmwDV3OYkQlZE+GJyozAW7i8K9izumNuVZAMWqiK6aTJmlzVBbhE
oIw25fA3bziymKfIek0aqvmZRBth5ezrAPdTB1HoAQLZNJg/ACjkTfk9/mIzErZR
8JZWXGAXUUnsERUjXfjhl8UM08oUCEtGui9LjUxlNNANyhgjTliAKbKOsfs0SNPG
P1qzb4MxkBNwit4LGQHXnw8IcP7fmLo/MWKN/xM/iDZYgJRWcaG4QFPR4Z1o4KAj
QGorv3tIm4T10+6t44f8GikMiPaHVEIw4kUrHln5DjnXpWP99MzgKnSDKKTO878R
chcZHskTBoNR5iRx7LEGZ6NFMiFg5gr3W7sVUu8+ocBPZL4tMFSgM/K2KUpyoT5p
WdgcUs0ArXNyLlpZfIXve1WCVfuJiwqdZwf5HPKQLbVUUITgf0rPUSJS8ZwQAzlL
r+kqmbKstzRO+neAOiPT5VDNtyv+IUAzLAIOxzHJ/kzyeP5zmTT+EkToESXgNkoz
obqtaxTtLOKR5PSQNNtoqAvS1xXAvlnUBs5vQnQI6abEzwKGfmuN0Lqw9sQMutXp
irPjevSxT18BED6DePbI8uTWsFujH3eeDjxh7HAHStb7bJtIVhUYBYAcnUGUZANl
qsRUUdRUrGiBPJE9Yjls1Y92EYIYAMciJLq1QC7GwLKHoq3FVm36LuyH9i4+ylRQ
AV3SxAIDgZksEB6zfP4LyNAIZwln7pqh8bcWHDjmgUXumU9UEdPtzLyaJz9Lduo8
vJHQ2xvik1a8voRatLE4mntLmp8YwO6gpBmvh7uo43jKK94e6IJjTvKzNzdcg0uu
n8loEgJ3GJfP5e9yJqn71Shz3zqCzbnJ68QJIsJQE1d9gcRHWkD58NsFdtNXQ5TT
0PcoRCBkVtTSPoH4xxXHmxqu2ZH1OQ6q+5fnkRxIPpkoRQKCRnrRH40O2UHFThZK
aHH/xjhb2wy1mhmYwoO3u6ZtP7ehhBUB60Nop+D+Mt6iJbVe7xSitjJ9DlzA9L6+
xbq0Tbx6DqdkHe0GWsnqsvGcPhA+0G5kEW3Oq4LOzEzPNk9IHjYUK374k3jH5d/s
gXNpu58+hFjytHj3pFpQV7vFWJ0h/CfmbiuDl6QXZikFQGLmCVkdW2KJ7Oz1Ln8T
I+p/uUlTFnCHz9ZoQHvHZPUdY+W4i1L/jBT7AlgDIBgwQWidfNmXdd9ysXh9Q8dk
bg1mYrJkdLZoajdGpUzS+ppwRkVkNK63t10vy1s5gr3B0CWD4fB/m7PNV2mLzBap
5Jhgc03mZU75hhhJrKtGzxU5zlr3WGJCJ8BmAG6Ji2UnKKI6xQmA3C3aCq4+7lKG
KQBOZdEKr17xILLtcBMjDoZOZNjGB2UVLLbsbOoHOigfQlk7RDSdR+1v94XOYQd0
1aDAtWSoU/CaZdVmVUSdv+5/Ss9IbAn5KBSLv6//KR9YomtFXHFWfbN8MbwwCREb
fLujGlSkgPH6Gbm3oMemjmORT903cyL4JEOHEHw0ti/rgaREkAtGDXdPcFKU80V1
g0OykZ7lp1Aw1culI1S8UGQU2tmYZkcrrJ9lZDGHuasiM9SSN9m8qMufv+Quw/99
YE+ytLBQPRkpYY2aiLX0c2FFPIOJVcbUivh9VtuaKuhF/02fSuMjXpcm5HI0+q24
WppsUDgbu6BXcsii3D3JxiOkbPJX+5oN+lRk1GBPCR88aDGm9d0aUfxR7p/z+Og9
mQ8ClCmehThtYHOa6ZUw09zlsyfmT7uxVhVQonDX0lWQSgL0BaX4zDlRCjB+lOUR
l5mD/GlWtztBbf6gi5M0X6H7gO70fZyB57V/JCsLO5/oypaTeq3YxPfJs61l1h57
iIPd25RlCFxIg3oQy5hIhqRyZPXFLAobMCMfIx0PF1OvLBoNmAXardD9RVE2aVXo
W6VQr2LK8q61oXOEE4I0giA/qrrKBYhrJu6g8o9R9TFwm4BZ3/gQz3TsAx66tyNq
NiGaPG4ZapxxJtjHUFhioyWY0CA83JLQY6Xlh/BK3NkAf9arYLDjOW2dFuCWh1tD
g9icB4VeAyXs1eiWDnQC4TLRZfzKch5nFcK9NwhJjMlUoGLVa55ykGch3xTRwIcR
8AZqGORo39NFpkulnC/VS94LA97tnccWBzwHihtgEMy3NfvOtmAK91XG4ahfycpc
+3mlRevoKA85O5ZB3Jtq+KdIs1IgbaiAcpl8tZ6jsTq/mD0ZomAIEoRUy/HoUUHm
NDMXG/X0I4ZCtLyqimUbAbPP7v7u7CG5LeAXW4awH1KKJ0c4Vh1sBKjM23HukjfA
MrmB9B0bc3twke2xTt92beRIdzjiyRC4+vC4PhuWeSqJqBM46xIHdECU/1UqEqKP
RHnv3v+6LKyI9TOXo0ASBZ9nXxDFn4VBVrhYKILEhC1hl20z7em/BwkWtTCvXAcp
Giiimk9SBJLq5XG7BU7EelUR5mZPOdFK4iNCRky/SO1eLcBVJqKAjfPy0Jd7uprT
0yFhT8GRNB+FCfmVJ6jzrECmhwnoOZtng9BDI7WPx6aQlgZndAYCDuXFkyx83no5
fJpkBvJroM6Q+sQ+JWbciF0varVN4uYzcvxRbbeIg3sw4kM740kIiSmieKgneXxL
Njff3ywDb6K8Q/3eC63EZZG+4Q35R3I+QKOjVOlJhnu7NR0FvOioOreS7/gkccD5
sA+3RXp149dTjOq/32lvTH2ignXqm0TG9hnqn6Tigyru1Dut0xAVr7duno4033Yt
ujUolAQ3mEEcJLA28Ib4Khnll/3yyDQ+NNnjAVcunF5vQGmXDiPecalKXcMg67s9
jz+oXSWQ9zej2fCjso0G+b+nF7f/CeH6D2EOlj7EJNGpJKHkalu0w3Y4pZiEn2D0
DKRaHktbbGBjzDWQ/D9uMyMateuS3wA2ADwfeffrCQaD3U25oeyAvM4tX0Ffbumc
Lss7YJnHYQZWc1O5q5f9uJuqIj+idJAd2BmqfB5iJ+lAS35Dillh1MqC4FBexoNn
1Ny3iRX9T0MpXAyJXRLVdZg9tVrAwnjPhXT7xxzQjE1UHVpxMhiL3WH3D8fudxrK
820UN0NQOmq3QBZRdY0bXsMlRtm7MiMXt8nTf4KIEZucqqsOzLtX3sPrunHQXKwd
lh3uX5/D39L3x80ADRhztweX5b9JvNCx2hxpdmqg6/nshHpzwzAmsJpZwRP/h0Wc
kLPOz4lzOCquQSJHej3GeaT2Ns9rSwYOUu3NDVozJpCGPvi7gvHjfQXB+SHcwgB+
K/YOqZgd0qW6XloIPHbTKBi8PNjxwciYtvwRrpJfnAqjh0VBZs35g2ewwgwow2RA
ZZLMkcQWsIArlIW2XnHoHNDiaVeXL9TgUjF6pmSV84h2SEQXKmr5t71hobJgjkJE
sHzwdxODoiE4AfqtQWZRJoqtNDFAPBgbd6xeLybI88CLnOYyu8vCygTzqoMMZhKM
9nCgul9ALq0BeP7CfynpuZn4lBjn42VGccuYLga42VZ8vtrR1b3NiVNGxh5ignKp
MDxZs/bsoz/WkevOatAEmog6GKSLDm2qYr3gM0WylD/VE4mWtO/JyriKIB0xpVkE
Tyb05dq4b4l3OcuDuFCt2PhFaVVyR3oZSETU29AOoFgy4a1pYYpsGrJSI8eNtz+G
71xg0/a7KaG81rk+6eBQPsz65FvIYz+hzuB0vXG3CJO9ffQeYo9lUztk7UY1Rn9n
bz1nxIznChNhMqtsWM6rA13/Kz2JK/FWDa+Ipi9Jvco1ZrxfxXIM8yzyGetsy3hI
7wvae1UG3hYwYyaSh42VPJ/BwMXrOuL5TuHswnzQ3bLRK3Fp5k6PneFTQCUb/MSD
qOl1C9Bwsz9frtXvmifskgulWisgmZjBOSTkR/n+clvuZ2s3zwQv9TF+lqCDcHrw
NS2ZnbyeY38yuU86UXo4kFjTgB7BYGv8C4N05lJ6z1eWq2DdqE7eSgTCx/v+qt6s
iJ9DTfxEr2Zs7ymmIhm2B2qSnbbOJ4H5YAbnlQ7kO/5fxvyEu8SU5q2xBEIuj/Gm
oWxX3KzyUXoB/nqg5wA3V9afzfKwfwt1RZDGDfIiGFXTXt7dWsojZyzoklOs1Gjf
ukC9gN/ug622BHMZh2vCBL37qVT+l5MBc0upuBiWficIf9YUF2lnKfDjNeQiqOz/
jQhsOKQJ0Nt3dZDfebaDwjaxyDhjAtOW3pJqNuGhI+BJHR5VFEqJK9+LVTZJlI9L
QEriWaiPdT8gzZHw50H6p5LGd7JPVdoXa24PQ7FTy1baZ9B5UvHeNJDU7OxXeuBk
ghiIlunpr1JaLF4chJg9hf5jmX7+8emFfe/++W4IOCZpGH95mgnNFBF/gDnMv0yz
jPDA1IM5vaK9452LREBCS3HIPvSeCrlCsQ5AW3on1XXgGSMPVI8GQRFg4bWZQKcs
wZnJ2KL803XUlOUR6xGoyE2fXenVy5Zk3SmWmi0XcU7e01mR1bp76T3pS2SHSLE5
Jk+6Vgw6emU4M41i+b1SosIPof6y5W987NafbDxaJwP2q3oXPqZ2OOIOaPQDdvAE
Gj5rHXvyzidIzOG8XX2sG6j4ix8dLyMO1ILpGwec1BqeK4eJhLWTen+3n4tUymwV
3gsSIQYH05kjact1fWwSQJ9Xeehuy8fqDtl+Xx5erNFWTrtMOxfWaKYxYWA0tI/o
IWj5Lbc2IJLe/XqIQzvb25eeGhP19D8xGFxvLmrHviaT3Qd6WDbQzaZEMnPvFoQ6
rtJV98o+bL6QXUHKjLQOs/D9diXQOJCZF48dfmGRk78V39r0K+JRwt0DBvrqZMMB
EXsL30Fw5REi02aMVKqPxzg9WfCf4IXjfTF4r1Em2HPAuSueVfiLg0Fo7RbmFOWy
lv6MB0G4b99xVdQd1fzqjglmWHL09LEWoi2N3fhNEKX1MosaZyXIDY7l0yCw5Dyw
6Cl7dVKBXDChtQivcjN3Vo7veM9lFNvO9V5zUdTUHT21AgPLjcH4B8Wf9nxdqR2A
/ByNEnGxTFVepjFTK11LjTMsUqHmYWvNAThho05Ta/SNkMw8+MPF3y4DJ/SR1DmS
UsR9bEZ8R3t+1nxJgmvJj+dN6u62+cxQFZ0VSBFgwLT/mw38q0p5QqsXpxh/mHsv
JnZiRLqGjRXjgPuYP0M3Sp65oDIlZdVVIwOT1nnsSq56FB5oE7Cln3xeBCZ9oYuX
vZToHNXWG+GiltIjHJbA+/pbWc1M4n8Hx82BDXY9vl3kk3kEdf2nPBG5QbMlJ0s2
Z3UZd5vmO16V2tO/vdrRAWVeZV9HUuAd04MT1cogbF26nuzCWY8Elco7hZZo1Teh
XBXyT24d7SIZg3QsLKKBymllEBoERZW3s/fn/1HLxoUsT1yucn/LmQ7+BptEN+X+
TfHAzN02fp+UAFtgMQT1MTgRR0MOuIXLNjuzkBiZlmmJH20UTvV+Gco2KoIB6bxz
VfPcP7/DLMSt4xHj0yVgYAKpvF8IYe1V7fTUwDsTMzG4OtZbFEEShI4q1st1ZyCj
UdtUwA6tX6VY0xdzYBDbeiACSFmYJz6yiNDynJoTCOWi3QF9BlRE2Zj5+NpsMwGN
aZA0iA8OsgxLz8p5ffvlg4YnX3d69Gs1I3qcKcVBI11hBOXisW+ZP3kdvOMLRgW7
r51AmTtO7bvcb1aeuqIj8ccxxPSXaOBnoR6a1fX7rrrzJ/SVenXR7NFPdxs+GA05
CpoKzUvMvIbX3YD+NbcE0S5iQqlvKym7EP7iRDhZWROS9uBpiAg+nq5nEYkIr8Y9
FBFoxV1ziAks/KyqX1uh3BCoVG/XqU59xDOIFbn6ghmJjYkcmThbRjVeg1KPf0+A
w28f0P7UxyZsQZ+nbLM236GH4yu8CdMpcyxFABJJX1OjdT0L6BzxtG1sqZHrc7K4
eTzkb60DUWu2oeVuZJo3vFfUKFg2sNuMMNBDvntAz4q3XGjs2589xoz6Lp5M9kOA
8dkIjr/b53ATe6d1N9lRn3Uhbv/iIfmvuoJNFK2y+YkexBWdXeotQDzmRS//Sa+N
4zUPOQkd7F276VWsG9ooehRfs0cWhLBhaJJqMerDpbrkdfKQLxErdcu9fqOBFLYA
28f3BI7z/mO1zOWjO8uWVLUGCmOVBkG727TQLoNR5MkEg3PDRWdAyMHzFDljzac9
jJrTSOqHjYKopHY/qfceQyEer8X0ZyAFUnphvd2qMC2Edos9QATZZw43LPiKCcSW
GnhLgHriKsnWhd5j0rleyImRv4L2c+y8ytpbIMDthUNYOxoOwcTaKffS0kAyBNN/
B5KLBKzMDhsZIKaHYLlf8kQuH0Gqf3K05QFbfr7WfO2/YcUycQ7k7igD5205NCJQ
NQEE87+Ry2Ayey61RbsVWk0PrvYBmS+i1R7MOc4WJFjpS/ZjKhwNQKlbO82dSMV6
esHt9xuROKLSOiuB0hIZnIUPK76CgJw/N7X83Ux6exnFrxubklfjEqrnzdYAQ9rI
8uPlGCZczvwUKt3d03t0tHAIAoENzZ+goZcF6beTapiZ0zh6nqikrxjcw3tnlGWM
KSG6JlMkO1Dy1UVV0NvDdCm1TlyxBYFeqsHH0VRxCI1poBfYCGBQwlLD+UZENFTX
rpJBgoP+IDk8BjHYlGEW92adZ3usYBW+biTYgxqI27Ba6RrDyNDcG6AwCJHsP14O
Rbj/ig7F3N/f1mfDrbmSoR9rZwXll+7XoYfeW2USVntv0Q407DXjdzGK5XAtS608
Q3mFVFlcrQfooh/dDg4Wkmz/N2ApbfZmynVrVosrLUrtG6mzpdc3bNfwVY3NweRU
Oo5ZwyhfKi50TycpA91RXgc3vfd2JIIY6uEZlcTSwIsjr1sxesXovp7Rn63a+sNl
XBr2pn0dAWnYWIYXL4qV/EQVmB0ppjj/7gJK/1ecOZ9c+rEjsXUbnAmTonPgiWHp
CcZQwxuwm+K/dUBo4pUdhfq2GCXKtg+9049pEZfX8cdUN5ClXtYS5erRcmpAcnvl
hDfoTTRsLZO0f+NbwJ0eSQ1XtlX9C700lEAaFA86UZ8LCKkCwUsku81fJeOphwTU
zuMdNMKWCQh9yLF4cYoUj6j/L3v3NCLPwZypaqYKmzaBzgLLRin/oTFMpLrBcVkF
FhVAu2KfANNaCVs40a/ELHDVPKiVmFYTt9Wofp+flC9WuXtkrW3mARj+IfCioFY+
oPOW22lQlt+Pim40CuOrwlaJp26lD1HYYBjV4bLklKqQj3wW76UKE9xV+K8UA8zR
64E/EXG+qOzuoYn1l2MjClL0j+18gJMEk85XdDTNeeBwWw5rvbL6nIexfyNuw1bR
eW+hKpozzaDf7oGkohsocIdoRQBWVLiyUkDJK34tA2vVtdYEOva+gyhRvv5Y/CBS
8Shr0AlQLJUbve3XoO2uRGlxcUeOiY2MriMW1uxrR9iSbngC2j/ZEAP20TCbvqMh
fnnPB6f5ICU8136wQ2H7PNIVYFZ4+ogRTuZkIEv/7aE2xiqKf0mPtmKYipyQx+Gt
VTD3ize6JEJg8IzwbVM8L4hreLBtNfyB6OoCxKR+Q8hZONV3LoniylqIs4gsXMrL
LOZu5f53HttdSTFAwnnihe2shB0qyO2h1kZS2ZTo4xEcmBC1FQWibA1miPJJEr/X
RhFM3Eol900LrMXQeT7zD6vrjn3Z3pfxMHqOoA77WnQ/+b22wp6SrmsFuD2dpsEW
pQwKZC4NFYeYUBu11qWziuuQES5osMdmObt93tvFxoSPf8t3poD+D86Wzp4dl+m3
glOgRlmftci+j0+reTtw0ALe75YDcQ/5mSV+AVksVEAK3Vr/lJGVInMfOBtEsBj+
7rsj8LZm36m1M9buDLgP+FzRkoXxU2/tbgz1lRNEGwk30TwgnRJxEbqS2h1uUQDC
4ei6a3y2H2SpLrx5qiU69CPnfUb5/e4W3wUJzufQSqJ4tgGK3zWS3AA4MG+8Bwg7
onzs71gzFVSwP1MMPAwXQc7Ngh1OvPTmSMqdyvV5d13mDqLhIRV6rKEb6+xYE8ap
kZsaNWF7yIokD7KC8n2j6dKo58fylWg8Wiu1TR2RJN/mEGNF0MOx2pF4ja1z64Zw
Wjp3gAPszAeVTdmfwsMEP0JvGNEQuyzM0PzDZy92J5V3YxF/DEt+9g816qrmc27e
AdHeQmo3ncyVgUJxg8jxgpYVhBziurz+oxRxaUnSsk+HfuPyCWyb/ZZIT5y3Cjxg
TzMPI7mif1Yt7UWCm53rgeqbtEpxAYi00ZHv9K21uKHJfHlFW8p0WqFEpYAfGsrk
y/Y2yuj313aVQDSAH9av4s1iNpNlE1mw/Ax2+0f+aFELCMv1+LY6ul/EHZMSja4B
yjxJN38sI4szZQPI6gdfPm8BdvHZsn6Oapq6L9Kbi4hFcquaM5Znkeprh+zDMxSb
bZCjE8ihQFuaWp3P86ml0gEV0EWxw8MhUJW07aaFV/P3GGeXk7OsEPWKWxbdWyXc
9tf/iyoxHfbws/rupeusMLBzn5x5djs6MO9TUxqvn8S6mDmiEHxEW4+zDWMD+C2g
8HQ4eIQyq3NG7BJyKk658By1KZxfOvl7RU03K/Iy7/OYixirQ7QZFHxblG5R8J/6
VH5V1qQBfGWGRbqF9J3qCDt9h937KMw4ZpuPzVLsOUiYpoOgfxDmfC9IAHyONkeH
NzOgxaMeeeBl5YI8zG+f6wmJFlH43aUOk4Vfras7PbaoD0Xs2ncTns9mzTpCZ/fv
EP0g1+WdCT74/zHde+7QjStD1pbg/gvVexS7XIGbbo+U61uu455P67F4G9SatoPC
QoyEbV0nnF8Afb6b6A1YDdlbbRE/xxl9B3M3y0xI7OwAZfz70iUiJ5N2mfaN8FNJ
R0WYyaUb5jI7VN0aZzlaI0YoF5fuTeUny6wYZMzF1BV9P4GiuYaOqRd5sakmCJdy
UDxKp8w+JdmypK/gN662R0xnFylF46CRMf856NiE185nNPXEVL57kvAtg7yflRiR
3GnKXiTYVrbMcCd8IElFXNr9y1eu3WHQ0ZDLVwBl7jnzptCToYTNByGw+F0cG8vs
jZHgNY7UDgsbFes5hVorF/MhsddutlUtShrenkVji8J1aFvPgEPvViwB+lnk5pwo
7ToYJq7JX9LUgw6A18OeKh3jFoO0gfbe2rwmLFs1hYbKSJUR4r06izhTaSs8ZMf8
zHjz+zOo6n6Daq0Iegx37b0whqK4sbYvhSycBszSxPLNIHNAjvVhB0HhN3CKAsRy
IaqvsqdnsU4/wDazi+qeeand0o16VzmEgCzattupuF297p8pPZpjcp+wxI90u+lX
Okn/Gm6vaAAMTqHZivMeBXkpfLXp82r0acndZk524Xpdb0CEEomKQ/LA+TjWpRKk
pOKkiQL1G2H1fIoY20FJz8cZ/amRK4WMuz+Fkc7FqB1fyk82E6XHbqOuVHlWRS9y
GqoaedxCNnHXsKg+Z3QwtKnU6zr+MNFlLDRDzSmnpMp4pwyRPLvQzAH6tUF7fx6w
v/xyZGkWg3xfaTrVjShS21QkL6itUSzzwisXkRv/W1mErkuZtI/M4OeKvnu3S5ZX
VkSAwQ1h6mBF+FOQvUswiao5WBBST7XXl4A0xrGpIOmAnv0FZXzjFKkAl1T2YpHx
043BsJXVL/7Yjna3GzGR45AWG3iPXXet7oyk2amMUMcMxQiTl4mP35syPjbhcI/s
Hykb5KIuMv6Fp0ZkW1TKQEGf9AfaO46vKsoT0lb7nT/0pJA+6hjPnp7S4KBwgTp5
HWHZMh3qFoyKeR9n1brmzH4OqhKjgzTsohon8FkfFwOlPZeszdzhYeqx66sX4XBD
QtNa8S5bl6rcGBJ0wnzYH9RaPatAOjTsl9HlevehPfNGLPMLUa+vOXCIUJ1DxEo+
bj/B0KByLEDlqR7E9Oob5JBKBFVYpf87zQj3J5BRsMOWqgbvgREzMSB5vuhnbnx2
fYT7B29eT3XiuJmRWSqL8A4Kf6r/RgDz8co/UdoPmQiWUvbFfhE9O7DsScwMv5qS
o3tr+/6iXQ9p4gVCEkJ6XbMblQ5u5/8OkErZH2sOrL0PsGtRP1F38RHEZDUusvWs
FHet7ddGamvLEtAf9hBexQV6w3IPG40bb1vpW3OkbJYbXKzVOhgG/tuQZwIEJyS4
J/rOp72iGCb0Uu5W1lpSeIE5uzW0JxtbgfNKQHYUiVuBVVKdyVLqB3ygUscc5Yto
e8b5AX2oHihYMde77CdJL6OJ3Vtyo46w4Y7XqvsxEMGw6fu8KiBPY0fgbAc0gBYt
y/E9cL3zP7jhanX+yRnkn40uax4ABJ3T2o4zOQK8Yz93fIYL2rnfgdTwpkCsa7uZ
urVSUjfMMCAnZNqQY9Rb80yAcPcb+fIVuQybFmWut1jiYnsHVsC8w86u4BwXKsgX
7Eb+ZUdJpYn+zbT2U59hx0NeazK97MjbrMUzmT9m58tF7TslrtfwJCAHtkoHXUAG
qalbZbRViYOm/Mm4MzfEPxg4NpgZGL31WG1Z7uAW7CnbsxzB04ZodCPvVGmdNOju
T8lnx93QiIeSfV7qdQyJZxz11sRw6+v70Sa3p7+s3uw8xQ0Hik8jCVHU8hfRY/eA
S/fB8EoJUrpzpBitWmT0GjD/geRnAYzkYqzL+krYoRGJkZcO+HfQ9ASUZN9iwiEd
GDEsvsgLNU+3Z44gH6VGOvQ/hXSyqXodJacEjTSEYTVcHzfFctubT/Ox4rRyncSL
qFR3EB58j3pMBL19Qtlh3AraywiZKon0pVPmqW5shhgTMs9mwgXSO2pj8Pua1TH/
MEwZ9szhItFkVXH52IpaP+mvHtQEeO9lQyg94o4aA0Y3LzTDPVEa4jaS13m2YYcf
CsTt8REELcDZzH1ffw+wM0XywCuT3eZkbV4ISgnJ8M/6BJr/uZH3nZ4PXzUHBsdx
rS/HfKt4IPQYIJio2ag2Y346fjSycHoG2pnF4/yzk0D7hsVPgt6wc4pYKpKU6Y6v
LxjKHReMvIQznqhdbi1d8Hd6w2lnBzGH1HN6hzGO3tvkV67+kAZ3BXTWNQIUdCNL
vLd8sN41MIbd6geLksyEkWtuiFjEJDmVCX5KPNpK0P1nLh1CnKNcCe/o+KWwFPpk
0g9xqx2ay+j60ziCNC6vpBJDLttCKt0ChIrUri9g19wwdWJwRRdXhtcErxL98yAo
0Xadbxj6QW90qfjtUkxEcZTDnsi5t/QePzGuaXav6sYTsWDIGmdHwg2xdkZdacAX
i8eZFc8njxfyhftbjSBGF8GZtOOlEQ+K28jqhKORpUlFxaYBoUIreY542k4xZMli
DetxvYQnqzIoswtRml8QzY77N9IgElqLeCaU3lYwdQdqofEl5Wu4DPHQukTn21pX
nXTGHtPJk/sF2J+urXu8q1Cezi32vdmELeqEErLEpYIbEqFwPjRWtsT2naY1UjSc
1FxO5XlRwj7/Nb1tOe4DKrKy5hMZbFedzbQbs7e6S6P9xsnzd8HLj3JltTk11hky
2aE4T4Hi/l7vjaCY/B9R4iq4Gtgp9PhBljX4fKyFmbG8y2PkNsBTOo1fTTRt856n
Ev9C3mdIbdfI2N+YvesWFZ2bjIoKBTwZdaI2wTvqFZQoxQ4AY2jHbznl1yu4OCI2
MuZjpP4VZ0oL5KqVjBowQJqAJYZIvrpBTwQ9y1EHyJlCFVNU88nCph7h3wdsCiaF
JWSQMJuqhCoOgvxIGqYv15lfmB0uKYuYLO3pEEJzZAxFFmffCSvse+9yRc2HrDXE
T+GDgaivB6D+gpAfeMz+yO/64bEywATzDBAB9dCanlUE4os9KTdKZyASIjcB7+LC
eHNZPJXl0ElNQIL6BDZF7SKXwPUq6Mb7Bg+HhpvZujwcB3AvDigwSltEfoSu25hs
jbZ4GMh83Nzqr+/pTc9QG2erRFD55m6UbJVzW8j5OFRPN7faqA/yOkTitKJf/8OU
UlbXdG2FXfBugLDn6hSjiBKs2JscS/OJir67RmVP/Y7X34fYLQsMc00Kmskg7ZuF
J94YTn6bjRH8gg0dXJxRNaU7r9FFeAYLmXN+pgIpgy89sdLEDs8OjbCK2IzRH8PC
O4fhe3zAmZtUaqNvAj4ipFRLk0xznYDs1DuzjeOUYS6lJbPErndZWUdzxaPv3Bmj
eKBE+MSQmzpLMrly8eqUPQZa6bSuS2rsT5n+zy6LfvvjnXW/bG9ue7sM6r757szg
0MvK4wj8jHVPckAx9P36FSkr22GcNWlRJvSf2IMLnQ2wf5/CfZCJfC1FOAE7k9VF
6SRiJPUb1kRDG+GNi4bUpgigr0SJkuiWPWjJLRtTRSJu4dwrNCLjfMBGnqEjfJJM
TxGRG0sKS5yKnUQCG7eZmme4/65DMGlfr3XRkIOmS7xuAAgmDfw9jHZSE/Ug6tsq
k3+60e/9Y7HezrLul00k7H9LzlBRTZyv+UgTnjGgf5rvlghkq+6q9eDlhgqcA9nm
qz2P8EdHKtSbYVd67u1T3NBjerNGHjqnCEgp1Q5HjS7v17b7DnhPVgWyNsys+O88
eSNhc0aGjvYheKGadz59Mu7oFDCjN8OVhR2ZKCwR/DLUCKAfhhHL+x98TL7u5lxs
+a/sHtQ+scnEHFucW3GzRe3ZkLGbePXSfzbmyrhInA+HNKCxje3mW1Ci+lcQPxW7
4LqmCOlCZmgDFn0k7YHF7FkLuKuR7NOY8a8LIWI97BgJql5CmtiBr4WGctM7mXZW
deX0iWFZomoEsHtaDaefSacxkj/dV2grxLXoTFEE+7HWDrWnTFvrUUkhcfxVOgAW
JPNN/MCR8JXOCK2kJXlfkdssFkOPL65ALQqRvWyAACPURfIZPhqkHnaVYM2UYhFT
wzYcnoVi2EOj+0ERdwfXxJ2nVkrSdTZSi/KgDbD56vQlKFIOuTJP7Mjww2ZyS7Bc
Kc88F+otFJCHvO92lnZEEziU6j2XZeHCj5gTYCPZL1t4TThDc6y+97va964zs4gu
kL2LSGV7DiuLtydTkNHMbw73rCETAOUeVU2Z55TvKEmHJEETpIr0IPmBtreiv5pH
gNVsVnkeDZKOupN2tvbrY/s3NjTie+U979e3AQ3Svr9ERyYZUO6UQKud0Y40KI2v
m8Zuby7JDAc/7zlkMyR7Vg+t/zp7vXJVm0JIQwtpsFilMA/RYXZWzCKc41GrPsBK
2YMuUbpL4PcjsWw2Cez9eFaTNGCeHynLilpzgfrNAO9gNvVM90+um8H7+IeEi4Ac
S4mERkn+d1TtvUR5xCxzu0oricYoIt5g+wjYpXj9ehZu6P6GXlxiX6JrCnG7BozZ
bWrxYQk+LfhGJf+Z7eBwz6L/6u1GwmmFCb/D7stERd7SjUo0XFbwi5x6uM/HGNhc
V+B9tsPJ9LxZTbKjf/d2Rv7TIpAA3jUZQ3GGGspPOZE3ZEwWziZzZtZt2+ys6CVG
XReesDqa6sG4+5pMlL81uDDTB0l9G2/HiQtKPtCJmSHvq60lfSHUvtWlmUgB7H4g
dkIXMRZ1lO+fxsc2W55sD0uoW/E5AFVYGdvgEIWIz0oJcSEoneLtaWDx1m+ylHnk
0VVy8ECv6FVK2fGDVVZDn6hMEetjlnBll9tjJmcHwUIqQMMtgCtLj/1Q4/gzWRil
nTnXwP0w1TRDpFxxDOOGERBXgjbp0kkE/hrMV4OOm1BmJ9c1LThHDFPFGVf9wrdv
gpiHtuejL5ylIzBVl3Fy7DMVnczoN+jrq+dC4PudLhNukcKJg291S/3blQAxm7Ib
fkIQoJIKu1TYL5UoBNK/oHZIuMOfQI/eXpUhQL/UDM16z8j2r2ZiaaBC8KbTEUnH
SIw/nJ2gp9w9Cc6liQ+CPV0Fsht9Lfe0RpkQEeZfPPg59Ax94BsadEwY9r0tREru
78JrfG1iq2z9X/xsZXhv1F0LEAgr7P0ziMqPhsd1RhHyLj4Bh7GI+7YYQp3pghA/
dmr1wJsFDEZlebicbVM4fRodg+IX3BaIrU+BoHQsL81nSECdWP6eS+7UAibi6VLY
QCw0id9FiBYxXvI3TDM4utPUtsA2s/X6I4haeIm9cYJLAG+gr5yWeTe8plUTXb5w
7+rfueoAu2nJhAAfUfLGmcgXYoL7v91ex8jO/2CWXZ6t17nM2Jl4J8qRzgLdWdaA
yKIdinPg/Rg4Dv9G5grVyutauiT2/VH0eNNrrEuh4OpXGMr1ytSc09AYixWqySig
huoKSyDGoFX7yoHW9GcGF+LP/qL5hwvnJz9XfOa4+wf/BEXuUZMIDUTDqeivKPGq
TXsazST94MUHqSBzFkG/H4EL7rMXBS1CyQec3QnOa0ZK6DkvWT1WFlMZ5CQn07dy
lfboyyvtoQTGOBLIZJAG6tXODoOyn5OoKE5QPT57933Yvopdqoofu2H3Jf0HCEau
8U8lZV8rlMkH9Q86Qr0iBFcUY7I4LiveNbHFlMOyX0wuzhRtIkWvypxH9R8E3N/r
Gq0l1iZZ+q7tbHcAIsCtjyazXnqzMA4pfhp4V9H7NdzQlne2ET/NFsjBNmGTX2SQ
1q8NJWzdTtwblkqsMFMMGfoffLmK5pVuCULOT0BRif3S/j5RW6r6suxSqYEVktRC
cHIo/tbnhz9OJGlumPPmwjdtpBJcqvSZ3/YXIr7DyyWvIw0CipTQfEa5/J8SDtll
0OuwAYklKRDmn+aHYqT2IOrx5gdNyyTmX+5YlxZkAcrOy5iJZtZm/OkfP4X74Akh
tv4aNPrLyKxm5mF1CWmJeDlQQKWnG257Wg87RUMZJG0fZwyAAQ4j1RrHx2uG7dDy
KJKbKcfATy0DfmBNX8g/lpbwxu0P+6DGv+YQZm/mOx74Q6AijihGWzrfqsoe1juu
PFrNla+1jZBi1ZVNdm1QozA6biTFKmYITrPBMunSGzELjD7qHCm9RForb4AXVxtB
qeIzuGfdSGz1kOql84Y+0Q7RoFgK+rt4ZPGG0O/ylcHK/T/XOOKQgQ9Od6RE8gex
qtqA/IbNmX+7aKE0FMzXvGbCrtblNb/ZNmwKJBTGxP6HhetLfJA6tI2Okgv8FATP
bl+4rzxqAEQmdhkCVm2z8lXCO+t6Rlt0mGWTbMXTvtVYsjbKFi4AbJRryHSufyuv
97gaGecWP41cky6tzXHzSXCqKZ5Le8gOAnja+AnNf7o4ukJsROdHH6COT06jj4Bp
HzMH3jGNtdX8XGL8Z1j/1W5FtpGKLy/MCy52SIkVGcaYxQbq13SG+hlzQ8DyvMry
Sq7RFGPxIc01YSJkoKwANfpKZG1IqriJ7VH2XJ2JqgFvx0kaLjtlYl24W9gifvKW
XpCV7vqR6L8N8R2t1ve06Gds426EZ6A59zY8Y39TmeVsJfcDkSCamANwGIuEPEsX
Sz7pRptRhz7qT7oUE3lzTWodRTTl4iz2dZT2Lc6bwh7gusZQ8kMfmVL/jbrityWa
Qd2E5jZGrGkPr3JqK05zxebx0ozOnPTYyYfNcJ+ieugZQRMNgEn9WX/RIqTixQkR
0SUoKqs4QEMRMAL/IDiMwOoGVt5PoGJUkN0aaReAQd6gQOGMsXBYqd6hystnpaB2
bsUi/nSwMYYgNFMRDwjcrmjp8fkcAoIBWnI0qB3Ygdnxb6zSYYWnMhkwBtzmdb/9
fnR1yDOf6VHxF7dS61Z6HPOKYQ0KFBvnERrTAzPUXoon7DB9yZXAUDxboIj7ZDob
sPcEKOAowCEoIlB5SNA2qgVDABRsqLWP+GZYdwfcIELJ9i/fGSdeeohbAcbE5p08
PNIwtQLTXRdyHw+0Yl7X3tiuN9R/JM1KK2FbA5qOvlWDZHO8FXP/Spc9h7d4E4A9
stKeToV22NgekT18JO1bCW3+Ho3NkSp/heLEzaoLcYs3vI719bQIyA+MfvXpK+Mf
YhLw9Jkt+5rng8/quGR6HR0rm5MnwdP/vvFdTeofAAgITjU0rT3j46+AtJJSioKN
BNlK5Rx2cJ7HOmbe7sLQg7DRgXCAlQysLS/6/AycBiYgY0UyYoyytBVkFR8RvvTX
+AYW2F1OtvtAHEF4Cqf5FkdfbtNs0Bl1fv78LNNbf3or4lA9JhWNdHtNQkNppt9o
XTeauwyEKDqvqkkXYKQXiqofkCsVyHxHb5lhGEKvCThIxfLry5nWz0qmLr7ZPs8Q
Qo71D4l1nNAx0QPTDnno0xEshc68nkw3DlTp6l53YJCAoEduMOcu5dpymItpJIz9
bCy9x4rSE5i1L5++LMhnM5MJf1Zy9361u2lDTJGbcfKabVRi0fGyueNYEdMBuolK
SSfpyYu3qElj3kuWrx9tuTziFSubflQ7BAGSCIYkiG5l8WxSMJFPEGEXo05GLOdN
obgWELFeJJ3A3YZMMSCr/zF+bdCgu5Z6dNUPvBHUiOuJvCLEwJ+bATfVvoImUw9a
BstuzJcFUoCUUmTURl7i6Py6rQ9pnV9ZLGE/adAfbT1x8bUZWXsdnza+ACYj3qBp
+t4luRWs3psyoywcEpvpmqUprtRJ5vXSsxC9/W3+QjJMal4+qEZSYGs/RSLuI9IL
zm5kftM0Qt3MXOEbeHFFmv0UKhrRyb9ypeVW+1yS1S5MhIP3rj+UYI4NznI8uKNm
EeDgtoCRkqGEqeQ1WjnO2tNCuh7spLFkmQX78gzxAA1vmGNc1GsTo2dUmpdwFYX2
GrlUsPvGDbIMMZB85szXJopoWSXJWjXBfuG1T436xUg5ugvq4j3HJ+4s1TbtxOGe
f9jHhnetnrFzhI84k9aswQ895O77x+JvedJYmkkMYrzCBEj7j7uaw/3szfL+aRoi
Kp3Lshrd6Y9F2N9T6eFPWjixhHk8KADab+zjfbCNs0GH7OHIKpXCVKr9PdILA6M0
lErvKAsc3odEM9UzaWs86pKxgr0qrjQyc29LcQSBIxIMFUtsh8nhCZ//m3XZdo5l
7ga4OndFa51ExyA+yk4YLFbaJxbz048tncXi+3CrvHpTHDT4o6W0PxX3Mo474Cow
hiygCEXB6V5yRTQAS7LHS0hxjLfQX63r8fpst2RwsNvhms/sbLF1rr4v45JJMP6W
DXXN0E/VjyoGX3Az3l53bUmySqcpLFoK7SplEMHAhbMLH2yFePwWX+IDlfvApXZd
zsny+Vs758ZyTrptTeSj+9FKJ8vuQNLdZpnlAEWyjpHx7ob40hx9uBJPayJ9Og0s
SAL3uhhN2PIvqKMXzLRB5JpJMzmh0I1PV1qGjMupoCpksZ61hXccJDhWjbrAcgbO
CU7VTPFnoEMtdX027wL3h8fioSH6E6Rmi9doSVfPM97uSwbzTvvOJ00nZjkV7W2I
8xc4PmWa1cNwJo0IYXFzkn5SJX6HlCD+3fpmPrueQe//r1WD7BYj2A9cMGOXstYi
1012nNmDWhsxgc+lT1agnCxGstOI4MjRotN247MEMcrHTzJWk0dW/F/acbuyPS/U
nt+zNqFq71hJPEYQDT+X3w+sh+Ex52BKoLbVF6g8cuKTqHPKNYOAmDMkSunn7PUS
kSVIvXY8I/NXExaB4P4k+rbmgdDleTdt9th9s3dMjOR9UUJYgBk6jHd87k3bwvoq
ToShp/Hdlc39Xip00myj/8s5yByxiHKEFNwJsaNODHNYZp9Fo6JvqgpuuT7amaIJ
STyPfMX5tCe32RNsfMZEkYxEsuW/8YglBID8R4r5qUraYoWfw2/UPwVw+UBeNjh0
cADhL7RqAo6KMZvH9LheRtv1RmgSj0I5b8+cKMbfh+2HMRiIscRfGRxbN3GeKN3Q
TF8r2GBjzqQh95u8ON34gH6da/Uu1WeryzlHo0sLDcfibX4K2GbJwHz658KWvtdA
9kghLENfbtZ1Kiz1dB6UyvNkxJHv6hX9tGAsi8CRKJBBCL94cnwwA/14yzTBEKfb
sDs3EwYFpeyuW2KauFI4Vua1i+GKrR9L/u4Tr017uKSlTE0ySCjUmo0yFs8FFYVj
HqcoP3p/Yd9MsQdUPD1hfmq1Rd+N4t1uBkVn4kjVfBMP48u7Fj9wfll3ZX0uO11l
et8yb4ooOELMF3WrMA4aKY/DhulpwoJwNEen+9dEC2cPELyl+LfskvTV2mlJ4yw2
AC3tjw+JYZyTDJ+s+1EpW5V28YZM8+UgsiZfdfdtZ/IrkGpr6iMVN2MXq2DQs4Um
7oFxk4G4wIcw/H1+Qk53f5rap/owKi3odc+kspEkjbu70Vm3keR4DbdP3NSgvVyA
dyYZkhg7+JhDcJMumwuPjHqjgrFe77ZBzeJCXgkZjvbDX6v1hiAEjaslOTUwxC0n
RjAW6QXdPOLBYxpNq3aPLo47IIAChLNTUw7NtLVotxXgG24zcNEreMU9oDO5S9X3
TKhY7GXfeGxwl9R4LKnpctPVdG7W5QXxrxQ3Hjl03wgmJzZSsK5fxreC9d7BGzEF
Gsq06zgRckX3poSi1o2pzjNzBL5SjdyhHQZ1NA9/JXMoxivwKCwdj9qj2xwlWcU2
BySkvEzY9jLUs7b7jcdGsZKMOVg5Jq2VEGyLtu1PvzlJ4sqAJo7imGO7YgKJUblD
UJthIcYB7BfWak6F1Knd3Apw1P9FfmWYmG/6xuAgvXqvi2R6ekspkTarNjPvwdlI
Qh/Wa6KKOnpaoztKzDZsgADFOXQdLc3cgFF39MNGo2DV0TJm7PlbuhDvzHg3xnwL
vobjtREaUUvo3jv6x42did8oY5Bt5ihuqhGYsninPSvSCEE23hoS8sXiLEJVCtwH
EuG9SOT+5K4+Z3wwQmk6ShcKa0t0a1Nvm0MyTY0ze4YAEEwpob2niBooMl0Lzw/+
R/HPfJhczTgBESdhRpy6M7GHcdcwd1n4B7WH2tk57fzt1mZRhWxsc4xZxMcne+yc
/ZMmr/jilu80hTcCH/qraBfno9NITQTbuLcqcYREfYj/ExXsAcdpyyR+cQEeRBHR
tV1g/q6xgIlY+kqolnEZvpAF3IeWaI2QoN7I9M5RfaFt9pq62b+8jH6zdlAbwEhX
jrc+FpTMvB2vOg0o24fwPA7O7zXndWQ2pshgeYVe9KNDCpMa4048L8xMX4Gs8yW+
rjOqkKQruJotLEplGKqx1Z1Y7++M4SmJZn5vE3yhZR7Zn9v5PBnSbMUejrCoiiJh
GuUALQwvpAcQ2NtE688nkHh0pUxrfKzj7XoQ0QL9RT77u4jKtGH1jt29uogmnohD
UbQSq6CrmJk9C0kyQdA4Mad8/jeQ3tyL+L99xppLK3sFTyaNYTjnmBuKXkpFpxIa
YuiOCe7qtdY05D5UWCjpKWTBTUsaWjv+U0Ae3AQPviwKInTK534cM/xm3aViJUhL
Kq2JM0kLlyE0oxXZZgtn5dwYtlwP4V4A/y2o74K/RlXPKmlvxrXtOcGEapOczzdr
ipEyMZK+NLwcKwym3bG2IoLrh/ImDm7Ot8hwhQ8iM+MU7yFI7cUO3J8Dw/WFFjMJ
Ilubcy94gDr7Ek47o5/xEopdCMd0+R7Bl0yjUEIg++eVaIbAJFiWbALrKFammZ55
43U/qj9hnTceqVWkMngGffjFEGUdMegZY79Z8Gye6raa7DPnIsWlBcbFCFYk53y1
ht01t5iU1PHg+H+UNn87VyfoRIa+vwhr0wy4GCcuBz0r2nog6e/qoWNVpUS6STUs
I2qFDQWXq4YUKK07mBDKsAZbnJmVv9Rv/6RK9zHMlyulA3MApLKghsk/d9D1v/Oj
1Y31AxWBNSkS1nSkiK4nEhKemaUT7AnUX6bGbUdGUhY1BZIiRQWWqaJqSWmtXaMJ
lTnGkkJ4il7OTYIpQDIasah/sg9191pA16tn8GBoV+ck9YK/zSA7aXIR2Hm5Ngt4
DPvvs//Jrx3q/95CzEF2JuE1GtsWobNk7Mie2EFja4UANs2SLjMuQUTJSpSSQF2L
wKihbpbDBYnCS87m8A7C3u6N1Q7L5E0h6KfpNFwuM9Kj4kk6pe1Lt4lIvEOlIgZV
XFAfxkObb5TE6QHqHuR+Mj0UozQN5YY2QY8t1kVYLcoKP+5KL3XCJl8cLJ0dKGat
HavoOumgHLTvlvP+Gek1djM1qw4Ahzcq4fY0e03yXbmIrsFPFKdoyXDjw7EKooIU
qJXTlI1IVvv0R+WvRAvPP3umH6UKcZcDJOz7rZLhD4oBZKSRTgws8NjfrUIcF+pm
oOX0pH6gbR+iPtapigmK+ArFqdDN5Spe722/H4T2nvPQzsO8MZe82NyTl7tAysPx
1FomdRe0aT3IeQp2n2EXlgpdoLRudFreZ5Z+bmiIMlPZe3UwmeiEoK1i7oM0BNky
juBvlqbSxzh/e3Ic+NJZsJtkWiTC1qnQUjzrJxs5jXMwKcmZ88tPF/GI2ZYdcNN+
yoblWeISpcTaHnJr5xwB+lmNNCzs5GxwMLmciqdBfdwX1LihackRAli0/CU1gcmt
A1fNR/ij975eGFBmLD1vXM3/tF1Ve+CawtM/HR+TolRwB2AvPayoJdz7uZj74tcA
P/issH07vjvZiC5OHuo5VZX+yuuJTvhMjE9dzthzJxipKPo40YBfjxcFXcchsk0h
xJRizqelbhX2NEZ3NExdgUUvxEoXas/rm+LhJMLV3gXscbhf2UAS+x9IVyrlDcxX
/apALzhQ/DSa4nRHEyU5f4jDT3jLdFztZPHz25r4cz+NPltNsZc27Obsjx/ACyKI
RYGfP3wS0LRCYZJNAyJqy9iDuBByM/Yo8njQKpZCbvTG7TfSnmzza1NnFqG2kmr6
BYOCU/d9K3E7IRKw6CjnM5drxpcO7uuqNF8ezSiXZ5ZG1yiT3hieLH+nuakTUU8l
fcEbF3o3ppOQfr/DV6FZ5MHZugUKZ1a7mvwxm19iI6VDuk4NkT+Isf1VVvk+B4DN
dkZU2hxG3USch5ub8SBKRZuFmxlGRlMFuSMob1hEn2W/emQ25z0gBzEwsOoSkbXV
/gj6AayBfeyKDzAmHkK1DobXn3dl/Nqu9cl/n7AfG67onjxCdrasgxTfGfgyUSmC
MXcFDBN6eUM0eE9QXHGqaeF7g0jB6jtnftCqxmIMhzoxlQNLgudLmAdB2Q2l3fuD
eg0HrzH8NHiNDZLCK/bj+cXaY2QX+UUth3Kv29pSD5Evev8+8P5BxaQUzF3XOZJU
oW3xCOaE+sp8V5FQGbljNEnGsRUsB93DvmwyxCzIumHK4qsCKMrjZm1sSuePbP6+
k63yrXLmkTMFSfRgmj1fx6RQf0W6lzib8VEitoVQ4oSs3PLkD1HXtcBA0mdN2hyp
W1YuhpZrh9UB+GoSNtZP34zHcmI6DrZurjEezb/kJC1eZy+NxmyN37hqxcJfVAYf
oIcyQiBDZ1ce4h09MxmM+BOmVJw7GD9sF6LrwBfAlic3Rd4y2U8mJWRaiioQB6Iq
9qsOUO28xlSgl88aC1z5iW8tUUydislKE4ocpivji9+FNmw5kr7EGtWtZZnCRfrW
5x0U0iFDda76tLVaVA1fDgvE4RNsQLhqEniO+EJqUxXY9IUz9BnkGBTp1Ygyj6d1
RTmmCv/vCDmuo7sIBC9/DMXCxpxdXJ17gDTYZrmSRrbLhUKOMRsMXs0JeeLu8mft
uA6rv1RM2Lev6wCgvmR1WEG1jl3ewpo/HrSA0R9qcRZugoMlEDr0mwIiHTmcQNHR
+ga9nRQG2dYZiOMfK1IARj1uvG+4jMB6ILX1crPIWkGbohSRKYSjm/iaWZxlSZ/4
me+UbDR8KbMCOFliNdU+cl9tmnp76QtFNjDDkbDSdmMjQzBsXYb2do7+2ylOSTix
rOkI5rI+8w5j9VtpPV317JfvmyZFH5bdK0QU0CdUoTRjgNFhaQa53G+u+tQaQ5Gs
uaY/lWRKRIkB4Dp8DaeQIfMTf4tgUm+ncU7HLjPEw67ha+aWKUlyHcktF42h/RXO
z6TPJ9TYx5oQOCdBuixELEZydzYvMkXWyncLuVE8WSjdM7Knu+FtCFCxNEskZtqY
G6oXe+Wwy9VnXQVO14p88ytphZ+FrPLha7La2ImfvulX4mXU/Lzzz8c6sfq0+S8P
OROWMLfJsjyiveyTG/x657Yfi/q1ExdhqeUQ25B/zcfog40GgOnkKCKqCTBKCXJb
nRueBbUxW/sEKSGxbAbxfixirCsgjMNnXEEqcRigl9yWCiZ2VI169JgNAI/mjH76
5b2OHKHtU+eyUtQArE4iViE/teIvma4PB66k73Yfh7NofK1XdJD59HODCYvIUvie
lJ9NG91fH/0tpGkSO57SROneo9h82cmi6SKzjZ39WGAqVwyvYtFjjia4i239L8Gj
76JMJ3GVkFEARCYU0MT6VXvUnVC7E9zFe6H5cc2V4Xxlw0DxrpVnjH1uJmqBG5BN
O5TJi4se0w5K6VNlVPntvaOXcEA9Y8hC4N0k0TlkNT9mKhCukztQxNVsZCmYDihb
X45u6ZMzxjbpQgHnA71uF5gsF6NUBUp02upFkZCRlNwv+b10W0JG6VLnDis/YsQ7
l3m+BPZF3ukwV3WhEyOUq8YTPN9t3tzy42Rh7CZrnGNI/1hIMGQzUxnpyB5jgXVK
KlVHYqh7tPM/wW8CZ8dHf/CFlOvrQBuKzJaiOVx5uZAT3sXwEiB4fdFwJ5LpIVhV
PXWGd01p47XSQ0UwpZP+4wjUshXlye+uexicplIocGOwPRQvoelfvjJtB6If0J23
oHUpdvt/1Z7v3RULA5hAYyg5EFNZBvKn8EzapGmML9Zj5gCEnPqnBTyMhytwdrRu
HmxgEibNkQsfTMxIHDAVu6LzTlUDS9MdmsPwCnJfiHg8IDAfBphAC467eGQIXzqg
CJjBFHYONUJltZIDM3YepI04yZbBH72nv46JvkoSkXLtigfTMz56P1ILzekeeVl4
oUcOElQPH0yBT6rGvMb5eWOUneWXXLde35jU9IfufSbh3OViky7N/zzp0Lw09Plz
Y+nHX49YsOZG0dZpY6PDINC2WQgctc/pLB4bcdrYPXoHQjTEkpDG/hNxps5ldQis
AfqTIZRnbOV4tOdjE46P7/LWvHitsljCm/8K0YLjnWXihC12GQ0RkgrkgeWy6pDT
/Ep88T7XddIooI4+eScH8R8eNLIYMLECWpVn4cnSHZhqYBp6r0Sr9Yp76VcdmFM1
DdYYhorwKe1dDiGYvtk9h5WqrR66OoG44hY3Vm3ucfSX6r97+jFhsQIS9Of9bvH7
P6PSBQz28KyYcFyKvp77fexx7wVGRrUTSKEHByXebujsQZUOgeY6Xk67WsksCCSP
9TT1HlSX3wU+WTPkVRrBGw4Jja2z9oQ3iiuKBVOqSMMANX1mxZqk/Di7V3pR5ySY
oeXqIA8Aj1iqxadhaYTu9lkdUoqmppybvz/EDxvqYx4U0bRz0mU+mE9afmU/WJK9
BWMzvWHJrQqjCC0Xc3ostiHFbKMVIkHUZa+yXHYBBDaUPqzuNSsGZ3zxod56fZdS
2yWRyuTPcVHzU1FelEFKMJIB3ZFqkC/GSwR8mSGtM+m9XwAHM9SS+z0QwQhs2oG/
w87XBUFQ+thcK3nMzSU5zDoLZaK+ghJdCAE0sXRl740XTmLNl4sJ8rPyz6stsBUQ
aDA+Xj+qbJp8LBz0QoDZK0wEAxOeQZUDVah0xuPZbeGkahj7UmN20bb5mVSzbZUv
9Od7ctm/5TCsiQm2znpsMozwl3JCa8VojuuxlU39NdrQ9dJSG7j9tW2BmJXEiABR
IqIlE4w6viV8CHNf2I1C6g8/3BePoQz1NxRFlT5WnYCFzJm7rOG/aC7bwI9rxGk/
0MrSfqKGEYQpPNhpiK17FIlYRvjr5x+ZvvPsLSmjVGPZeqjbXmQqn+VNZH+FbX+Q
AHPClxpOrwVwQX4zuVIvPQD9en6FgHXf2rcMbTN+NwpLFNbJpy/dxBu9XpstyMA/
VJrMrTbp8A6APXGp5P7yPlMbnalE24VXU2myPMrSnbT+0gVEy8yrlSLB4BXOOQN2
xUooK3LEJOUvp/n/7W3coSZYKiJpBMu3AMiKlv87KYskDIW/0TNPIc0L/VbSzzHU
K0yHzO6p0ySbBpm/50oDTo1uTc2aUGFRgIigIXa9POeRxXU4TH/GX1hsGxkODXFo
QnzYyQy3wYbdm9QIPrg5eRonwBnCYoczwz2OxdM6Lu3BZL0Epqk8cXi499CCtXfP
JtciiDxyyObGdgFgMdYOSlKS920Em1hgxj1nzdyckTsqORKHvBseMY0iAKHKiwQk
i3FeFRtpzBxNZQRWvKHvHR6Tj6DXK32YflvkMhzVWRh3YGhEFDt0/EVcI6XJdYmy
7/nbsoIqb8kNZWoIX3F/DHvK+Iij9kpRZloEtYyGizUARUK5v7rVpPbJyERL3U3a
5HzvVYKp9sf8roWfYreKimv9gT33NKNKK8XeX3/NwP8eLdqrtLQHOv0jSPwaPgtY
b1E3Fdjw27Dn8UWDfpodnUOC2qfKEH3D+nbTI3c6EnbmfpZEz7Nk+zU+Z459ptew
zLTes3lFgHMC4glKdEdOGonUyBfTYWr1xVRbEpc7hoNFHgokzt9fQCwXoW13CPn5
5AX9y12yxuumMj1epxpQ3uFdrZ5tYXqkcveBn5CdZJ2rqmlsaTaYK4kgGWpDeK4X
4/fM67WxpS3Uv2/vFF/Fqx8FZDhw5Qougo6xvwoJDwLrWxXqxjN/ftrsV807D+mJ
8kUhz+Z8BwIE9t7oeZugpVTjeekggIwVaQ3e+xYOSEbckNaJ7RELEt/U5M6fIbl0
4Tr6nyYBr8msvLcGFf/Xvi/YCh1iYa2+D3z0A4Dj2VTaFAAfSx/ryAhXGU1zX52N
FesqaBsTF2PQdleJqHTbCG0bYT4T4RLpMvhB1CNqEAfvdbt9Mn4BE/lDfL1NW89t
uy2C2O7JjXzR0mQ6MIhvVyOzowE3D9gWk/6HsOL2wAJl20ckbf5um4ZrNX+zzLbd
/t1nHUE2unmYNhS5UNH51/QkD0kjZjadVaSwz3bZ4kgmPvZP2Ta147Xg+KKRf+jt
s26gsJb9+3EudWme78xTz+XaJ6acwkRw7HJJmUzDkTIDF6ZYUfWCjUaI+Pw41Amp
qvQVinVE25UWOHD6dE1wnYcrtc1o9r3vv++WepC/fc+EhCR2DuUwJpVw1SL+wQRi
Z0C8wcvE86R1djhNf/TVDLOf5WmBlkrkRUhVHquY0IROTkHvX0WfXtsYIfPaygkE
EZnDHXtE15r0TWrmLRtziYU3cYA3FLFUOh4pw5cQi5eR0MQfESO4Ew4GrIo8MROq
dTpGWc7XMu6a2nHp4mnjWPqHGgg6xHKkmvElTaqEddNpDUrPHGPTL+PoNcgxwZFT
iDjIt+ITBjbMYKnMxvjsEpDYp/+7UXKD0fFKssrDeLtC8AvAPTz7ps2L7twkdzLd
jRe9VcByNtAy2dg+e0p6WUsO/BiUd/2cl1AlN6J01/JRSyfW7B8TdelO+Z/GJAdM
Fv1M341yjbACGTgbx578KXJ2j23ciAoOZRvq5XYUzrgdbuQmD7xJpsn7Eex17oBl
HD0lNv9ONAwzzS8/Wwp3y/OBE+Rd9G4V66PTwoVkxBdc/DRRNKPF+e6/DRrkRm+2
ePywozEqq05SpRNS2MbMKTwUtYWArWbP02GxdLS1Uzwy+IVlKVwNCRXtvrp0Pvld
YtT/ha4o6YZY9x0WNczyPFU4YaGnaO3QdO88BnBICOyfEMy5ftoLObfNfqKlCtZ7
Fx726ZmBMbgVZaR8T4uqjMtnoQPnkFaAZmsIgMt9NmSW39j//l3FyJPepStVcRUe
fD/eFxAVEWMO4wUkdSh5XlrHA9+9Tylfn94dHPjja/ds5OR4FUS+Yen3XzLCxT7a
18rvSqNxkywqI+NeeYwO3qFiN2hoVK4ukw0EnCMWr7KLGXHQiDCmxDCiiFHL0IlG
3WOz/R5hyf80MivJe1Txv7jlzKsmbLtcQ5xylQfY33ZZv0AlRb01SL4rZNMo8NQO
D3UM6TrkyF4e4EplTVR5Hc2fomvLj/39M3riW6CuunAGKWlFbpGKYbUysgkUr20n
v/UB/ss4KhQa0WjAM8XSfLd9edcQxrYteEPVxfmUDyS1rcPUp2Jqc4H8Z9rKKoW5
3OjUL66Intwm6KH03YQH5hEjzIv7JsfzSmfQWVhSK11vgDFIO6eMK+DizA5RsHff
p7oNdMntYXG0txLzJWWogkvOob9DCmPtY7ZPVf+27yPPITwrsjsRaFA8RWUrfIXu
vqAvbUNZC0+AZf2k5pBmRwvULXP6kvnOPuA6/92eFKrjujixRtCd3m7/DYcRYpPn
t8afTA3vG7sLmXInJSl5BQOZJy2NowFeZbwvdr+PDjvr1LQnUrwg9SZ6AjvyJIfn
C4PnTyn7lM05WcAVQafUlOI73Owe5zQKzO5J+9qO+deq+TOTCOGr7NcG4RaYvwFq
Gw2q5S00d581uE74qQHFllxCPfXeGgcE3nHkxoxEMKOdh8e6/MtreCeO0JSlqeXH
Xo3Fr5IgrNJwPELTXJyVZJ3ZrZTvORGuM6Azns+lVn1sAJK1wHRQhijGTY+AZv0p
POMnahVFzC8E+DgjOHD8DjIgsyeShMqcCWBsb8ZAsPBr1nAqOmELyo7DXfQMigni
wEVREzDmsl48gbhanekEy/6Qeto2Hbll/oZcHIkdRLk4XYWBf2kQcOgindn+i5bF
e+YC+ZOp9Xid+lwj88TqaduFOBaWFkGQNTb+egLmml71ezfCm7YZcL/wMrpsC+un
Fmo9ju15DgwKCPnLiBQpX/+NBnw/CU6u8pUSjeqlQ9d6V7XOSjrvSfbMNxRPb4tk
mTeRo8PpIGzdf/n465/TNPM//CmFwpDJMHEqO9IlY4r1x4rR0444wCiQBiJqP/+u
nhKQW1Te0aGBVNjs20lKKsW8D4Kdg6y13SvzSZPBNcuclBj7Vgtv0qVw2J4LbiqP
vFP3uhY1K2/+f9GvV2OnkK9Uh1Lrkx6jR4SI5FbZBfADHstf/YFN8Dc92k1HHX1O
kJzprvqbEscxb9zcpzDZYNbF1+imwPQ0TBfxzDvF0Q6YpjAK+i6DONr68SzOo3tb
YyRAj240X9iug/b6UffCgHo7ZI7wFrNs5e8zT6yYo+3IWoQ0+LPjWyQr1hUXji6f
T1bblE+BsDxqFCI8Nv0a7i1av+cBCkRXJe8OplezsPZboFhW21oPE6mQYl/zpwNV
myyCVozatNdtBI2U0JhhBnUnskta8pj2G5znjsOpX9J8sYay5eSx33KOFsgTexVk
f9zy5VhCRdirXHIXNwPDG12kcDC+ORlsIG4AZI52JlCfHAyHwnTp3lVt4GamHymQ
HdnUTvzzIEvoAcwiM8i72r+9/rban/l9Yo3va3/eVvG66KzR0NuEjhYPKmplobjq
r7arJqEfKPWuXjOs8LI4CHVD/UBHkv8s+qJcnnpFSaEGNSZTcm+zQXNTo0KaK/T4
cMhntb/A6+7IWLLWqNFDjjKgkSoM0zFqUOLTO5OG/7rQu97MqnugWSz9P2334gw+
oA/g1eqYdGfh/fgrkumuTxQmMkdaCkCBoQcuHbGSsmcoOg9FRToh+A/RpiQEMUa/
jM2ms11Ce1ePlhAzQZqIVp9QSk5E4UF4Th1KqZY+c2tc9fCaKJRQtnPzjUYekDjt
OtX6xuBmkvyt5pQGHJPCaJrv+VXI987HyzcTInUa4JU6AS5PJc1UPwK3U1jXBQ+r
O267l27QfJB31a/HQQCjoasvOb0XDxVSQjXFSuxv+yIHj3x8KS/QXWwmao3mQNvk
v0lzyXaPGYeN7XcIOmwJ3Nl9n+pFLi0y/yfywGkf+uokm/lAMiasLHfewTsym5gS
SeU/LQqaQ9gqM9pcLPVSQl0rHjAPKNzXZ2Pta2FufTvj2SBrfTZvqRyG3gHXKFwl
g4ysA6OhEd+tK7wYqdfaq1sNCZqZZS1HpoXCOzJdhZeJHB/xpDlIfQeU3G6W9tZx
vFNob5LcISbfYF0BEvqlpjEkKX7zAYDd8L+Uoxbxfpm5abhvitxiQC9+O59raNN+
YT8DMtrKBUrYgePmIGT0PHafwW3Za94Y+HG8TseYKavXOhHQK3ECllqc+5pWgwrH
G0ljCHCHdmVfQ1QQeFX3ZxH3ibkWEifJApzKLRdE6sKd9JOUGVVwFJTrFqX1MoPR
Y7iWl0IZT8JgekiX36Md6tKG8nrvLFwRcljRq7e3G7Zdyv7lSRdyHNl0HGom1LxQ
ac6v8wgmDL0qg2onJw+o4R/G/zCXO8KIDKfdnqMJ9UaFaFyFvsMI6TtPLuJTANNB
cGhahmJerOlHrDObOyDin6Fw6pcDamvlSFVrvTf4JQttB1+xSER+/RoxW45a1Pzb
WkuN01YUsQ6rs0/YzdVcBFfSN4u5DyuJc3kqZc97Ww2Vvi2PjAobPlRR5UNxBhTx
HDEdSGR70UfPvuWm2eyDw8wALhzdQYgyaE77fxdlIJ25Akg8zhENIk3wXgJRwAGq
JhmPbY14e17nSOGY7Ps9s568qi3K+9EGfyrX0y8ic5yFVvu18HqlPGGdoTu0TN37
jQrkTlFln7HkmJ1T7MejEDFRdtSOb4B0UR/ZQpaVQlEJ+dyK/47JQAiDoBauPj2w
68qNVTUrLTdGlMHg9rn9eqF9qmSCKq/u6YbH/kHZvuHxga0WRkvA0RALdXTegcwy
YVm7gLPQCY/5SGxcHA6uBt0LUTkP6Q2CchLGVN7CAPpB/peTet/8x0dQChUH80Kq
7Cc/WiBl2tg41NXUH/2vf4yRvgcdGQLAvHMwLt1IpTqdmJC7k7Q526xxJOY1fw3k
aUtCJIzqapRbzI6YGmc2HXq0jUIgK3HiO4mrcZRAOSOA+bDZaWN6NugKLnpNjxRy
ePbxNkjobSNCxoHPrgwO79t194YyZC8SOjUcnM2EwpArX/Re4Em66J0QAF1NsNb3
1kE6tCXjdem5J0Dc18EUGP9rnSobHVghAkIAGLwpcrB7dGSS2emZJ4klJkR1SFMq
r0u+wodrzRVkRDU1IwlCVO8l5ZRPHc+5vKKoALBpiQh9fkXYCbOnMwL30qxBmZZu
t9DK3K4xoENL2LVuULlMUK8tu8MOhLhMUl6H7i5yXUMAgshcYFDvjusWHq2G4Hth
TM7fI+CkXzWi03oyFhRUQU7H21+98Jwad5eZNVHkHcO0l+XLTzqp+XFlcqAUStJc
tF9UiDuhvC5N0evF3qX+TUl19X5FDukTi9FLjqFkkjQGIZGznqS8dZwbbj6rOzEo
5U2fzXN7sYpg4F/DzVp/PM3LdsWCCBvG5qsOzuGJHzLAPBhrpiM5phjDxdcwhYF3
YurnPQ6xSFwuOrEEoqiQtUwrLfPNb4Xw/1/ep3jckEgY4tPUMMxVDtyYWV8FYq6F
F/9YJhF1A+3YJVvVUc5XAbeYTGLGOls5x2dpGOrJG5lSLjuQfxxCPpeXxmtJ293j
9bYyzON7a8VelBQgFLtLEAHA5OV6w4lG1LB53Qe/Ojg3S0iiAasGTLQpWzPT8Ykt
dF/PC7tFXl7mQ/+AKuXxK/owMKZr0e5Lchibli+3A1jQgMXjhWKbY8tI2pCsRkhF
57SkVnMLzQTd1TPuEnH2L0czY5lC1sS6iTc2gBX6hZhvRmCfvWt1IvZC2v42c1ad
L2MrWHuddGZvklu58vfD9TS5J5F0kspgRKf8dIIRXbzHQPY8Z+BReNm9lt5p7DYT
41k5DAlfD7unjSTNjCQpXD2e1RuZys7n83ccJ39WfS5sVPuaVP4gJvfusEHo7evW
kLEtkmX49a8oMW8AZI+/gdA5cWd2CuaIsDGFxFPumxlBBhgqEqsfCnY3QLfDqdsJ
VwIpqVVxL05mbxhzGyLFe5K1nJldWuHtixDozaMzbSrZRsFbu1WtqhTG2HXZFyCc
dOs+jFWvuCr904zTUYSthvBxfZTvP31UIi1Kj2zy1xU62R7eDyIo5GmD8ulFrpzZ
o/DonrmZ54fKIFnqE9ue3iQmxVfr0nu88VyVF5bcKgrt5q/kTEr+Gd0LQxXS/fzQ
wanoflIo6W1NWbooVSznSibWNepOxuv6rrure9uiNBgb4qYtmjQ28ULrN1WPXin/
JPvjIHKemC07i9/L6s7sldI5O1Y1BNMzkU1a01+hM0yyunMLA7pAMG1BANxsHA24
ZdXFu37tKWXq/itWEZiVn7mwfNKCph1FIjBlDTzmEBngsRwByhU805na7GB6b1SR
XdxFRE2+qWC8XuGz7ym+mOp5XWzot/W6VK1mIlR0EdmP2jGsq0xZO0pAqYbVm60q
eCYWpX5WtZrU3cnbQMBPp2I9s5LE8VDz3SgxE9rJWqeiZLGiiWtKj8THmxmkLCrq
PKsAtpE14UKfQm0QtKXmT/X1vvn6qA9JgTcRGqdYUbOA2qaM1mHNv8xQB5zUOZAM
1BbAVBVAd2Af9/zE+0NmCPOJDThcXVQSoXcHwxRiK0hKxtPQUnBvC7e6uqerFvat
uagC0dvf64ApH3GJcx4xf9/Sqf/UuNgcSpR8gjEEiuMmnHRuANqe8sCRf2QWReI0
yhZd0ak2xx7qiJhJ8/qOlERd5AETUTUe2w+xlekRjb5iyG/sPaXLO/ww8QSTAsAa
t5cAuaMax6v5RPGjvXIeynSQ1due0Lbd4JDXgWmWTkDl+w8w0P+2XiXPH3a05XX+
LI95Yw3uoVdwtS12dBfeVRHaSvHZGI5I9GV4v1JQa9HmKEC/NH/TbWhl5e+cdy3/
GhiP2DWFJn9Y5CQxOH6UQXuvOFvz8jocFCGVN9jzlaCPWcB5JRtA/+Sa0nYtX+ns
Ov5t6FQ9NEmAbNFghV9hnACUwAW2gmMnMCgkgi/0K9efD4raPkTDzR+9CBqDmWSm
7plBkGRrwh+K7+uW4izEMUk4HA1TMZvxoBf8typKFB0Ksd1cAXCHuIrvp62qAtxe
Jisbu32iWq31nerBIvlM5PAIUdnoCajTbtEC6qkb5J+7A00Wuv0j4Zr0eO8rerey
9B1db2NtW/OSkVkYsS/pjQsRSS65vT5qB8eWHZ5aUtONnSJG311woewE02ZStVMj
uHnaFi551vitD6Ybms8VCzfmruaCCPbyZ4olNgDDUXMApmx+O/emzXu+dsa3xe2Y
0zhI7VUger0XakG3jKKPsvDSvZzrt72ZcM/ZfjmKfK6RIPlk5FWMRfsPd+7CXt40
bXkS+t/5oiRTR9HevcSTEl9yIkCDn8HwWaLtiWgir4TD+5LBL/XpqOtfr33I27qc
JqdGwj8+aar6u6J6x7Q1WoaKOTYn2HMEwbpSjjoJBBkpyt5OTrAZVensuAMTrTtK
0hcrqi2DGuXgtDP8MgINS9bd4wnMVuG/IEqkoJ82bvCIPHGHT3wdi9nFZzxOO0Zl
Qdtcd/yakYOsTJDoR9PIuoVQDzV/Id3keletuBguIi1IIvdG6CBV3wq4GFgNbW6/
smMTckK3yR4RHbHEX6+Gh735YWdxwOwcVzCgkB0wCAZgORewMRFMHEh6p9cw/QTW
KKx+JIlzy81c4YO2vllVhl3sNUVyyvuEouQjfSW2e56tCLVNpHdEUhcgwqJbxUDy
hSiVrBIsjqfrPKIcBXpdvIkrFT2BCVMablE87UU+LNnrWU2SEYddKI31927Di8Ha
JNp1NBz4m7T9SEjOMwMlM5j47VWAcUbCwcW5tYcdlkzS78AcrLH8RG3ZwNbvgyjI
FH8n/hZKw48L47CJX0yuYWuLoIYI3BOSXqETkEkxBJzcBewiU6L6zAejcTjGBy3D
HGLY+W2ehMSeryFJe6Yka+yFp3i8QLLyyczzRqgsCD8NuEuUA6ei/peflcUudIMj
yievCh0EzrwPI9QzdUsOx5R6mlRtb1Crux5Wqv/aGXJJoO45rA1lv49bOPJ+kj7V
qE1ft53/kVC9hSfYkt8mQlpW0wmf0Rv7vMXlUD1HV7RZc3w4OGJMrLW23vIty1+Y
pXbm/xZuvBz2WqA9mW8enftktSu8zbthI93O3UDOailnk+0rwonHfioyQ9PVEU5x
OpGRZJchjQNpBB1kj7cpOkP5MphQ8qVCJnJghhCnD5Iej7PeBh/Oq7SR1bu8Ymjr
GTJWIdrdjoKqSHzQF8aLnvXQDietzd4dPAl64ELRNjMpxoEMUviunOB6qnFnHmps
Per6OxA5Z9Rsh3rVQfzp0/e8oE/WthSg0DbmkMnYfg5W7MZFckzMLUFtY/OA+0HO
AF3xEhTgxWAGrU8tJ3rPLwhfLkpWF4Bdeqv79YkqZJzZoVbjYWVDLgQTgSzes+pJ
jGU3ZZDnIk3qLKAyQKUNb8Juxn1FXYtWJj1vDbeXSgmlC1je0VADynZoBlHufQgo
7I4GlYKbNxQEGUdi+8+1HHUV9RGtLSS2D730/hpdzeYP/Y48HBqOZDbYx/c4QJAM
+7UWB27/kt9yJu5MoANaa4hGpKOoOqXkl6Q9f2UGjo5h77t7xABRRqBhwU7m1sU4
7cUZapJduChyfAEpVdamcel4G8gKMvpqwaRAUYtxG717H2o3WP7or+a/5Hh+VKRA
SD/uYo+1YOp+ZI4AzvMU7We8QPOzrUpsr0/nA55+2V3fFTMTlmsjbI9ynFhm0uAz
KdNokPlVcFbH4zQj/D02EadMOjMHEm6hl2wKY80NXO1bJlXr77Y+lNlfG0HxvQiI
Pf0T3UyVKHqoJ8Ee5oeYWad/LRcgxlVAyb4wLnUiWkM48F7M8muLR+qV8FahWZYW
8QnS9+j6UIWp5+PGsWYgIrMIfCIJ8sH3ImTuN3ihFfNEHbPqtbrZKchSBbfRU7Rd
H90a9+f7jeoUERSYMzA6gyyJ6vD/m+SnAbP0b2b0AUMnFIyh9x+FQptLeZaZspN1
QKFnGNXMZaQjheifWF1oyyNg47oKt5a9dTiwizP5CKc2azqOdDHOUAP2OWwlp4rq
K5xu4utwyYmHjtWob0aBfbgV35a6M2sVERmEPsEMI62NxyW2rhWFggMlUQ/uv4vs
VyHblmMb8v7Rj1ai2QOXvpoSpW/rwG756WLVQMAr+CIapbYlF893dWoZNXUBnfHn
wE3Imu2T6UwS5I1qX5Yhq5cJWAMkxIaEfcTFFdD+r9FY2M00hVpGEcvEaIcKd6/t
PuqvZ0uu/+TACRTCSx2pJ5NrNnCKYDDrkYIPbkkQ3cOnOuE9y6DjlxDu0HvyVqRj
uPzRC1liDLXiPXK6YRUi18MC3K5UCVdqsTnvcrI25oyQjG080F0aXHoAgA4Rhs8x
oRNzMHmbh452gdrs0MjTrlB5YDBQoCoDjD7TKEsIpSnCfjR69WHlw7J8fgVKzzrj
Ho35NMgQ+Cf6TBRV2pxm1XrN/MQpn7IbtBhM4brjrG+ShaCdSXvk0H4goEFNW3iz
PERI8N46/exDLKCS2FvnajQRaD0WbW5n52yuwYVbmdZpTxX7+AzjJBTkNalgdHSz
KMU6plFXo6M7EoH3cJuGxCcnGJNBNTT5lntediZH8w//eK9dNDn9sEGzCikzEbME
/YrjwpkW5/aqqRPv6jApeMbnUfWoVc3cjMyZKIttMEMVJIGmPQsGde0SxCFdtVJS
qk51DCmaU2XKBEgoL5goasLhZYMT7HCfN4hOdS9YdgwXJX/Seki3FaHMsj89jgc8
zj2dicPDo13MleF6PyE5bGvwEfQcl2VOQULiXSPvbuLAPgc8kqlQ3cBvve0xtTEW
IQZkk2UVLhMxmxKxO7TCxXAQMVNSAOQstO7kAq6qudT0XNH2Sp/owJNrIrCNiwAj
gArWGfmoQb7nB7YrW4JzNqRe+evaF0FPLt5NCCq5wCQCmtrqoLiBGOo2YldlyUxn
ywwbxIt0NmPk9HFGLcUp5PE5wFAdWfohKf716/dJKvQAJLBhmT8pe7/ru5GpJ/Yw
SkfQSHHeVSH1FoJp8P8m7GlxNUVSGlbGLv6KyC07Ind63bigMHUMBO9mjOITBWCn
96+wuqIEio0xhGIMHBG8sevxsLBPzjvYLF+2xZbIerml+7xXeD+9hR4CGuLypurX
F4QkNWQmyWC/JlEjCv10cBpfI29zkW2+Qdov93Q4sh30Z42PV6nzhqtQ1X+hjLMY
0ewmdJGGutISvhGsxBIuAieSjbWyDCsxq/Lj2NFG4EPWhHMk6XLa8ZWfTisvE1Je
FZizYLssfcO7i+J784Mnt4t8CYJpVJmzfCjq175aRXtc45G1eylogU182if1E9fG
LK76yjzrd4elQTSJY+YBD/5VHo0I2JBOPCITbIcdR0i5h+tjjI7BcsLRu/R2eTru
tsSxpeZgO1SAkrunODjTyOkcDvKVOajJEsLKMA1PFzS9mFy8QY/Wn+zDlIjLjfBQ
O2d2t4JQXPT7o6eQYTwsKV5Guy9HVl3lNRHPjwIvvIl8ZM6c7m0zjHvNAgUzChQC
i2+HDtXEGH2mFJXTFsUrns+NE0SazSsWB88canlEokqeQxiFzFkts1spxsBmoEB7
E7wfoZ6nllDu1ZVOju+4ZxK4PmbS6JLsyne3/skdn4RdXJoCc7z5TZZ8ytHIlp04
Z4+Dr2Mf0G9oDFwEnSFynTVqKQGW82GFzbvpHR+VrIVMNT76GkAEs/Dr6fNLX1jD
IROk/6Na0VdmXXgVcLtvcDK27rKVLdYnp+WWJ+5Lf3wVmxOLDxqVnTVYAqH6CbNi
a/NA99iGDNTrY94Icbfd90IFCz9xz8BVMOiAT9GQrbi+spModzaqoSL+nO9ZDYyv
IB5Hi4kj63025nf3Ihd/+L8PEkSxZXIalM26nBP6UkjVxGLZR4iey8sxqDRDkixZ
I25GKTydGmyE3fUq44Zv7JIIfa4k64TeOnwGsavF835GJD+XJi8ho4iJABsqRhO2
VAfNHQNn8fwcidZZ7YEEbUTrH7iRaG9fCIsvKwWxQt44m9kypK6T7Nr82/j8rmzZ
EFSDuUBHS655Xuyg/li3beUY8rBXFd245LuSK4MOOhE8KvBaPO73ySAYeZoAkJEI
3JDs728MSzwTaUMSzoXUNeqpS0E5fn2QsVxRvZej0CTRcyWZ/1DqhPgRsClHgwIt
lRXfvs+oFibSqIBWKSY5NytetieScGIfuTgJyZPq+CWwTfse9i90/pS444geSbhy
pKCxji+baqJHCy/YG+M58SLKZyqaHNRYh364pO9xVVwhZlP/dmBbkJr/YJ+7eJ+M
55h5Y0IRhoGauVPTgeH91raMxQY+YBswrzw8PIN4BjfhJCYeeSrM0TWanBkoRhEL
jrSVw41g0Ob+y4jlp3fkqDCHJe78yTC3NdyXMppvqWXcsKgLPAFdleHPp9jh13n0
g7v6s4gWZ5fW/3O3yjrKlCOZmc8J9+q61R7C0tK3k5Gnva3HcNBEvvdgUan0WM56
+zIRtIwgf4bX27TxfoyH2ggs5+0SDjZBc/CdEzz/1AUEhZ8/x2wg9rUimQQ5VlQi
xBJvHa98EA9Zn+lwLD4VRlTwczsba9vr8O0p63HRqq3FSYiwpXTfL2SQh6/gpxp6
AS7GTLn8gu1oBPvAqPNN9XHsR4Wt10/v6c9T+TQx/aqQ5U9b8fQ2EzLGGWwCwjpA
rniiMPiGb7AucqYVEW2/7nliUxUuvcI5D4jTcYJ1ziGAJ1Diq4bLZAlpXzhN5iI0
ByXoJqkxa3siWCGGIsO+R+54+rIOA6fLYMosJKU4rJ255Ccp6flC8IzdoRPAg0qB
QmJx4iXoP3w9c5yTdntBcqyA06lC32NQLalEqXfuuy0yLFCcSVZZH68Z04SckNF/
Yrg4N0nhA+MtOXjmanPysocpK4LkuaA1Y07/ERa8sHV7XNhJLpv3xLKMSlWMWvyR
J8+a5f5xqCS6bl5B1sllqzysk7hShTI5p5mkTK8otLikS4WQjxPRseeup8j2+Cg4
u5GVpoj5uOiy2n8m79Zyla/EFyD2g7p5mHdS4AvcVHhElIzLHOWrIg6sbg1H282u
FGAbDW7FDYHOKyeeYEG2i+wVNUsY3+445Po3eZK0wmdwifQ6zQKqQk+UnRll5p3Y
QEDIqMo/jkfkm2AgplKZ5zI9X5IDgMkh9Do3G2QVrQnYiAyLppG26NE13TaTMcVm
H+yzIrFCLPKM10K6lCtNO4KQN3EBL0Hn+HA+6CgYRyw2mk7y5MVDiWbuCJnM6FzG
iwHBbALszToRs3SPOvBik5XR+hJD9MhfxDxk8zswgnsF9GGYPiFTz4Sq+iTOrAwF
a8JBP3vlCv0LTi4NnqAG5haa6UWw2R00iS3vHNJ2OeNoR9ua87m5cRD9nYf25k4w
zt4PXfCW2oglq31ktZ0jV5LfjRpJiU25iu008Zh8HD4cGoyDFYibXMtd0metskCc
2JZ2lZsPbyfZUXj4Xwd8BrBjBfpP25sSViBBjQiMQ2lroolYi/U4j08wWMU7JwkL
GaKVKCEEcrmPHoycKYRkXnAsTHSyQlyhe2qikdK4NsudFL7Vqd8Zm6ia2ncEBPbf
yA/hY++xJw/BAlVFbCBj5PNEqY4ylpyW+8aR58wOpjDZew0WBtRWUPtCyFPZKuwf
bs3hTCNauCupgq5dSQgUpScl9ZpoJUIskQD5MuDy8o0H1ynCu+Ma0Qp06JuFSZav
gNvIGW/33P23jVKJ6UzdrdDjkvp5KmtUeXcFDnwvrMk9lib2AuPARxJztfwfgFPQ
v1kwXtLBzgkFe2BhbciEc4einuqlNnCGlj/d1GHDE74WUgSMWR7R7H+2p4Q4r+jp
/iw/k6cET6z2DR+cIgX9gn4c8CT/qxb8kueD/gxcm8md698dHB4Yb02PpG9nyfI0
hTg1Ydpt1vclFegtiKEqiQcVIeQx9h8pwn8Rlu7MzY8OQ+xY1feG0IaDJR7GwbXs
yP3cpDcArWR+znLVlqDuNecfRWG+sWotoYeKBq9msP1mAUBS3xc/gaBVzk/LIzHE
tgK5yJP3vA84objnbRhn5Lyw3v625nXmZ3k2JLDcpf3KThXt7cHXWxUhm0ne1sur
oEN2MB1CLEfnOvIM5/zNqZd2hoIdjbC5ICA2gNK7WpKoKPNzOwJmsZkObkiwTfX1
yhlTFSK0WGYZSxvwNAx+6yEE6Kbaf0m+KxZtmvE6O4UCOVNiO226NEih4i11I/tG
EnJJua7g11XACFmJ7gSHjAf/ihGaK52jpSwW0G0jJI+UndM6xwvWpiAV4rRVYotj
0DOubHzhUd0lJqbMGQJRuaD93YC22GH7WdZ9vn5Nko+asIErKktjiJLoVgB0VcH4
I7EqRYdskQUY+R2M8M2abC12OHUVcU1NRH8K75Jotp+CEowVffXapQHMzCcOXmkH
6rU6/EvFaFEb7csWkbUVS6aHlqnJ3Nk/Un0q1e2L2s/a/JdrSc/Z567ep/3yoz6W
ave1SwSkzMHmgmhHh/IMKrQo5oi3UN3ZjF3R7jGiPyCZvD0S21Zl7go1s/iLSSHC
EW6yHFjTVqOK6lJ6i/DTdpamAQehUIeg+u9IrEi5xxfxa0o4ct70I2PhO10RR8Rq
jHZ6pImqeqykoc0MKd6S9kLxUL0dGLhW7RIMAUeUAC4GOkgFrZfA39nIbR+RJJH/
oGbgiFEcxQWXIFdBxMf/8OAE8CoTz8/J4OfxMqqkbTK/uPNIh2XQM8Jg5aQUi4su
os0FPOya5PywH6PAZBxwBixKgrLrr0S8/M2+4pwRatEGcVQNZWk3wujeJNdZuUa7
XbFekzM/TQIMvU83M+rTTYPi/en6gm2AAAu0wPofKkSP0GahWnGmvHCbiJ+N5WLx
7fxJ16jJwiwSNdgvWjB6NUumnYiCpHzAEgaK/6lgOBwqpDZ43hLFof20Nasga9VF
Wf03BEFwgjGENRn7Nhxh5quiwtHXEglfg7NQQZnunUJaIjZiDfyyXPVg8vtkXCz7
+vAYh79MNs9OHnZEW7cG0RzHDZ68WTByZfNS5ELQBHXV8RggzUSgNqk2WeIx2b7X
aiThcglwADD5vyEY1IqVc8y/eZeIKkhmh7J4tHneAP71a0y4eHwbaWfDL0Q1Px5M
maOUalJ0L37/exaF6pLyF7oyFfubTNxdCKtgpeQqtTXM6G6N1Zfg3n6uvQHd+kzI
ijEyGsqPjcJkfdXMYaHE506FqMs10yUdVwtiAiFVTxIcowRmtWp7QFnTYOaUbOfQ
53zT1Pt/BR2zARtkyMudt4zI66oI0VUdVpizkFBV+fXbVzA7RL2BPLYu8XzKiF3d
AgZ5zXYYWNCDcN7d1BmkditcUJ/7zySaoCzoryHZZO7vzIWb4JPzfc6Trb3KcSBa
4UJwAOOwr8NigcpHmiekRP4e5AT5bwOuE9o0icD8MKtN0myEoh0slzG4AQTSlW6w
RV3jIGBlgvj8XljBZJ5cB4CCFSx5/fpUEdN8LJyy7RNa2AcM9w1ZCxFLH0vsgMrp
jhNS9C8dV5jcQFl59welKKWq1cGgEQ6k5QxcOzjA0/jKzbSC3GRh7jPx9Lrmyt3B
P7BjuhXatTHlj1YX50x3HCdtXi5WzXT6y2gW+qbC+tN7BB0zYn6/4qeVPulXIFyB
oAblGERsRX/wzKjGNHU6OhMPrnBnWIV6Qd1wttQyz1BkzVodk2lepNukvjxBygcS
QPX9e44vw+2MMiaGaAsf8D1QgTBZn3E/rBNMoscGqkQLxy/IZ9cIzbUzrC41djv0
XpkhAimUiC9NecsAYEqjsYLJK9ez/WpA5kVFGopLFR7cF839Qk5hELBOXcqQODws
B/JoKbPSPuhbrpN0/6qlJXgWHAOaO3W0hpwcCv6LdkjNMAtLOCSlUKWXGTiLay/U
A6sc2+jy/NynJuO78lrhUxH8EGXcVGUefC5hiCHgRUeeXo5bck2rC35Yl+Q8dr5z
+eJO0H1dIUs2T4nMZJ2+rKuxZygkogNPnFlkP3yFnQsy9LoKW2E6+JO0UUBH5Ake
PQ1lzBzXyjZCutmfVTI5oGnAY6HNcEO1JY3ai8P5xUSMq9NJT8Is6KtAf8loNpx0
YF8eizLwO6LPd74El01V0s7zujo5t7Sph5F/II2WNCepyk6zTIaqf5r+ZgVcO89F
+PbbYFZiZJWi7jEnykzM4khANmwzUiNaM6LRDV6qY/aiVe+TTwWDAjPLGSTqx7MU
/WIAX+ClKR4Pag9BcdX2pWnVX33s5DUAHQ66lAF+QDprf0h+72LNvaSN6rsBoHZ7
Z8/M8JZPyq/MVWnMVwLTEOv0ooix+ntOqcz522JxEtd9K0PBzijTcqbjZt99OH8u
BvLdiR3hcEHFIdzmo14gMawCiVoStbviW+l1YmcLDVxJLHLPId14mHoaN+vOdLnn
CmNrBJLBRlno1tBswe8iGSA8gvLBCOPqGGruAfNHKIrnZe1T2Rib0qYCR4Tv8xKO
vlLKcyzab0pANNI3rRjmpDM4ztBNwQiNRdk6cQuhaYpO89cVmIPFYxg+nNo004fL
uGv4by0SGFED4zdUtLXcQAoWoZkwHR36ALOdvr9I+hr9u7qRgwX+TjoXbclfegRh
XhbD/CEHHhRmdv4fErWlAz4VpPL2Zri5nRH3vrlRKxFV0B4JcH6M9s5x9IGF3zU7
z87DGgffWy6kHWgO/Jz/laqKHGP8cnTsdia9KMICXkMaFkmn6nPX5OdFkL1AVhrS
mft1hQcCWwhPGJnPFMWw4vDdMzAr+w6okp4J5ZMC0dKWyI+abLiSpQX3Mfv/6DbS
y6KzpwwtPka+0QpPahL6VfUAKfOyeVVTIAtvOGKRaVnZREMJnz3HCxGlFZ+AhcSj
3+HeZ2H/r1S95ImlFkKDTttRY08gBGqsQw/icibFWUzW3voNnZkZCeHmM6CDb7MK
AbrOeuFOSmDzHENLLsq36HAuN8WFrV7QxwsHlFvPs1vLM2KDth40+9WUEZAUpKTa
ViWynwRrVdPAxyDWYAY1hcshIiVfSevkVlo1c5Nz08NuGslUnHVATG/zdEF9XmH/
h36dJnUDIcYLTi1KKyFDeHvz3rTD36121dpTaqCWqi4vRsNGLDEDuUaOB7mUm0R+
Cg1bYjItS5o5ZeoEW+IVDacLp3YudGLcGh/nymFdnls3bay+OCblWtkw7t2UgAuH
PMDPUz/6MIlsgGRIocWs5BFEroUsJMPAtDkk1qq5j1OXIzf0/mOtxct3XWNwXcY3
U0x8FqL4M/ThsWJkNxovhqdFGyuNwQvqLgVctATZ2sP13sxmZzbBdJmgM4r6SP8F
wMNxAzRk2y5CEjEJ60bC/pGN0SJK3GwEPqCnGta6L8hNaYKTR9Bur6g6Tv3UjDaZ
K0mVC7ySjKyRdxme/3mI5NT5QeyqyTKluWedj4pxt8X1dZqIe+1wuKbgksW366xH
rNM9kMlTFJxo12rstKr3TYfPove01tbTC5EE2PPGLFTwDuBUqIPfybLygYPhNCxP
suFRchxYYFptbV7z2xqhLP5ciyPwgP+zf+h9vKj/8Uk16kz3x98Q0aaAAelxJwHM
Z3vIH8tBXdW4E8NP7bpsESEjbcY4HGqyonxd3bdlBAcdRXuTu9DkPqcvxH1Ehf8J
gUtpqXNsw6hW3C9iXkUh9CUpDgTHdOT/VIz2ZVPo1wKzM2u5UGV0kH8xfy+EtbsY
modWLyP8gsq8AY234X5ffeQ9hFtL8JL6gfvAYYBEo6CHRZ/sD++lHpgSWzh2vRJX
NTL64soWebODhOtd/ahFTyeV1CC1QOHJZ04AH5G/ihC5mWrtXCh4+Tm860LZKD/6
ZRr+y9ZlgHFI6asPQUxPV7M/36TExPbuTkNy5XIj4U15edw5QCboeK19rrRYXGos
dUs1WHVDdT2IU5jCY4qXTT7C0wjtuKysGCY7e9iIq9pbHzazLYUyB8s/C2kp64W8
cZfpnSBcJaSYUDgueHqjz7vq+tIb0acfSq1iFuEIzmvZfvQ+AORdAkA+kKiTXPZL
3CTEl7QTmcmAFxD+KRVCB7NdRgBm1zixFDS2WyQ1Czdz3OQV/02/KJKlTniK0OC5
YxCjgTVK5G/m4jqud05J5MrGm9CLI65WsSq8Fd0uqVq1IOZaj3clAsuG1z+UbNMA
APwErLllVyQp80TbE4f1/X625sPchKku6yY6K0gBsmu0+umLgshzifDsgl29WB7W
uu4OLvHlZDPeM1bNGwJdVR971OR/0nHIDdoeuGJLyQyoMjgsussgaE48bp6Ar3S7
BlGASMKySdDJGzUVCST8T5PbNJbdPL+QbHm619ji5ViZhALBqV0VKMyvr76qyAQN
LC0HpFIDcXZ9+LaXjUsqi2raeOoG0s4h0XRE4SocCjkwOzcCB3O4SyHAkE/02Vqv
pPHCwrfMyAJlCLZ5HJ1B4K46+g2IqWKbTvP3J3/uz5AYbfdnKFim2ON4dAoBuQS0
K967Br4V0hPhu1noyItOjJMF2jiIYNdKGQoJndNSdA8HgEZIw7AD/o7gnDfbl1yt
+nckIInKuM3S69J2rGvlNl6S/gyweBBm8b6oS6F6QEyJYuN2WipHdeiCutAXSn3d
otarhXXNDNPYQ+4MsaEnalOKAQIgmiUN/8MHa98eP/RUTMWj5CMlkOE2DCntM1xF
z8xai5GXQE9BoM2e8Td3rI5Z6EbEeCwMvbMGRYZ3zjVDW52K/bXcyfJoRVsYmG7w
er1yTaPykkARjvt5mKrM4I31i+0aicSjzRa40reY9IRY+X29ynuDcHFzgutqnCw1
OOcNJg+oLjf0iZRthdlSBcJDeZeVahKUxk4DPSJKhLDJ0thYgGwDEIhtqI6siDyo
V6g6KJLpTQn2otpebrU1j8muRyJqyLTa8Tm0D9HQm6OcXaFksiGU1sxHZ7rOTmqt
q4pS6Hxu4n4DyzUorF1h6Gxs+ejOj3c6i1WPT5XHv4Zox6yCGJoWX8F3xWXFTLDL
FrNE+0yYF49CdDD5lD7TyBBstGJYqQZb6uNU0zMjtOFgvwjonaK0gmUm9ZRV/hWD
5ZYPfcrFRx/W4iMbsW5xOQRdYAxvFetuCjmNxw0vP+1xBsPL9LfJKh+l5RwTbPyW
EY885EeFwhtqbqDHNVgHxpX9fgkX7eAc9AW/EnCpRBrytxSFK5hfQGE5Mavg+nwm
d6O/Kkpj0hSUEUA6/I+chJsksMYu0gCKL0kP7Yjogp+KWNlFOht+/a1VCe08s2Xw
GluqGFQNz24Z7KXwTWbyHJQjF4DtdMidCATstaryGhkGNYER0RypngPDaGPcGKWT
qjYIgK8u8DkufmFkk7jWuhnBscMKjmZv6YJTrY+cfZjIlIzNMiv2e2xW6nqFLChQ
14xRpB+y1lYITXvVeZB+EMkKC/1yCPWR+0RW3nj7Tm9ofqzvhl9iFhUtP/P1P6m8
m3Hy2OOQmbEhTlxO+N58S1gYP2tgTsxw7b8Y1DcbEFwU3o0vAuVnOlMYsUceZi3t
Q61eEfno8yv9NfxdnfQqgmZ3/fuyhDAkp1ofdcJl7vEBFV1/BbkJC7ksv0LUYDUj
1O8KF5xbBjgJ7MqdLRii6aKpLVJRt3a98rjFnVvNMc0de2EGWCsAEnScVeXtzxRD
EPW/EP1yxkw9sJGPUko3mdAyjTm5N88jUh6e1ZMKdCl4ii92RueuIZeS/TZIRKVw
9H+Uzw2HcB/vueLynFVslmfzrXbrV5dsIAGLbaf0qqAQfY1JFkKujJ45fCjAInlU
5zQ+aEQgT3NZGXrzXV6OfwWIDbre5OdxNVSQrdw2EM3GC5MhfCc7fpl6xxycWMi4
ZjOTHY+lH2laGZxrxbktTQWgQKFDiEnDLDAQev4sg/3s5/mA0240PgwDSZxcd9aQ
h9SiYuU+/ujwXRFXB3oX6JTj5xWhqjswXHi2HH9+v0NBQbLOozsq04aJwg/GHDwI
Z55dlnzdG8sxwTeTIfV8eALtIOx3NO+XDB+kNWPr0KBH66ahqzrrpt12+owVVlG+
B+93CBH6qFbMTCt53Gq8NwzXlFNtxus2ayh4O7sUC9Arbe/FMuIxZPeru1SOVnOm
0O4fSmpeapf0kC5ddGSFBGZvM13u8L0CO5LX5+29PePGI1hTThtpvOA+JS9tr1hK
gY0s2dCyCMpcUihPKFWoHTHLljQ3+/LwwCOnHYsmE7I6YIhRVxK6tDEcZ/3jG+/3
EQ2r27whtbKKAMU8ILZKW6NfymEHPFziJBmcT9F71sk8mI+wjM05k41B+rlHqcN9
jTTcvSjDZaIRZ8C6HpVeheKOXdM5f/t3EUD6rTV8jZeXbfRpwAqDI1Xm9+3hgJvv
IO4gypfK/a/4L/R61/72UZyVfaaV23NBejHpcFNs7/qXlaFrN6vbv51zn6YNmXAv
snb2JZyVeKcjfhZ83WBpPMA8hmtf8rVQnzLNW5mWDne9hHbgVCO6YC0N9f7xL8zD
J6O7HH/D7bFQqvoEWMtKM7EKJZVa6iMOGCFiA/YC8e4uB/4TT/VkHxfA+kch3HeM
bKT8N+2Q8l5gDgubi4Ye1wm1WMsbBEF53xcg8g5kXd2lCwFEgL6TFTdmBLHDjMal
cxSZNWdVofJ2lKCLOw0FT7hp+bLXscciJtDziXUySo/cNkTWKRxmJ2gQwYqQXTKo
EAWxpxmKVaCwnwSDepmvz4laE4H50nXT2M4NsSEP9fAhA7fO91mIS0GyTspvE3XT
mspi5WNr8dQhaVn1Ktu7STp6W8Dq13tXnAwRTeBQrf0hAT2rArDv1G6icwy+Q+0c
MRcV7RbUfx8P04EsP2yTirkzhBJsFchScTrSpWEokMwpMCwtLAf4c03clS6qp6Ui
SyIuibZ4K9y8NlvQKyJ1UW5GMmr/p0E9ng2tEnirQ1Qb50WZnipYbIjDhDTO0evv
cX5Mdc/mU26y1D5tGgtN8kjX45lBl9hJ+8d187pIV7052rBxvSLTR7Fmi4JGQROB
WDVwl5LSeFSd5m6f5NSaHYIN+ogOxLTAwyTqt4PM65YoTMAu2AwMLnVLqaADL2Jo
zRhoFEDXqdSUr+EidNuABYgfM6+P817+eFBDoPmDepmnD5EyiBiPj5uxuUSwZcG8
L7NaDrVQ5Hez8Q9g3xcY494cIA2kYgMKM+bvfTPTrbtbzRrydVjSePZ2td7nemS7
EukrtFFHSHyziNcMM5mEhFjGzlIBboe3C619l2ACo9qpedhvdJ++MDbRlqg+3szm
dcULcpNcSoia9SpMMSyqL/31nQiEaOfX1OcHytSskL/f7xbJOCsZ7z0u592TjOIV
QGnXUxZQpLY7oJEdRQOyM0qBYCvanNYYfCug3xR0XHtbqxOD7px3ROCeJTJnAKAK
2OpJ4lHMjZ7ldpDAViigIe8jAnrtPX1HKW7UlgEMV/ylFEASLLoMwUmJj5Bo3xyS
oLGrNSq2b5WMMMX6jLNEkdln94gnyDrZy/Peucbc8NgJvl/0cUSCzE+34W2rDEnN
iDISGPE8yVN5NSeXjxMk14uMxOhPlIn4EYx1EdhQFta+yytnuOUbYVuvC+3XrOW8
+yHx4gY/yk0tdyAZEE3H3mQC6HT8r2zr867TIngXAqbtts+ACqLn+AZrpKdwSB+v
uRh+xSHeSdIdR9+HJrSuKubdOz0etBrfU7C6C0NUgj0vh5RiuFQfT0NNwN7zVAu5
DppMTELrHuOi9OPJG51UWDTppPpObgxbp66cY3jsREeZyn7e5rL3808vbjfWXgF8
DKrHX5kVkLLM2WNPDWGkOZRXXZEWW47EY7osjv9imfNSg2prfYQQb3Br5yJAP72Z
RAgtJR1NTJXR1u+J1IqT5ljhq342raYWxFHfl/HsWDxWGfIOPVJMXXAw2EH0jXtJ
D8ncDUJ12Z6KEXJCVtB4q3c84NlKTks9A8/tPr0IB7eVizy7mbymJgpvm9z8JRvs
5e8FTroabUEIfbUh+hxO1O0SuP8O2piLO4gwNgZ8OOHA73rpDULue1+LoztYiro3
XQSof/goSU4LCRaFxmO7FI95feFw13G66y4ftbGQG2rQElStXpAEuyV2uMTUovN4
SLJTBePmztgrae3+E+FWMrehSCOP4EQKWoBKbf6x/71oVeLf6SPjeOFq8ovvw+wv
ZBKts8G3/8PYdg+4lQ3y41B6MCEvwcOT0aNEksJwbvoTDX/kmrQ2dVJ6y0MVJIxZ
2yCWdXBETKZzAQQmFcHBQd2Pt9bCnXs7JfvyN4duWBY55icvbuHuFLq6c16BNdmh
nw+D2Ju/mSBKiPYQiQQ+LKd0jO8hgJSNaHYlepDEd7NM48xezMkhPV0JpJW+TzVy
mSjrhY70/6m1Kr7ndTmrw0adCeEqGO4mU0dVY5LLSX4rVz8NXXp8hBeXHgo3zOJX
XjwVPZkavrAzxzbtpoFIhg9KQl4ovsR/QwOxlEdQ2gRgqUVVX5TixMD8OpfC2aeG
Pqt0OH07mV2ddrSaWbCRqggs0jmSljE8GJ/D2GWkc8kOQLFHBkuM7U8HGXBrMrG6
UemjXGUhG883Cv6OY5tNt7cnxgUUGAqTiRC4GvFDJdAj0hWuvVVB7Iv7MgNPAqOI
onNG7scJ1XnGv3BJog32rvFWQgFv6leZLoj0vsi9H0R7iRIePJvDzNjvk9FaTIpx
71uIbGozpkAGJWC70TT82aKzRiC2EtMjEj6bdGmJEOIv3CidAH7HoYM5fgqH8zd6
XutdufdKlnkBlxbT0DOhqIPIs4gfnfFiUrSapJdjmvIpE0n3l8DU2jvU1BtcYEa3
baVgjzTTxsD97Qfk8OHIh89CpfT2HXUjvI26BXDAH+S82uwAqJf6/hRZN3inqXZW
ZC0oBxUa8AbbfOZhe1RFl6sUmzgJ70oaBWX7MxQkHhk/KDppyAu38KwxuDmB1F4r
ivX48RXQRugGzKqYy0aCAcZJ7EmejigD2g619SYJjQ2bion12tLu4p1xRVb4U5AW
NB1vZuExMdKVAtnKXMdrgZ+N3sct2NLe1wDWwNaX5vIrsaQ7pDWV1CD3EpdkTDAr
ao7q+vrM8YYXpdk8xJWf/Fmdk+PtTc0dxjqdock36M6vudiIpuJfdKkssrluEbk4
wq3RbM+rc4WOJrwxB3vby6wI+jVOsuy9JezsofdAHd3FSzVVZK2n3s0jWh5Fc52r
SWVhLu9eIcFU75Gim5LNATMQmRAjFBhabqia5BLXeWoH9/a1spnpRio52d7XHr3p
RyqvlHBMKLknMpeErEjhJ62OZhwACDI2vXCyB1yTjSP1yiBX48wlLifOQMyzRerh
tp/g4nvAQaOOckolY5HBk1H/3QpWR1zD9mLk4dUsVMFFf2ci9I86IKVY5bZisrqY
7D16938oJGxSw/VyEBhzG6jynXTQZ13gJvyy1JmbOf3lxQG6CVNgwBQEcnQL2Vis
wPGta4ET5DDTxbMgxq2mkwlUJxJVC5dehve0NNcytnjaAdNbdCdVyMjqe5lMFKIS
R2OO0TT8tbChtAoKBk5382Ue1ffPUZNBGuCX0CspU5NDzRNRrBbeSMXEJA9FnQWG
CUEYpemj6zlP3bNbxrB0RrfWPgqDNqmJSiOaGEyYFd2nQnO7JptNQDH0+ieXtdlv
if+wSRu+Kjcf++Paj4iKc4yJcOHoJeu0RFLU8EP+hkzWST/V3zwrkzAY0XoXWyps
Q5HKYHpKAEuto6ZASBGpX972EOLXxUJE6tOL7rL/JVDxw2epo+0BZ8sKyUKEbXLP
QndiGNHfI3D7rqyyLOPg9soqNQNu3l6gq7akVh6kM1cVjW2PFsGjMlT3DQ1RBF8L
sGvnFvXACI/A60RVHDhrZ/YA849G1psmJ9HwuxIpZqqwEt+FpRVrsoXAPUe68nCm
5/1u7K5Tjm2IzCaFNdexy0eyhEI9sCdSoPVExGNRtDd8f0GbHwtWjZXDiu7ZWHyK
HN1L0TWP+AnSx1vtswLuUg6sOo9NXA8leiAloXztfIRjCdVnABfaTJo4nP55gXtc
2ACs9cmjLsDwIvZNsdXmMxy7cQBpuZljm1JtW7PqyS075OeSUSuKnrYZj2oLZWKK
kh/5nSDYUloC39Uy3aPKvXvMSQ6qjfTYk+UKf9XYxfHb0fs7IAQ2q12FWOcK7I/M
fnXAzPequlcsB+UtDk7wmcchCd3bWgniVyLyjIEOJlcDSesSREF9j8jzDDRs2oSo
3EGr3RcBhOU6l0m59MrnBvAFDZrm4xIrzrM6HunTHvxCfOYwYoknXnOXxR8bhMKe
rLLkgdXl0B8frF1kMJvFZSQtRIyItP9he9kWtof89lTqAtLGuSvE+JMXpDa0WH11
ccT9MaHhU36IH9onxTnihRCzLC9ylDkUJy9M/sBDS8dvVvtMH9pKxSiZJ9kg4H6v
e8fhHWgxLGA62gmSUeGcOis63DyJaLgOoCD0r8dJ0hd8TcbpUvCiqeuceYYMGR9H
EmI71aTjMDko9oUUoeSzVQl5fc0IevV8M5KUsC/goTI8bGxa3qk1/Th8NnP5iGku
eoaw36T9W6muK0xCkWmbNt8tOSZi9bF3bXwiJN+v6W2st7ogxDKTdEZMTFTglUWF
E1ACXTlDZ38QV+M3tltAMqYrTNCC54TcUnNfuK0EDTQmad/A8Cu/UPgJaYwEkacf
RGVwhKqlVOqen5pz0CI+dT+yOuW9V/zdqD44jfd/55ubrDsmVBjqIroIA18i21gB
tsXhUJTDU6s8Jlyehbc8ou1iQj8kTIjxtxQjLI6y/Grp+Y0K4BXWZV3ErXW3/pHn
LboNHYBRymXZuMbOIwTIHhd7hJqj/8m77InvDBI2s4AnBqrkgTmC1hkRFHg7bSEa
VixbI55tffifLN9S3MFtqPYvS6IXmR6HyUv8EqYHWW54DZgQtFGxaderWO4aAFrO
dNWfmxoC/jpkRpG8KnczPrTRjnl7tPmNaR8n2g0n8zJF/GyMPBEKGgKyKguFcfIU
qwyHE0OZF2r2fudVepN3t6RQkb879bMQr7QEFNx/ZAh5CSDSiTX071jLf0AH0vCY
cPRL0DK5D23iZCRwpuWgyjG6hi4zOxadkUHO8vK5QDdPvTO3ZYU44OZxsVRu/6t5
3Qsg34RjMryCOGcUc27qf/3couGbF0YrTfTt9d5Yawb/cvSvdmkNQ0eQ/2sb3KVx
Sk8Z0cy9ReYeTIJaBeqXp9i7cP+UrFgDEynDmcnD7ZtzYL9gfbQqQvj57GmjMcHi
6/tH623PFEPkIW+Kb8Z8+Ie3LCQUq6NQUi/dn+KdyE6gNMXys6UPaq1Uns28yq4l
vT/gFa4SNtetHCgVzzgkQ1vwTjdUi8x6q8GmNX9+ssdk9XARJjsOYzOAweSeDW+6
3VlTDsNj9r5pEepkFACAV4i+muZCicINSYiw8C5qpnVhqRSQyTGj5KHFq2qfRYH/
K0CJoDFUhulb2iV0078fLF4oKt4Lw8CUPRuaE30U5+xlYA1vzw6hGbstCPRgNEYe
JT/+RTpSkT+2mW7LjNsBa/754p+VfUC0vsQOIhWbRd75ceP24sOfoWHchgU3JIxp
TOv/PG9iceS38+Cyn4f/au6bH1dq/yFCe1vhe71mbyy+tCFfeoOlQoTzntyKDcVa
pLh4w3KsvBNJSWTAmnKUmwK5AzahbGTp0tbkKCQkMIVoXPhq9ByE35NWpCOCiBfm
dsgh1qk3Ud1rLYoyTlddII5FUHU+5NmcOW41Frl0rZSYw2ZLuyGZYjgf74/xeLY5
F2XRBDsjWMuTnkVAV/zRVslY4E4F6TlUh/uVKQW7ggf9ITTyZBGjm1+OebjAnBWd
VHxzp+5l3WB5h3MTV2o2HALa0ueiXVtCzfYyOufSIXRvSe7pOxSUjZqMKFWJrg0O
9v2P9uXuCKb8Czd0WjuvlmTYgqtQP9JyqeXIWN+G4Sp+hfaFnTAYr0Q4EGxQS3br
XHrbPFlONJXKTtMKvXWWkcdixYC1a5CGkSzCtprUbn0qb3eytqkp6FvsIzDGQBzS
jcNJyfnJ26DJlbvDFi7MOrzVSKz0qDuDN9jeuoqwam3AD6uzq821UWZQN2tZQSPl
CTiWajQ5VZ85lJaraS5svPymaxBRfQbyCR0wvitpoBVbq5U1kGGlWKTZ5UF0yGPu
Ic8DpB0vRaIkBgzRHX5i7lXVhFUs85wZAzS4AA7z9QvLYn5m42WSfnPSv8hvePa5
rg78T9d2xyYyG/mFgDG5Vx60xQThtyUqk0GoK1dShhUpC0t/uNz5zmx/ppNr4YNg
Z9V9z5VEyy9q+P8uOSM/mR+GLqZeGtX3cApkM4OfWez8aU4G8P6bH8aecnagPFCX
QJzbg7C/zGMdB7UHYa+QOLjrKM2lTHWptaqlLhpFPdYE25+YB59WTWxWJ8OzSbco
9BYWonkUSqz0owoXldzHKrRiEjSUnAV0korDOrdF3MUXnXVJFQA3FzVcLmQOWuV7
D5jgoBPpobM/X+SebFkcwElQij17em/li0uHwhql1tqOxm57HKePiLSyM+RT9VyU
NE5RG8nR3iIKlAlSPgjjgdnn88BEM2bT47Z1Xs0I+4Tz1OBLM7py4ST8sapVwvzo
sYcVTTYetP3XLXNihAFcpQhKaJ9klkMz9JuYbwcVo2twik+VGMuG2ExGObbnQQPK
889n0NvHK3mdCeLka0L2iwTUtg72bK7Fk6t5htFysDd5gn/nR9TOoaLZA3TgSVP2
kc5qp6c/ONWpO5hfcjtL7e8H7MBxmjJcUZFmXMeRvhG4YT6laT525L90wxqiAPM9
7luCYQE+VeePDCAhxwlZucnOce2sEwOIFomRDQ+KT3ozrM2kiSA/h36Kj/BmeYZW
2Np80flaCUrt24tEdmbrxciZ1UUEmQBoVLvgItNMfVjtzRNMORMcgSYVNlsCgxxE
ZChOE+EWNUwHwBygDEjaGNNb2kif50HfrVbhsRdoqVRSgpibDcJsraOPji3qRvSL
i2RHi75Krdlu9xLgN7bX9FHCPQlCidgSJlpmHfRhplWny3kBJXnEbieb9I1MdqCW
6GVtZqAHmfqPo+75I9xY3T2Xo799w7FxgyzOlQtopbLuYDTCPnJDkP46F5clFFfQ
yd9vDISWeXtfrilGp3KZZ568wl19OtIYPDFcbXKKcC1IsKbBz28lory6aj6yd8eM
x81YaKg0hXYuVSq/vPxBgWlxylLCbLjNKlqWCDSdTR2tU+vJ7iEE9Xm3+SdXnT0Z
6LZcaTn8dsfZxGM763ytU6yzwppZpzLrZXdxmj2+RozxpxerLzwKeioo9N1rvs8J
3FVavbBc+o4XvQg2qbeLHAMZ3hHfOhJCEIPehX02WclYWIJl+atfgThnMP9Cj6tg
iZaxRP6kUNgbdH3IRV3ARhU7Wj472AmdxEyAXO6ATguZeO5PUIiwLCX4o1uXdM+W
P2y+9Qv/fmglzsYWfAiw0jzZmUKSqWvNRseC/ONfCxJR54emavoGJhPgv6g0b5iv
f+ckpQijn3nTQciDRuY73IgMyULq5Bj61CaVd9S6+DuC8Cn+VYkYouu585H3HlrU
OZZRBVi57A1RFjRIvKTFhlS9wFS/uFklgxw9FwEpZpqcL3iv/pIa6usQ2Ic+76DJ
c6RE4+dsAcsLt6zSk7WIV2QMxHB85DF4YkAcRjSej8Hw/DHdLOqhANVybbEAf8Yv
azxvv5XU73lgxodqEX78sm5je/LGMOtYSqIaEpS5YlQmujanIV2CqF5NA/P8X4di
Wnm94qkDH9ASs6pP+W+Oqk09r4vnU8TdAQBXmbj42Ab3VeybhF4iaLY7I+pM7tLM
oT5S06rXkyQKLin54d85n8TP3/Y5belImQLhZ5zSKIp+mvsW9wgFSJGaWLbfgzwP
rByUvrMuJjEH3Fwq0zWowZtgoxAOAHqdLodHZ8PeMxjAVS6eEi4YfLeoDSpx0Um7
U2WOAQLxemwOwUrwjveOJHlwVvLKVU9tacF43FRIEKX2I70FbYC+50pkwtjxl7WJ
`pragma protect end_protected
