// Copyright (C) 2019 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the
// Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is 
// for the sole purpose of simulating designs for use exclusively
// in logic devices manufactured by Intel and sold by Intel or 
// its authorized distributors. Please refer to the applicable
// agreement for further details. Intel products and services
// are protected under numerous U.S. and foreign patents, 
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 18.1std.1
// ALTERA_TIMESTAMP:Fri Apr 12 09:21:34 PDT 2019
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
OUSxmmhnRtFtFgx3OhLmaS7E5G4QMGmdeJ2l2OQyj95DkcsOLtGZk/ePpVFBBho5
dQs6CPxuh5JJ2pwzT3SsYpirwKFRXCLqgxjt8oAIS5Sd4CD7TiDkI+H5IRrcewhh
YWE4u6vogLjw1liDlUO5paSpFTn0DrHdDFR2OtQg4dQ=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 37488)
d+xgwad8uHMzuK49eCNaa+H05LMtJwfdmHUI8y4uj8jmLdXiM8hyXclyNGvWGKXm
2eoQFK2G7M9kyhEULgJN1ECGyvHWxMwIGu11KJGc6GdF5guruDQHe7QkqeGKtjTa
A4d0mikAP7OH19Ad+p1IR6qR+wd5Ca3+8P8dSxX5hgkVw3m7x3WaRq2mlRiA9gMe
cCVbp1Ubo3fDAqBXkUUx8kslcOfgh3VWRda/zkhPzp8AJ4pC+CdxnRAQURd9Vfst
oJIUIYWeb9jGyJICOzDJrL7HPzPFPfdJhOHxS8Efi2KKiYZDBRFXvQpsyo0dn2of
oM+LwjnZyirtYxhmkjI4RJ2qLtgJC8cq2ApMjPaIyqp6pkg9fizXDt7q+RoMbUB6
9qIeMMYTYBJUghhlHTxf3OcKzqvVL5HcL7h4bQLCpE10GPNGaIG9YlwMXkYk4FgR
YVsX+UY8SBe1v3PVEYzrPFTz1jnN7ivuxuEzzIFUsbZLwDusK4XnTa5PtB0ZcQVo
CnNmZw7rSV2uc7Zc1tQnmIjHdQyyIxQ2krV0ARD0GavkMHK263vbElwyxaut8AV2
tMGEaQBGNJs6s0dyp2wvIHPbnN8p8Jbs4CsBnT2ZLTMbog59Rg9LyWp+U9gn26ur
pBh6a739msbDCTgV6kWvC5dv4HWAkh9Q6zmDuRc61Mo1pNVXM6MaPtBCYEFR8N5b
23xrJ5ry1Wl47COPB+pYTq/cDZ+0DOHVUuYFxkjOyZoznQeZFMHEWWgC3Q7oKgJZ
vRNJkFnuZsO+86ZlzKuVE+mA9BBWPAlioM8q3sNKrXFWJCzeDG3VXQWcde+fCngB
hLRT/o8/S4+pHX70W3wevEAFWEy1u7d+nFaxceqkvMjA6GHz3nGC7KnOX6Fkugej
JlgmmmJq1kpANs+pYDbsJDnVjltsvHh1o+9Xkguzzy4bzWkpW4h0v0T1+oVuf79/
Q1iXi8TpLSFjzXue/ryv3Gruicq1WBcBFv3h3+JhCdaykmZpYbWFwoq7+ZGTvzzQ
3kIQ+jrsIX7nzsMs5CB/SIGTqhJz3m6WiEJ20YC/0wWicDagnyeJDVpO3OGfZgO3
wsMHUNyhvKZ8qyGRdbXHX1XGUXkoYngn1VZfO0tc67A+DLvQs6WET4DSuv16azls
5PsDxlHYvUG95Qz/F7f82vsFw7UuMtzgI+1HuDVe7MOcnPzqzMh/zX7HQbhnOnyR
TaGPNUKZ5lNRD12JP/aYY6cDJr57iXO7LYcT+eLFs+JNKJSuIXs9Y4WWG9wdo39F
7WbepiSoTzo6eRLpfZcFwsVOrRqzAzSGAsXhvK+prSuUMZd3If5rYkSWv2sBZXpl
IL6VhBgM6qCYq7xp/YH8/ubnxxOsBtz3ptWZjazwAR8jZcIzIH6AKDK9yjOWSn+q
TfD6zcm1JqWDd54AkKv/tLMAk0V9KRcxp5YWqJHG+ydTsAVjcyDwasXr61FpDKSA
EjdsfUVSCo5miLI5Q2tQ3KIrPjbuS8sRc7jr07w0YkbXfh8XGn4XDSfa+MoDp56Z
5sbIY1VwnKMvfnBI/vmb5JJuD80wYmeFeH6zYecY+EuHa16VXSkcXRK6vleflpWi
4HUIDxPGNoZy2508kJNaFqk3TMTJg2oaYHeLYpXyRbRvgORBVZ0xo4tkfkXGBc+X
OexqLPZ+0AgCLtk6ED6J82If9iC1mc51g+k8JBpF8+Ba+ljFv+ZrgZosIWj7m7C4
rwFsMtcxC8r+6G2otTQM/A4a1MsGkO6SPq1+EYqodzgPwoLHpVdkUmZjQXKWlVQB
1lFcpw1shGJx9Rp4d2jZWUBDLpMiEi/SbH0LWVdlb0lyWXbO3jThGUwq6TMe0k+T
hhTtHdsBD2IzZ/e5+qwVchQTaBxMyiYit7T70cbgfzladyV0GwNEqRYUtQzZCD52
/cE37sSsKwvnZXz77ii/9tnBhKwvOuQKLXVAr48wktquMP9mvCTD6O2qPehRok6d
ixt1OEb9wcdwdQ0ETEj8e/A7QAqXSllxj2mYONvKxPFtKENo6EdDi3EDOmwNO87Z
S50yf4kNMRdTVz8mna7atQzbVYBUIuDLEm4nkjLUHUOqwWnewS+LHCtS2LBYerct
z2a4OamzUqtYJTUTA4zOdUEJAhL6qHasfXTfeWpDjb6Cuy+SnPpjipJYmr4lbAXO
A6lO/AcE6gFiUJMkS01yFebOVPsilMbfGWPvsZ5oeEsAcvAOzWUik3g7QzABu8T2
Djw0az4UvqHN2gJ1DxGZUHo82TEc/1Z1dw1QxS73aNSArw2eHMK1zKE0ODR7DisP
IGLEXd7EPiSjmWHTnI59nayu+ri48qKiSbUscnXbXphkUvBq+33KKQv1b55AK29u
047MIN9W3ugR1AS1KmJie4WDdLeAYpsYHA7053fWliQGrQ1l8sCC4zZmvhgpOku8
ocdjIU/23p3N9yCTxG6tlUfuksx+bnZKyJ8RhHAO9zuHnOUAyMxUIr0ZGKI74J5B
mHxGLRB3AL1uH8PHU8Dra0iowPcHk669/zhoAeEygq+bx6xr0ESA76yUFTfsOu2m
lgXCCDgPEHmM0WQZ9VINpj7eSn4QV7l+NOdaWKUa1JHIdd8aZfONcNvKLJOWZXJt
MOwnDyXatcSKLYF9MQrYD97v4E4KL/M8VGgUfMhMMncpkJbJnCYftWX5+EsHFSMe
TJ8LbULc2jvgV7vYml2Ep1n3ZVi1QH1xbzcgesxomQOiH1C2lNnwyLmYnwR/d66q
BtzKo2yzeBW1qfsMc/SWspmm14RieANzUa984fNOzGbRdTPOWLEZh3XiOpAsVOZt
wnqE5I+RhnnVYISdb0DoeEiKFlLvO2HeSdMqh0Vhk2ueo9i493/luAECBQhwAV+5
1fvo8Girfu9CibpUe0vYI6KnTsg/p98hY14TNF0LXpR/n3QSNQUmLInmaTq0naYp
VPSY+m1uZH5Vt1IyE4E7kWoKsrrSMh6KblgEXb5+ddEFrf89krQWji7ED33GyCLH
wItHtKlj7/F2SVAHZnHY7UF7fZy5TRieMThkFbqdArFiRVzfHLpb78+lhT2DlbgX
py0vBmXCEGsJ22BZkVYMSu3Il2JhYty5AqJJweIqeJfoYGfVQu+ehyLL009JEfSL
HgmNboW9rP4wvLo9+IEbD2xHP8pdRwqguG1MNYW94Z/zv5h2vkNdnR5RVXyYm9QK
NfcHXRSSn0On7uixIyZ4TDCSZNWFpVcLS1e249wBDOJ4rUbq5gTZmESMR1uGXpcc
EjpFA60EFixecm5hjbBMjhudMmyevhTnmiPxC95Wk9n3YfYPANup78NfjyUpDLc/
K9ypDifoPFW72OjUzuiS0XeaOwjfqlIyNxKhKUupIAzlRZt4jDCLpdseR3gSHWBF
THH1U+S70wCnrW89VCbCcrgYD/dJDkyS5uABxnGD0wElh4fEMlDybwlBpCqAvSrX
B7rPCp2AS/zVaJFBMsc3ARCvI++U/7wCWQ0m21FG7UaZVTXu9Sz+KsOgU4OFLrBH
N1tNx3ClLZjQr2PwxyluwmRnssctFAW7zHqPfemb13iAEmnWaECbmHTI7W8417UD
80BQKlLgZGs6sheLwtxZAJuXRw8DZoBjfi/UWMDo8YgwMAvGuvPlvLZKmFXRoAsR
SswtNgBRP9cJNr4jvBSR1Eu0UNpbE1nkq8h2it+sJZN0QO99StXoDipAj07pU0wN
eM/fdtUB4lixsVaZvbYkCat3NN8+85XYo3ea1Qnv1jyIy4vIYYOgzFflgDWcag2N
/icfWF83JYLEPo16QOz5O20QET/QOdbUf4Ze71U2XOw6rPeYg2rO4JO510/KiNeJ
2V8F9Q+MD0maAMT14qSM5gLFPnAXSvCAhclyNNENoj3qHHWf+EFhj3MSmR3eN6mB
QbPHlra2lRS9r8VqFcLCWa1NV4+CwZaRo4eQ8rgGJNX0TLd2muoNN4Ce4l2juLvS
Q08/MHa1HOSnjlMlI+hy2MIVPVIU5Liiq5UJJw8HkXGH5zIMcLDlacji9BB1hyO+
roYu+vk0fb4VQf+aidQ9vrv/OTAjIiBIDqgkUFkJBos636tgv3VB231EoYer/t6b
icDCBv5lfOw+o/jWfpggyRUtNHD85JI8+Rvc409FokySAzvssrXW/16oafX3TDF3
XcIlzZjdHBcC3PeBKsDGvRZ4HG1vo6WDY54yYEvSOEGR8pnM5W7NBVBwdKZRkO+7
e7g3vK9+DEhPDJqCyATBPionRgZBbZ2NjHFPRLQub/1Zen0b83KmjigALApRl8Vc
fgIfhjcB8hhYPdfMxjs7hwQwJsqwjnyZi+kv3u2jr7Xe9FDYs1Y4LW/OVhPkRUSV
GrkJOLyNhgbzgxzSnm/c6dQOlxRU12BpdlEKsFJWkKkptiDEa09uzuh1Kcb5xXpm
yQowqPvwDBMbDimwwmhqEfJaq2QIJGzDrZkYtXrovApfMtxiks84H422bbipcXBh
DROY+48Ai+5kYKkxKmJmjuyAWkvFX8NVDcfwhkAAYEnO5LuRfSiCCEUk4mBEbyMF
trnqMz7Lx59LQqHciKyKFa3+tX4e7U2OfbwknSZ4+qwfbrioSh0X02f2LA61+rs8
uiAP1Cex4DS+y7z5bICwvsjqPt2siE1eGpt8jp3bOkZgPjlbWVWKAP3L+I2l3wlC
q1y22JfzJogeWjgokNtOLZC8WpNHYkPjtIT1ZvbXTdbTRvQZEpwLGvDyAT6APy/d
wX5lIogHhbCphrCB5thp7SxvY7IcJygn9+cHghBlQXMLFhZU999U6YpFEsvm7lMR
EDlcK956icq5my8ZwQ2pRD71sWJAm7uP8izS7jX4L/oYVmUXv9Qyh/6Ycpodc7Vi
R5JuLBMZ/TJ0aY4SjKMvixzQfx0nOUwT39IUFCzAkVhijejobnoJC7MxOCxFKLtN
N/JtpOpFOrh7LctBkG/FSSTknRKcrwwQlgFxUdEKQGQe4x9gRGvmMt1M/83QD7/X
RbCHMCsNkK65VGGB35NkAgEiHqnroDdUvC07pdZBnwIfpl2Cd2WmhDJwqeQh0ALb
dy+vVnyvQIAZkDpLY2QK/Qt1imw9bhwx3pdXGyDav2sRI+UJjK0vG/6t3Mv8JB5h
MaI5h851aPhGv+blvxVbcFNVQQFE67KW23LNPMCBSac/XxErJlSsTyzWw+flqabd
hqsd+/c2QDJvPOW+f09trlNZZ3Mk76Tf7OwG2/ZEg1V3g2m9huKFraYCbqW7xkDv
D7t5VjuoNMDEV4MrWe0El1mY2Zw5RotVKRF0guvJaxOF29ssaQZ/GIVgoVM0cAzo
BZnjoIsDROk3bXnNHPq1+F+4B4wmQbPIYlvsIFY+G9VuVq9/siwjkc8ekxdR9ZYZ
n53weQIvYzB5MGo4JBWGhIpNOZBDrH/WlxxhvC83Ea7jjQP+YRJbGBv15Gi2sl8P
SvgPAwlPA0tVzkzZT6If6X4hk8GRLON9qBCKF8ABIUJMwEV2u1tb26dN8HXNRAc0
YnAWB6Gqr189J7VO6IkGkSgWU3w7/U06GwdF70wflmNhdt3NgrFGX2j39m3Z09bD
sJg3pefzk0ljNtm5BPI4ze14+QkZ7jBd7y74q4/7MX9cthTzD5HB/mzPzJvzoJ6D
T/FdIKgksH7pwYIFsygE9OYZIYOb+VXLFXT0phI91HQk6Q5bmo06OCLSjEDs5bOF
a5BKoMf3+UUr9Y3Dfo9MZq4Z96S8g6dNJUmGSrrzEQ80dAm5j8q2NY+MRmkkm2dB
G8Q/HAjmhE7fGgVfcS7NfddgcSKLsEbas6ijC3vIxoWTWKBFLF61VXy5DBgQjY34
ybcsLj+6a3U+KW14CECrAo0kRO6LY5StMqATlhuhOb6diFDaluY1adVxWaJ8DAZ8
QQKDQWUTV0VtlPAplDjZtblaIykUIzhhfBM4Q09RKJ/Q6CF4ZB6pIC+xanCpvgvA
Qyg7piJfzQZ69LGgL9boju6HK+kHexrNPHYJOwFfYzn7tnoADNnEwHThxJyq3bIS
oawUTgNW4CI5SmhQIsppotn0yA8OVS17AdU2YSZ/qkGpcyC84cWF3crnhiq4I9WJ
fWTF2zwO6MCddNrb1N+J4Gz2cpiSsMRRfLOC/hKa7x9puUssJ/zVaVChVlxd3+ct
WsGX4QL+tdaB6SP2uHzYZhaCAAIts/GUn686WAO1hXd4r+nPfLipWewVseWHxi1O
i8R2ZFmVTyqZKpzhFcyWqdFUkZpr0BMiSrNRUiI3qqtJEh8N2E+g/zlR0hE26JtT
u1Xj2NRke147lV4c4UW36qcTA+5Uz+CqltSF7IJMUsaZiZuOgS3AwUjAXgH0Gq5Z
soTISfyEnhaYxSO3ZOkl4fJPXVpD3uJ+mDab40OI0QJQwYavaXybLy8NXc+eMnlv
YDTUUxEP2L6Dkaj1PlROvAgAUigiPT/5SnbvhMpB74as+Rqe6to08n3pxmnrFK3j
zL/uVXx13g/IvAGBoLmvxj+2dVRS0ABmHUvejohLAlZmm/yIoSveRUlPzSQOEUdT
xhLbueog60i6iB6opgvoemibTEP+xTey9EPwyi9vM8dO4XhDVgHBquGkzIFUOq73
SvOve9zOJy3LAswGEmEBYivp2+ZNNiNyvuoWya3ebJ2rhmcRAfzGEJOUUDFuXPiZ
KLFVuCoR+aDmdUxn43EWO0yT1A2rFUtm5eKjpVC8RBRnaLjMt6DYpgtqCVT6pJdj
3KLckdDiXaD9kX3UqF1ksUGWgHYZX0EdWRnWK9zmVybXMWrFGLvAwcxLyyib28Xx
K6raXZR5sDkSf59crWYT390c5z1kl3QImrlNN7XkYnjfB1tWryfXJMGSv+ZmOaOg
2gN1S3abTZ9k6A3IX61O63Vtqz+w0M76rSBwqY7fPKEjVL5rNH0Pv1w1RCu/0v8m
8edQDab0ymVZd3Dxdcm8SX1OQki5lTd9RmrQrALJMz1xl+LckWr5V5eewEuu2rCK
7U5dC2iI1Xkvf9Gj4GYcdAzecndCvUZUVFFVct2z0A1xIcGidhwNybVVntD+NrO5
S43vVflEMZu9fruLR0cOfrG1Oybn8jFShckSdVPwaRQY4SJ7QuS1VJ1zVTyCEER8
y7auYgUp45HxCfvsH4O31GqVlseAhbgRwfcdOc91sszojYB47+Hl4Y4vUykhq1gE
NegCTGJMw0J0hDMngA3cN+01RXDDkVkGhx3kC/maSYrEquQ3YDpsGlz3X46xXnmX
lPFYGpZLtOrz+XDCrzR66c8bLcvrc7CkJl79h6emnWxCbygIvIEj4uIk3Ws7pSAu
flymB5VfIMEVYCSENgBPA+6gUKVyhLs3poB5BlX/cKBoqyMJjntH1ZlOTco/FFcX
xuNfr9MWmGI6Fv9jMCfCBfW7rHDQoAnuCD7wMMaHDMh4Y7UaMn3LB2UcC31DXk0H
IMAGz1wIHjhqT+CSFQhTQ8ABRBUr4MTh5Uhiw6e4poBWZ6/ZFJPKxKDaiU8/Prt7
CAnqUYVMN0wtIpyuvV2VOLz1/+WsYxj6ttKsuxpIJhIcfXSL3IYDa9B28WygpuRf
ujihq6hJjbZbBqGuiedKB0kiEE7OXOgsTHxQr6v4hEfAqpHqSR039U1jdBXj+pVO
PQXYSUPmQLuykPtsfvNPqyc5rBQP95ZwTBuWI2U4CNOEvbP6Jl9VvF+XJNNUYyo2
+oF337mibgEP94p74uUU9VtbSEqTCGY3U8buu61vV1YTisN5Y7FCSE+o0kPoZQ+h
Koo7qG8NVlxlDf4vcUkJwsbG5b4Crkd4aoEB+fldxaNwDMh5qaEIeaVp4xgvL3yv
Wu/w7UgiRWZzFZhKHtgV7q5nZY6mD7y9VkTK8UvO6exUQHffhl0Z2gdn3AGwAqhq
YrfnqnvKFdpLKAP3r2OvvjFTjNOzy34mny/bnddWl/pfEdrgcxiXBbslvTDXYzHf
Taiga26NjjlAeiC2KFjBCfriJeEBQWTvn+l7BsrFBylogEsm4R2IZVKr1ivDHUHj
UDNevIpp1Yhq4GIATmKWLWA90cSiHWg+4IJOZef7E1HHbJCkZUq27QUszYXUI6II
huhwuU9XhYPbql8SucKjCdToWffAd36E7RjybG9CKJHe54ueR24fb06MefRqb0Z+
rPOATsRsN8rVALab6Hiv2sxCQhg6b2KYqf6dPw4TRAKugPnh9bSVq1Ro/g0ZSoyN
apcFWtW1HYw5W74KW73NfN1lfGde32oTEevZDDQXJpoMs8LfmNpe/sSwfOwtEpE2
k+cZt86fkDnDfces+xuWjL12N49nIrtufOhF+8CdP3hAHW3GWraDdSsttyUc+P0W
xR+OYSUa6tWF3+e19ql2QSjHdfq7cw+PfeWH/2qx/WKP5NrGfbCt2DrJ6eJ+g5bN
Y6EkorWKMRagEyCktbLtxInbQGHTuY4Rj8k5OPDgU0teE+YNRwKZpLO/KbcoTP3W
PY/BRZcEX1R6vEWPMi2PYRi8fFrXhOLImYuryg7drCB0kd/ipZMECXxoATfX/j09
mIWgjFfVDxDG/ytYJtoRKE1XhtBtkDdtYxOHUbe8BKGeXypQdq6cCt9jxmY1xhhO
C3/0NByVlSlt8KSMUvTny9MJbixyiTA8vRftyrhuCzpzK4lUHw1hg+PH9JV02ag3
0/gTJZ40HJtm0kQdQ2Js90QD0ReDuTpEgQsjHw0VFLTQosZP3BYEZCNs5aXRK+Lf
7eyeK+YzitMCxPYQ+5NOxR1JfXQTtypZ1G9+Jq+91xjBKjBlIPOla/kdWXGM9JI3
AHIrpDMjIgXyhVhmoLVo+D6gu3kqxaLeXyGtp+XTDVgijHndjZcb+7YCQGCJ0Py3
Jw60sKEujV6yEdAUoPal2wM4WtrovVswQWhmY6lAm5GhkQv5HtaAF9AIA2axs5/6
Vk2YbfEQ71emBd6uzTVndcbNxxo1OJ8H/rwjvuGs9KzdGCv//HyrLomUNbYb2v2j
/Ah83T/1HOojv3HTxmWh4xjZLsuHqroK2fpn6ZUtzaAOHC0Ltp24y0rdz1V1Tb7u
qyhoFSht9tzxqtgsEHtoqF/2rA75A9aMKGMTGO3tQKHWkM5AJRT+emU10lHXLyy1
frtckpzr71on94aZJC3gC03OPOsHfrEiJtQUAguACmCUUipRFi5O59vIb2xGKonf
9bvFWek1H/WIqPGtPYn7G/Bv88lhKjjyCT6JIot/dloeTXXvrmFSuKdRDYvTjs3q
Oy+hAWicG2cZupDUYXfgpVXQ92doOubUwX18sFUNf139calDcMWgCpvuSI957RSU
A9deYtb9XS4hOVGftavVtHH9zlKtL1BIBa9BLHzqfb1AtHLSa9xZHVAnG+rLXwwB
7z5IWQikBxrn4Xf/acHGoPUggA3P7Cc7lWd9pcAURXsd1jr6QAVvcpLNih0v867V
5CjmF1uJ2FZGz8/mp5WotTCn7ghbrMXn4doDmat7TGdc8nPZ0/QgCvbGODfWC4gj
uCDlf9pQ7KpPmUFEaI14NQx+FoycLlCNsu8NlETLI3h9P4+nWGc2ms4CHVLK6RxA
bmL6jOzW69+eqUcBst4UFrr/rIOqVcDWH+c3u5/18c9aIlhpHGREDtaRN+XBUUr1
L2r7z3xu5DbKgua9Vg0h952ObyxrK0hi8ZoSNskxmZMBUXTaSJUPaKbZD8FeQppq
Hx9wOH1YchIwLSN0mzck2OfREXIwL79kADZbRED2byN0FjP4v+tWO1PaR01mAvUZ
RaXpPtpz6kQBYagJX35X4Ub2a1NpmlUxaRojd1YHrckOV5HS5/Wd15WMKDjO+xdu
8VRHcsPyK11gFR0DTquIUOjy+TWbQfLyOkZCKPcEE8M3GPIasR1E2GfDvm7AJ2HT
wm5dVvHk4VHdIXAkONpR86xQTIULtSxCPg5Szg3QMloQN70CXFsyzrJ38AzP+Hwg
445MLfdt6BF68ydb4qX7yVkKeypHpy9aHS1WHzfLCZElUhsSmoWtXAmGVkj0kvmg
oGOPobzbmcA8oo9LvuqInu1WCz6XS5s0LKppy/pt8GledoX4Y0xf40VBCRhhqvA0
JtOvz2E06wC1t65xc1cq2veeA+Pb8wS+WpFv732CswCMXyH4qmAcVSGfY1A/NEid
kVSPZnUJd2CfohEqLQHtK/ITrcfoURzHAv128AKU68gs3xYgN/wGRMqpteXqM0p1
Z3TaNWhl0Vdwu+znZ1xa8ItWk3lQHYEnGVfDDkalYZGm0GZTfYnjw/cK7FwLG4wv
4G2aNuebKnPKBFVnNpsAbOwkGFsm6C38F1MiHoELb3wWOfLgG8yCoQH3mBnLUMKT
HzHfjpEo8vyphb52rfnUa6wzI3a0etsn8/Qi4Xlm6ODN/3QLAGFGVFDdgr486az8
y9Xz3XGkOUK4boOAC3Cc1RTVTv2g/DH+P5SOIY2GTEnJjeNZNuFOvsOrQnmBO0yl
hVMZcVs7kW0onIsUXLrfrgBWAEZkT8+zZNe9XXgIjdJkPbbpkU/S/mJjpgUjY25Y
zxRtoz44z0gSDUm226J+PaVLz3FC4SdiUg+QHxWpEHX36g4GXdmWivUEAW2oCNKl
1dmFg1pONBqQbC6X7hoCkkz2SdKuLa+h72lPYphBf/BNdiJxwBBHUH3F1y0H/J57
0ndvtSgoiPLMUOq/uESBXREknVXSICZJiW1MR6DAnhPn4AGl2t/vLkYdPqTqYl7a
g5Bf4J5bH0SA9yFsr0NP/jaR64gOTz5RiyQHIgC8m5uGOQsQJJyktRupHyBgFAyw
h0FMrZAK8sAUs2Q7Fd6hc9g8xttYpkUMUUIDqCK/XPQtmDqM9AGyvCEA/UzqeJGg
FxE6+8WzPPMD+Q42S/EI4TZF21beYaBqGUZ0tUyvftM51/iUvQZVQygvTzSxxXry
rn9jOBlXbImjmSU6isyACLxv04gAxYT1UCQE7BweJ+iq26TasNatGW1aOMXuX2Gc
hiPdFmTAdOJxADPkrE+PEktl3meDvgCHxnUHuVGi2OtHenbudGtDRjSM5i75cwaF
tpnTSb/APlam89KhagksWMZLm4tlbsf04XYASP+8VPAnjnomptq0lM5Y7xnguVyS
Q9ymw3Vpfdxy6LyLxvfNqHTgzC62gYEpDzsnNVunuR4rtxKkPzacT1EQDmC1ZBcm
7uCxE22EagmnAMnPkGfWaaHeGjd+VDbYjSrWyrXdSaLOGlUkOtKj0SnRLItnfsnF
7k2QNHiV8UQoUY8vz6xIR1JbceI4F6fjmTy5Q/77HkRG+KW/jTxLZ6jgfZsekwHm
s3jZ7zDo11xT+HoFjVW7k63cv4JMQR+q8yPeyUAk6557xXjnWM2qYKVNVYr9SArl
FnSgiNqbVLqIFUCzo2dNqSDyXuAKO7qTTTEQTVrKyT9VHgVLjvJML/tX4BzkqiI2
9RmS1aI8819odltxe/j95MFBpJmZYvich79GfMg1Zz038pw88dvJZCQNIlrGwAUi
dIo0eU3/WkZtUWdo9guORZ2LaFYGqyd0VN0X4alUhjJ0samDohcpRLiMG7c+JYAA
fMIBrQGCV+dlWKfw36BJppyUpn29Qo+Sw2NpExdJX6epA+UO0AgSgLfQ5hwYxcxA
aKSpHTq/XXGNLGuRBzRzrWwhg3cpZC+jbd4/y2RbgCvGqWFmeNVqZfDbKhiIvOOu
2e+hRYZ6/p0SgRWp0YdlWjyY8RRMY3XNJaNeauXyBabAlMTndNyDsTOKZjZgkbhw
iY7WB5MvlwhwtBRbW9s8t1/Vb7wzsssGWw0zFAOp1XpDXdAnoZuSkfWvXBFQE4iO
i/PMd2KVi+O/UCAG6eHq1B5ubmxe09GpAQpkciqeCwtqu1/aODVBkh87onI235EL
PR4sFvfDMf7AVCt4PgRmk6zBGbGb0Z3vMFJZesar30Kd9pBf/qhyDOdLI6zqxCrH
wgSlWDQTqJyJI2cqEhO/zUYHoHqzctjVaCBrDtap2ehhaoIYOkImwA+nJkhJ9umF
ae3wM4UVFFtJ96eYhJoVLmmovSxvhfZM0dXCWdJoYSlLC5fnjTOIeEb1ENyR2Ynd
E49NbMuP9rOQNoqBzzMMPP7am6uLLS4eLpPGumvB3igjs+iDvkX8EweImo0fK7j7
wfteTxMgLe0IlhCedFkTYIsvBcD9AoqSqDbB7eu3jp6WBeiJnqStvecNNrLdU72f
MkzKPSUP6ZOXbjDzPmMpLiOQPQ8RG+SgiH0CrjDA1dGWvM/0SXcKqoMGRJjtrl34
c100ttWtaYjxohDXGYPghz2GBozts6IgflTK/jKa4osaVVvqBBlfs9JlOO6q2EsT
IZy9ZETB2EcNDQLpREjgkZqq5W8lWoUlcA/MlvZTE45rSesKVBmcgtleCL84TcUQ
3/Y0FCgnBuZHRK2kEayJUMbeGS2jzH2RJDkNZ9XRtOi7SsIk8d1Q/UvnKE8Srgbi
yrwcLh8EGQ1YIYzP6maT/cbnL9v9AoWNMIXL5kEsIExF1XWU16Tx9xqeJw1nYWOV
II7ORqq5YstKXKsLBbf2U/2iYj1yuW+JmQ06eJ2eLr0hEwU/RfcS/OsM9/RloCVa
F8Qn471/gPfryPP034mT8aTjhnNVeJWA5mzpj4rVEYKoQPKqqWiOf0coFeBa6LD3
8h3+wL3n7pCHOlHZIA4ksV4nv2SzqoRA2HmmH3OEGQGgsxtopaxlGk6iBMlD5e3l
X66rrxvQCw0XFDqC+LqSRACx0ppSVcCY7Qfg5j6Z9E2/1I8UM7hpEhOgo20eDi4H
piVBJs8f8jRyzo1fdQDQHkbnDMWodDycNClHk8d2ay2LzUvGkCd2+GyhsGVqzLqv
+MgmxXypjPLSM0vY2xq2z7GDnBMAj6dw0Ls+VjZ5yYCU16ZyOXBF+Sy1kt3R3rDw
rmS/aRfB/fcvHsjyImUXWXSGA4VCZSnSGdAKKGiqbnd0sZwNDsujtgCwwV91ZSze
eL242JoEEgLyswFQ5Ety3bdK0kdNzRP/gE6NbHOzxUsmTAQkK11GxilN+nuR4y0Q
eT8vUwgLeOiJ1AmGgGiZN5DV9z9WQBOTgkT+laTDXcQW2UjdM0EpftLcnrQWSnAz
Z9LPyD4tfuVZZXbanGwK1+jdZS7v9forzpM1JHNfizpyHP+UkdqhkUevpZDbNd5U
rRjmlhEjBSOxIC7DOi5O1X5V+Waej5NjkxCo+6yKitIrYTdCZmfYkMWI+BARrbnc
FAP81eUCmXfsNk2+NlZX+4GHM6m7AMdl5sXJcONIVed0IdsLpFlo1nqLDqqt6oSD
L3U6Wb+HGvnrSPVaJ5++lSXgT7LYGdYqTAUY9jd7b0kLBeMph2/3YAZMWofI2NDB
d1bgtjA5S+enXdtwvSeP0uVT7RVksx3+FXcmaH+HPyuz4INMq+3b/M/dRBWTAStw
ISsW7cNjqvXXDStHSlGMncrdEVD1c8DncxZyb9hzPVKl7CqefvWn5Jt3//wXU4A8
d+rYVDVW5tc0q+8Bujho3FH0IXLp0i1WvIl/gqgW+sEIz0cr7pHlnq+pWp9N4ASs
hnmfTsVzrsYY8F+ZR9QGACNT5UFCd9oY+/0kbyQ75rSuO4kATImNI1jgw74nlh79
XZ85pt/EpS7Ua5yl4kvHt778VP08UlrDlxC/YvHJs2MkjcYZnX+SEn6ZMWZ++bzt
7KLeHdUBAi1UR1Xh61b/cAswNaeLMpJT10g9ocuDfPmL/nCkwZtUjpYroC+BN1XK
ZK6QfV3dYWzqCdw+nP277MgCUA9PD7uO4pSsbHYrxlRt2eazG4GIGpteRUj2uTo/
QYnk2JfNBB4pWB2j4L8InYam043RJxkzZxny5h+/cmIe4jVf9TNNBA7J43HQrAnB
5svCVCuy8p7HCLWiS8l3iVERbZs38K1ZAJnN0C4fQ5h66ZyGIcwz7MjnSMbIYaTe
DBtmOjagQQh1ZqxM9cA6YPkfVI8cOy5kjr+/5r7bh1Sk21UaIkSgkFReFVgmtyow
X/Y2SHthhxBos8tzkd91Ct2ssRybv7HnNDRqEXQllBUqKbIt/DpYNW1mk0kyFyhZ
QcuEVgGf+buhs8bbHaIpdm8R3guRF5msV154kaLmWpq8+pvX4QLE33wXxFVth+V1
Z3MG22UE5eWbz7DrJMsKd0h2DqSBtdVlrbppen2wiYxEXl+JEtbTyO9ZdMHuyLE3
HBODAVfv61XqV89sc+rgsu9taBhRkZLPs5nSpUqcj5AKeRzC4JS9C4J4AIQzSOmg
LYucbKiqihkhPvib8O5I8FVXB0dLkZqRhe+uOh1VBQKy5g5pxfVwWZQULM89c6Ix
vPgJJfkA9uwB6KxqC9zdN2T2tpjiVZSW5y3OvOLaMGp/GT+vPTBEWKoiXZMOB+Xg
qfEDUMuTuOGx0YBXWL1c4xlJNYth/KbLHZ8Lp22TkyhwqcilJEblDjx8MseIG4mW
yXt1nrEsHRPREM+ypDNSAkpLiP7yzs/GrTiSOH8u8eSnlT1N4yQnNZ10HbNY2nTn
MAc2gdRguG7JoQUqGVkYUVXGPg3oDsiRcIoTpdd4E9IGP83P0tGSwigCScHcFnL4
kRzdL3R8XnH32qVTUkLVsD4V43om1kTBUbTqhWCo238UwXUKnMArD24gFku1sAgo
VMi0NFnKmD6MftvouGYkZ9Ne2zyzRiVpsiVnb53cN/rG6K5o4k5Qn94IwCHFldBf
0a9TTShOlRhXTc4LwSuQ60iLEzKxZ0jIx/xumZmoQnEMuhp7hfUHRKfNWM3JDSZ4
4nHU4aZkR3J/0aYyjimvMBxpALza/wA4uOyTv0QZvTAR+YJOzX9q5AkelPniiR+I
l9k6nY+Vp7lc25PKHDZrSfYjXocpn3CB+THeBRYSoGYXrUnWzsPLwicVMgFrl50y
9Uo3xDc7u3kA28Itcz0h5Jb5oENkMRYTF08VoVaSDsFqYxXcj0R3+PpLN4QbPTqx
+g1vGLaM+ArPgzS9cNPlmpzYf5uY8IYFt+gAEtoDuv1y2PvwZQ55IrP+yWuGOt0I
iklOB6wo5c3IYIyKoE6+aswvZr30Q/Yxb+x/+xdUM84HyjaTIWhOcaq6pKkTojPh
rG8ssblAh/hq77CxdAGUpxDZNKWxKkd6508Unk9mlQtechb1g42DqpH1ih2miw/U
30osk/Siv/jcPvoS1MjFZycT6PCym9jpVnK3XF7HUopWJMm8ugtolaOh5nfNdk9H
4cg7+lnHID5CGWeCPPCL7TQK97HvqBcRJTUo9Ulbdyv1MncsUSMvZ6GhcUIhkIto
pJ1Jmt5uTSPgpFO051/S9nRa1vLRBv10KGBZTw4GmbTYVEecvTRGMJUoIOG3Sa7w
1/6hh0D8itS4PGjUUpTABCCO9GseZ+dzt35jmA0Pec9HdhQKGI78CeHb71i7LK9y
CfpY0aFpm2qTWnk33ojPVbTa3TcoI24rv/cly94um/mgOJZ33vHRRSN66qOVzjYc
EkINSNMy7nLUm0ulSjKU4aNqhwFJuK+VRtqGHADJgfnNn2I8CBP5aPUVIMNR1hgI
ythJcQKskwJRGsybIwwg69F7UhDVWw0PoZdsRGDHUdFAjZEsUQ0aAbvRJZ1Sz8S6
aikhPuRUR5vbSiFcPTYe/QloV1BEXrjyYoFmKQmIQ6PVYeN8p44T/AldI72UZyuo
X6UZeSAop1dPM0qb8QRb3Tf5UpZu0QbUtpbOw+9ylYOijnH3V0LQRZ58kraIJ5T9
vyaPv4gkARlrX8wdMegCqGZ4kgnvK8k+ziu82FrdeAooqvvPZoUVCJODis09tMW1
ZFwnYGuwHP0K9ilg54vwbn0w3WWtZlYLYGR871VMXFogH43dtSSGqop4i8PFPZUx
vgo3Pvg+xxfmEBu5zuoykHd4Q/h2Q7Sk18xulYmuorV0ZXbVaMOTKEj4MhCaGPHX
6lRMcV70/4x8bU43UACUi3vxNenkg0k4BvQgwg9fhW6tLRcn4evTVtwpw8LqSiGm
PXDl42oQGjq0Z0gh0PABaheOIcDf8f6J/wU2b3RILPlOWPp163x9aVPm/E9mOKT4
QZnsLlF3B92gbaWnKLhwWwHb50mu6ppS4kt9Jq+ETxM5EzD/cQ9cHCm3utmz6YUS
afo+frG+zn5YfC1fVILbzUSzvN92woC0g+enUSCQUGEGigE73eV4BkpFjuj3VJYR
T2Kr4HkEY884gBfLRAt8cB3O3LNtve5kAnR+ORhpgyKduH4UJzGxyhkmTsr3b5Y5
SbwXlbllD8Q2BYozKacO5KEYR3Pxvaj3RPI1QwVKWIp8ZxFT83Vpwdf0BZU4rW1O
UEZEMTakFfPeexSkTGAYdTiWoevxa78awVu8bPMTQ7DDqhfrMKatAWtSkZ5G6sAr
gsuvtoIKjNqLT5z00HQqc9LqK1Z/zdp2HnpiEaH6Tm2oK3AE6bEtNI3vxi37Yb/8
+W8/S05RceRn6sMW/KY3lfqelqAh/vPFCa/gPyteVD2GIkcr53prK8a74+R+XyMu
8JMXFUwXVvMneQ/PWAkG+iDdKny/yvXhe/f3SalbZb4QVoQ0RsPUziHrZuePmocd
6St3cXPsAsXqBv04lXx36NykjkcKzR3srcTMpAZ2j3wx/vrKU472VR9vCesExkI4
rpkUy7F69SEZLk7oTk2jRbPOGMZw49bhxqTQH/IwkJJO6px/jGrkQWkdzyMPSPOq
DpuHYa9c4RpExnp/onXqs8Z/9KkUF5z52zq196otSxA3ID1ONT1wmdJbCjBNf2w2
Cg9Q4C7MAP8gEPxiHFxdYX6LQBUkdiZv7JptSGGMGbSbYtc96Q0U/dKzp7T47oJ2
e8S//p37vQM5ZyLYhx1GN8j9kZnkP7SKWBCdNh2iPAGmIMrxWVlUYrCXflbWbBrJ
PSwKl8Sp4kRAUINUumoXnEu2Y1y4Nxs7iO67OAozRbn4eAmPjUgYf5V/ZDvU2sfI
Xm/usk+IBjiEGsK581GS52wr2mb/2pixh2TEpELHxPaF1KPNz1OqQSzfdH6rRBTH
ljzuQtXeSweSSTJgBMsG71P182lNRo212s9KcDBNdiWZDFawH8ijapz18gi4oT5j
uOPUiut0uwSzJ4iN6vPb6yRm3Hv2PTEPfkWNncqESLqBF7ykTvNqjO1l37tBnBpU
vBter67k0Bg2clBFyMLV28zJQ6FK6NPpZglZQDCVm3pukndLBNPhymqbpqOOd2ZB
OrFNzJBxU7cpUYOfIZo+xINa+DnNcSz/XOFODNM6UH2aazCdPiKbVZo5ri9fsWvW
QwO+Xg+2mtXh6FoyckQfnt8fOjxxBr0PVTs5wAOISbS+sCTJqkv/o+g3pkzSF82J
Ek4437TM4930G25VCMrDylEB7dJ7V6E3VUmUMv7+bPKYd9Lo2qiPsm2P9p1ZP9zc
ulM7vwJZLEiCZMr0hva19BTc+7x6NWFqxOd3DhvBmFSgJNuz3cpCyKgvgzA5laE0
JRomIbrdt1oFN4DIPjfVMJ4ghxs1sMlaq+5+4WYg3s4QO6NQdf0RDmg7PqIjdDh+
pOgR0qmkRsud5AfXOumPML9u7K1UC+MtoOFt2js0pXLvne9jInvOq7J01krYcX9K
hQDirPNa9sYZsVv2/XhIuxwIGJqhXffrIjsLDlp8CDfCSSKynpl8yrYthpGM4sap
pVYCrJJJz+MOHgu5XGW0KanW5+pqXN7nSa4Y3GX4kUiU4v/Q7mGlhb5UvFMWQE2o
P8QJ33pDLitHUWq3NZeHOhCa5K9yWWcgn+NHphOT8IGEvBYFyoyyW0yYGtWN4uoh
dP8h/JjtLa0gR8q2YVwd/O/bZNbbwRo43jwyWjrZz7gQldMNBHn+MIWPKKJsW+IG
itAz89Incf34Krtp4c3rCoZ8JZwqy2Y6JeS+11YudoHDb/Ov2zNlBGAYeusTsNhz
nZjESTtw/6g/s4tBn2X4ZDNdtSVkFN8riKG6sefXrSKaonoYZVOCvBGSuSN1Q+ed
jJFL45gNOljHugW0cH/9c6iaOqUA4OF3gsrAGc/ngib37UDeFvkVChtEMDvVGvKi
JMIZ6bz3ykvjq+VvvEOKIv29S1Xm9owzXW3+SbmuLOL8nEVArDKSwSO5B3BblSY2
tb7D3XXisk0D8w3gJ/x7Bk4fRrLYBF7GEgbh3lXoUVhrr0H21rwrkhfTPr8jvAB3
aVs0+zhBl+MxcoHPWII+cUjzAsXVx+hUTbcA4hHGmyAzaro+4Bv8pEjBnltydtqw
z4t4kuvy5//4hY9ATer3mowqlj2VW/7Ja2Z8EQyGLaF8YoowqVNL7uQCzNuNwyMY
ehg8AhQOA3ixC9PB4RTjMTERlbw7xBm7ZUHa/7hBlgxkTYkNTmfgDZk6v3cqw/UR
X4UKN85pASFu3lS4KPEDQaFZYwhRpeFLflYOssrFjtFQwA1gt7GdzGhuGWoyGgAM
hRqacrIaDNZWzrHfTtkNWOU3tBUgRd1uWgh0fZhQY7HbQP1FZQ4uVBweJQMIYxtr
dr20ZgnQZD6UpDziMttgroILliXwJUg7wYaXFnZ0adrF0dUGMlGlZlqLdJOz54Ga
GLo1OZ1QXnN2WcuhBO3ZXDybOa9tlTdPF4Cos1DEDmcWwzD3ecLyLgRssRaNIfIs
gC51HcmpGVK99Z+CLcqGhb/mkBn+I0oq5KaQ78D+DFYeou+GceG3IrDQrp+bIhtD
Qu2Z4E12piQ/w7ULnY6CIuI8JvYt8HI3k4pCpTjGG7ujUyDElBgsXAHhhrebJtvY
diRQQ0vgwlr2rldhxZQ4BfHONOl7ojftsQGLcfpQtFnbP/Tm0IKyFFjNwCJssGw5
j9/FkAX6hu3IU+Pmjnex3UD71wnUi7WlEl4jcxpR8xbR627eY5DG7a5ufrenFcX3
BFJ8eYH369zX1IJqRLju/c8L77dLPOalKu75y6v+TAhZcf06PIPvfsaKZwh1mtfU
LW0nvbha7wxU8Ppk0M1m3lTJU0ZkUVTWkXJkJ5VI/CrL2FT//kaFx9GwfHF1uYrj
Nt4RcBJW3Rvv/wuRpu/j6ZMj7KbCsVPcmpug80RkeMa/9FqnBeEssnZf6jJNj8Qi
Sxv9Y6mUrsCRdxxNxN4gO9GgquUk14K2dJQSFMFL42R5cZn+oiAoK5G3N6wzwwxW
RDiUqKHTozwICYBX3BMSq740pWZo5Dl8aqSuzp6Qc1/fjK2Z2RtKKxLRxp9pjIdJ
JzzQmgi6RFltidQ6zvTWBH2wzYprm+/qBjv309wB6iwT/pY+NXJeVA0qHo2YP2L6
KZewCFpSs1Pje31Qes71gqGQ8FZSBPub+KNy5Fb89P5yBVxaoJ88fREi4++iVi9l
9pS1ps0kenqtriANu0Y7aq0bGkPt0Ol/NvSoCMo/2RIvXYYi/hwv4N2qw4CwY50X
PUNWMfpe8CQegkEmknG94iLTp7z85OhV1j+9MGLuxks1yO1yO42Noi8xZpXxgNbe
NpDkTtOCO+HJqNB/4CaKQzgzE/ZZPa2ba7jhODDEL9QnF5t1vU3GsT9McQECG+Ky
LzOMcsXrG0lD7iep43pQvJVkioEMdb1UgxjAXulUp/siJHorJ0mLMfFKC8QKGgT6
8e3Faq20NdWeeJu+4PSzru7qXzsdOGj3o25sWhpXBtk5TwxmrwfCqREXJP3+Tkhn
ekop1cWDdH96AlC0dP1dgRcE1Ghs5NWmWqQqzEkusfRtchWwhtLY5TohSgEEY/v6
6Z0epk0B/7WYLCMzzCy7Fe2ZPGTqgqgIC/WSckHYn9vn90jEfl5ddxmpnQYLwgKT
way3aFoGuW/jtK401Rrw5SXqNC4/Y7e0XZmIOzNpEILkwhQ+EaEQa76atsJfKIC0
76h+/eAEJdsOWEQZbHqAOXj4KQU8+vhqaegGasHuDPfDkOxEoaME+ym7aD3NQbm2
x2urSLW5GRMNRBcOQClNZ+stIUYNybFwCnDU2y8GaLspn8Cgjgt0ZvN13Ei7YGju
E1svSUzcigyRQ81pC0dEKKOW6gROZiLOrY9o0g8FV5RagIE665/zaTjozKZPy+PU
UQOq9Yt6vmFFhS4BplYQQKDUTtNU0MpylzkzRvBiBSQnZpTDrPdXK+N3lQTZ3o18
vdsPOJiJLZXn4HnChi0xDsT3fTtBdYoqXcqGinXJwfYJMDaBPeYUUpjGB7nJF2EY
2FLKBHBleWdxUSIbwKlrUmO+aoPg7NIgJBwF/b3Mx2ddDLb4kZY4/HXqBBR17Oo7
FzDawBuvLRj5xPGQpPK2Vpx/GqkIrp5meHQeui5df4qVutpqkWAdAkJJ2tn2Yl1S
5SpUuuqVcjGU1ngTUejf+cTczCzjUIvvtAGI4G98bH5noqZpjuaI6sJUuaTMzoN9
dxnNTEJHinC473NJ6SYbv55jjsANp3rlglPyMmFiRXkdHonBGZ8ixtxK1jcw8vON
RebnSptJ+h/9o/6SZwME+YjLPMOigJtuvgofkBdX1umDOe13NU1qDqFr8TwpZzxR
UapMiUvEpv+GpCxIIRuYKJh5F8W7+cX+ib51BoCW5mcS8XuZXawMmZ3gFjaowXJt
kwXylySl8hljVet4Dp0bHCUWhejE+r9tzEA/36lRZSKuvSV3F8pRF+GMsZzRKeZK
nlREJAQujJ9HWGRuMWDVc/tWG7L4/K1mj3WUFiKUHzn6MJ0DLHae6suMMnTJH0et
uv9O9ZfaHyOWV8Owa7ADeNRtvlvGv0jNi0gZVdHgndHV2p7nO2mCqEi5XXaprbY6
8OHhyOCxx4xFEmO4LSkPIGvuEbK4UkPWvJf0A9VB9ZXgogH7ISIt4ddO9NoDMUTE
RWYCHj3HtiRoiiyAri6nlJKzze+gAjcUQeeP4n4juMAB/EClRjZhREd/G9naw+zs
1O+xdpL2rSyGwhDIsoWt7MZry66r1DC8E9SbWXxZRCmqqp2ZtvqDfz3vfh0tVyWX
GrGTRleuhk+Nw1akbCmXld9VVHFi1LCx/mg/K+cDHyK/O/McgE7/eQyDTPz/TUHu
Q4Z9FnmDMocX0KE6D1heGoGyoRno8cRuHRgn+7pEaBmaJFwF+cL9ulHv5qF4vIKm
RPkIpHaohUNynWIO/M8ncxSmiIJPVZ9NuPxjj3cPL2QRWUMfZAns7Ly7h0e+FcAh
sD0waowmHSl+n0fjMMbMQ6bVJe+fHoT4RsQr6v2DwxQdNxEcD+0wAy32wFJGC4xx
w8M9u/kdeIMM1gNZoqNXRJtOpRUz4SOsNNAvBJ/y3apJtcMeQ5r9+NmQA0+AFdZ3
HdA6wCvCjLV+eoVvqz+i//GnEAcPGLjjBgvAcAWewWm36FHkrkgYvScAs/IHkpw7
7DH2Ynz5fgNRGA7nXM2cIhjZubz/cB8QIlMYMsJEwaHSv0XK01h9a/tVLxmTTInM
8yWTWyymLdGV0FN3e8vnZEZwW1pwV6DWxCTUf24ny39i15TPmRO8sO8Pj1w97t+6
j/xIsRJp1bohbIuOKxEPb/mQ5Wm+vSsJ88c6wLySgnvlIFMvEy0Uph/CopvS+d9x
Ix2b09ypb8EUWKyNKQhpD65Cll9YR21P6FxgAWB0LWveDvjdm1nMaq3I1XMF+P6C
QJ/rFGLCjELzCIRhcNIUSXwLmUqme9JRbRKbWh+dAMNEdDJZKBR60oGZ/aU+no56
TBpTgDpMGBgNbCQi9hDZXvK5Dd0GiVzL/oAZdn4OAFIV/SerkieswhjcuWA5YfZ+
wve69xRAlc3s/OPgYTBNJJrZlLkDGAfx0ZFD7EwOCRBdfaODV0GQLTHgkWxX6WDk
iTDkwVPyFIgVGMk4m/ddpSGUymSs0D4Y2VApIBu9XVXUqRxlMzB84l8SMKwTWK/O
V2qLzNNbe7hEG/8d+tv6/hMju1nfJK6KJJnrOQ7ytZy84R1V172THiPKaArcrM5K
QUATnWs4ZWQnnPVmYTXYxfrTtQ6XgQy5BPBgR0jCV9F2MIi2ybD9g9hiq0SrehHr
mZ9FfN23LJU99lJN+BEt/eUaEnd2FWh4+fxlnFaEEP0YMddNxRdb2CJF0MJ8bpHr
enV4V+t+D2VhZxCockVE1MA5PX6zI6nw3bq+e5i1WjPqIlPbPzNPJ59G6966BqBP
+wj0r6q/RVpTUGuELhP768dqcavjzx0rgOmQ/zhzeC3CxkKV+0txtWVYv+DOUFzL
8cBHl9WoTn5eT9GODmUbLEDXv8aCl4Qe4MbOHE9oF9Wuip6ike6OaMeMsY9hn+jk
7tia9Tbpi0AciRIKQU/Oi7HnKx9ONrk6Nfpi5FM0fT8UDGuZOPSsEjtl20ws0pSI
OekadkOBWnqum79wJ+LyMm1GcgubZmdIQiP9VGheJiL5RWNc7esc1nSDXSvN3Wg1
2sodtkrRa6E9PByx9dHHrbInSI7sK8kbfLysCtfYn/s2TvGrQqROKzI0+aqmrKl8
WnkZ44iGNqDL9yZTTWe2ovaYd0gCMKTGeC01PajXoCtQJumZvTMP+/vcpmJMJTwA
sIh5HQzhFGpi5LqfRpYUYM3lfVIVHqUnCpIu8MAxPWnuc0s2jQuU4QTeKd+oI5h5
yaqGSSrU/OAd8jQeR3S/n/qCgNA4vJvr8jl5IK6GYnByATNRDsx1sYbOvaMBNHZY
EFrtyga7zWocNFg8eJT1yq5+GhIG0zFxQpZFaJgTI+Y34qfxT9p5ju6GLMz2A3kR
dATMe5U1g2+U2B2Qkx3xYpp8mQqKT8r2QM1E/ASY3UaZx/Mc/7Tg4oLO3q1902l6
Rh2UCI+xbr97ZqiYvRz6IOimrxF3d0KJJ/7ibjC6vsupVKuw0RYMLCRp1c1KBWvq
s6irtHMPcNxjYjHv7UEu8BSDFE8LXwGUCVP8z9AR55OPWMkHuV3tA35J+hyJ/fBU
sDxE3eXeAZ54Xuhxw57bvQ+L+AfBxj2NmMPYaXwei6QsjaHtZM3SYhMMR2yMC1zk
era2WsD1GIuuKJ+VkM3eDlIZnZwRnLylTY6CH34w3Ki33CgNtqoKnCC4+VV0oH1E
CCHXvLPCyrkt+qdcQHMQzzp9Z0ZXl7lRYVeU3d1wTdkExARepigOMOeKDG0a/us2
N9iRVvtIU12rBvae4mSqPwAeDH/6kvC2nl44EfXrP72W12jMIIB0HhHmSsIcvVa7
AHGaIcqTJ6nba0bW6ZHq0d3/YkSd6w+TcYmnaojypX9pk0by6mF2ZXT19JSkJlGk
IC1MXGrIrIdvQKIv3IxKfNKPiHSvCs63GURYudh/rTrd5okYqmPhHYByKy5VFqMD
wRUS51VGNvjsBo+FZab1oevDiUZDSf/yhfwQ2Byasm9kBQjvHQ6nof8AXp+6oBQJ
P4SLQB4AVn39kMzq3TKHmscUUFcFlE+uJhQLzDH0sOHgExjLC6OTFB1ZM7f19Vex
kEzgUoTRBnpSKUJLBxGc6XePq0A3AtPAbuZY5jwoyPRf/wHbfo73Uc6/flxeakUU
kW2rdYVWrcLMpGVeqJm9BqU30Zi0oh7zbHysBcbQ1mR+g6CwR1tPs6xw6LJkCpm9
UpSnQJFfqvDmJZsVxEV3OITZvS2HbXvdi9l+xLBIfyshvRIgnVCat7KWiJ8B4J/A
nYICpN6yvyLnzZRZfBOrl/f0nDfYpEEM6v92q36EL1oPp0RVZPF7XaRheWGDTvBy
WAx2aN8jJ6EDbvSAXcWTYneD0Ud7KhdROivzOAbTKeD00zxHr8HnRwxL4DeR0/bi
Ylt/kIWb73ufeConDyWmkYi9zpkgvDNyPjOM4TtxJ3597lkhqv8orLYS5ePlN/ot
F0kq9r/aH6M5VI4JwFXUQcT6CUJA/KPjuScU9T3ZJEmfHEZmN70PmgvWXnarToIg
8BEpZzi8k80BHst6eP9zb44Wb6p//y2WnOgi75HwFmbwNTlt77rqnYIt8WEve4Ag
hYCRfzJcTmarLUVxrfy+WDfPH/G5lJ6QsNcuPZUE/1JpOoN5Yij8X3vH8W+/qjwl
sWE4RCQzWRaZDFjzJo69kSXpzBQtSqn8F1/wQmdOIVH/c4rrZNXnk4Tx79rbITUu
6IRNVCsWeZokw43kCJvnI68YFQJK0GMK5yL65RK8rGOGgM7GJsy+6SMWPpQYggex
xpPyGU3emGSgaLgdAp5jUkOs3nrO6WZe+aSYveGJOgxUN9ktxkLj/v/LgAPec36E
3lR7e1T7jaxbIHzTCo57YrS2Rr36a+LMyo30lr4leZIfowBn9pokdrD2P4scK4FD
ZuUMcMB0oCBycoTQY444fGFmiWBhM5o3fuMPvv2oIfwsrYZZx4e2kXG2oTktqS7j
4EbPk6n1eeBU0LZSO2gLnBbYmi97olHGO1etf+Gp3XbDzIAlHTSSiZ1OFipgzrAI
mTMDGTzxnmP4bRmbpl7sM6/HGdKXLIQ8rVSfdLulsxn2FKh4vrROmZT2mu+XY7eO
PIpdGmx2KGqH7DDMxeCLTYHvKPd3n2rnnMK3SACaDvjJuC/8cJmc4QV2ErrphI+A
Z01byt4DrfoxFupEX38fXHzjbee01MZj5cK8k9oJxYEVAhHHtyNqU+2Vcoj3YeCw
p00Xi1LJS+jo+HmjRyUNieO9FxK7RnOz/d+ZbeBDJk7Sjb9l3zTgoH5M3A+0Gvpe
Zfcw+VDcanoQ2BOBvMVvhgGmTz4/jD5RqLV+CxI2Vtc9VWpUdmrzM8qNzjpCItMs
bgfX0e9Q6L5uJZ+GF62fhVMpjHIxJy19xyVNbIYXVSTyYXYg5Rwk8JwvbWkW3DBK
w/9Rgxt2y3rD7fTW/8m9sfuIl2Ugg8lSgRk24rBikSV3+hhEtEJlujfl+KpmBBkn
QQA42QehAB4DetZQYSl+tzLZNt+oWCyOVH7YwV5cSmETwgxuZsNvJ7MPxuQg9NUt
Ysg0dvnY7DKkBtBwEKWad49A001oNiZzeJvJwF7UC04TN5B0cYcjhM7Iv5F1lbZY
V8kZ+LH+77aEoOGPsgzCJjhnbFTGLmqhyexvqk6iYASh7MejwOzh7j2tmbCMxpiZ
rDgZdJK/1PjxUKEFca0X23q/gsmo5Simc0bJmBkWgFixgAsU9C53yqnJEKpdE7Qp
ThuuVIFyYABYiycNvCRLD2vvevJ7BKK8lGR55bFn9es1oC7Nd8yz95ZBZ4aVRc25
5ssgyG7QyPym6kO4OCdzegPY+0aAsB0Gm4oZSMDxUZ+edMHAeDR8dUfAzVUtu8//
rOUY/qrglbYKruFkd+vFQ6vjFaC6w4Zf25316JbU1Ysr8nAjwceXhUpLX12rbkki
x3ynvECBGJSmtQ9Gah9k6C9lfXLWwkVIw7qclSHzQo+iry2Lox9VCIXDK5vRphYD
Wv6tK4NnlPC1qdKx2QcqQsPg+DYgrlzcpElGmrFD89TQPyzdwm9hihqs2RWQrh6l
XTtqOEOVhtMM6mx18MhozWUV41TAhqEZAU2Fw0TCWbHKXAtTBvWYqkfA66vVM0rS
GdhGH05rMwQG7XlS3oPOBINJAAn+bAkNtWpkdITSO9Rp2q+w0BHaZoeLtzXDcsup
lc8XP+RqP1XHCvT1Yk4y/KxGqa+FAqgLKg1G86/d1EEafWKDZmc2sOHyVQyFJgqN
VtVcF/+NNp2GWsyYWPCE8+uBG/L4S9+lVJ7JDlkEeHZtxclYT1T5qtIpyfbt1xzq
LbfELpIb8XFt+QW3M1mGlk2chFeO+lrhnDvlcPpgLmAGvjwC2MPaYXsVJc8Rg3sU
UjSckSAMBBmFCuRGZLfJKwyoyC0fNEbpj9oQROWmKmVtJiGU37cSHwbeOJ5qpbUb
Rs33n5s5zqGN+jtz82SvLlvvi/+brhV0Hw1eJukMTW1tflVSrbaYD1hwHpQlIBMV
ZSxQ6Dln9y1pxLiN6aB7G+Gd5xDGg3/eQsxYAYsMDuV0ht+3v3FB9UsStm+eZmow
wh9NQEmnMydArgmzDGr2oS684Ab/DyvjxMWFfrECb7w8fPkZkXprP+gWXDkSVYk5
asEsnt2CaLSL0X997GhgtZmVUPi7E8PShzMV2QPIXDgsL15C/u9uLn4fxK/gjB6f
R8J+y6M/lke6sBZsVhekIrQaHq1x7ktUAVEefcCLnLsrKcHBh9RtkBg2M0/fjTfF
1UP1P5JICpFzYSNLdZhZQ7zNWMMSoAWAUShId0tZ0RYa1XjPjmaHmJbZOQOPQUdb
FnMW6WJPbfcJk3zNZn+1Vnd2d2KiTK2WFvvJtqr/y+0UbDyve5uH0HJGSdmnxiVU
oFmNVDBP83xkzwiEe+49zPvEuwwJNGJCVylowk8RPA9W3zHNK749Mb6iHdfbHqgJ
4uufFM0QWGxDIg7BIbmbjfGKrewLH3ecsBaBUliaqT5OMj+zPwk0la+xi3p3fgS1
pZ1mWhkL1uGurTYRViE0OFcI8fPEB1mNmtjOPjj9qlwU/9ZpbM4pMX+a9An9CuP2
RkNksT1bk6+9mI7/b3fQ94cavflHnGDmOAxFnSbMlb0+M+Rmp1PCp6QUH22bXvOM
lPX285qxs0K5IhkoqaYuOK01RmU6kCcQefodwRPFKvb54N6mqFW1Q3f9yhpzu0sI
fD4BV5O3iZ93NUlMAEcnge+PSuSEAoZRfV5DxQ43YbzMBYtJQSXixxZffwkYGXFo
aOwkDc5mZ7H+OHbolm4CD9yQSXw4M+hy30pnyxpzdLnP+o0i5QqOvBsOEtL1D87G
Uhlz6jEmu4CQb/J13kTmXHkqGY9yIwixydkwiiA4bsbhtrOaHyKFEMsubvodvw0M
2firTBmhkcxmoClgCOZGLltZc/kPpVFmZJMB7z8+RD07YgDinX7mi4/JRbd5c+h/
Keh1sYzsS8G7bEmWagrgMXRuJziD7QgQPXZ2BVy++nCB8OHPXpdrTQIizZx7lh0f
l2DhFqcNAg9+RQxuMpQUXtKRancILoWzOrP12Bn2Vlls3PMBKsl+zmfpBxj0HAgB
Oogqp/vNStxuMwMLtKd23pdmxGJTs1U2ThFQU1TSChBHVGDbQiKPgz22QkaarNfj
B3UgFjdCEZ5mgH/VUOA8iYiKqVmnF2Qz7Sif/1QZoMcbDi8Qm1Bskkj+TRhR+7D1
/RuOapapHQJNIomz/QP4IHThmcSHI8LO92DuRhAQ894JD33rVune19NeLlQY0TgR
23z4nYs5ylpz0www4gptcBt/42hS9hEpDIvyOKXjSItssSCq1cxvANlxQ+8Rt+KE
O0dhYGRUoK4riPJdePwA8Fl5DWEcMqilAoaDDyYC9Yv5U5D98P9C1yXtEuQyJEId
iTSSkVj7CDqwTKIoRF5bNiz9PmIXlxgZ/So2+IAMJ1kCKasTc5pd0zdlNqYE/Q6W
HwNqrRrCaDciXeH7vVdFPiPPInOFgIMOz9Hh2IbOmy+j96rYb3TPL27t1uzdgOZV
hmTGsl0Cx8oYBNbs+wXjhX5GpPZZIN1/PLEML60CRuGnLA3n5/UQ2TU/F2hsyr8B
tgs+N7gfGyuL++wu6RRhAFRVtCuTCNbWVLewzB77MA+1pb47tpol8r8T6wtcSa0F
MhE4CEQeEOfRAWdfP/fgZm6uV1sI70JPkPYTa3i5t1ESL8NLruCzb09pIzlmhbGf
FnG68fPXRWeO9T8uBcAqldsngSoF5qD/wzBpvtdHO9+LY2W+I3vfpICNKJLrMkCy
ISnXOszD+6qazoltdqnF9q332Y//rWcww4BpsGgtejf/SarS/Rw2MwjygBeA26/4
k+wxMqSNfE9XF/E2aUuusw2Fc5Tf1elT5mcDpK+BfTaG2xV/v/DSpkDNPOV+rkp2
WB8o4fWor52Fk5OAzjfSV5P5o7Ki1YYMUf/OfTL6DAgH8ZK+fuYmQfIMyce2F0jP
uALu/eK715jXTWsMQ84JJLRKnhu4tZDjBEPNaFpT5HWHZJhD88p+pztVoFZ0epAH
Mbor3awFvlHNJ7sfCYOA6olN4v1lIZdK4fWTfOQtQZ9ohlFXGP+cReTw9MUj8TxI
GqJfBVBbrppD2M44mvtx6KuHGkryO7QKtI3Ii3SN1NPaWXCjyN9sqYxW8VFJhOow
wAWiHZA50n5gfqbhBewMKHgb+4PXf6yrJ7phmOPwdh3yp0mKNyjwKzkB9wql34Jr
FuyXLj4qXSCQB69m8YSYeJPRlNt8zt9jXdex8zlFzXhoZVAbKCw19nMRm4MEe0FG
H1FjvIFvWgDCB+Bc26oHGT+tVe9g/Ppm7Z7H7rWS2BsTdebsVnoll7foAqfRaFSX
ElxgJ/u7Phbycs/vkX3J+zqRu0uLDsM4q6OVMCIDmGxRvJVLAZmgMLymP/q82RXr
ib6lsaVc5iB/nCIOv+xXyU0npRnd8uaGYTJuB0nTBpKiOU+4zsFB1xGzKAM1w33/
3g5l9Nbvod0nDZbMtV40YKVx20s7Ajs3OBxvkBvm367+tYXmX+sGHU824OOixamo
efFqcCNhh2t5R3smix0+Ur9fGDzkhtl+4m/hqW9/VEIrXL5z+Wp48zKjBxKs6Zjp
ra7SRNK018NIGewk4oy5Swqe7qnAQ8VyIXHt/djfDC288QVQRgPeDifLeade2J6O
heXyPH20PdE6xFgrt+Ez1wldTGGRn0cnGatAwvsnzUuhY1JlueXRUbPZ5TkPIlXH
oILc48//chhnIoqJOUSBocibtJXT+OCo9xxxNaFbM+ko8xdynz5MmKKNp0hmoX5v
Ph5++2ZCYLXIjebRwxSi8xjgtcHW83NegR2IplSj4JwqJMrlN0a1HCa3ivxy+eMi
FUa9YhhtT/EzBz7wE+kg7LANIEIHfDEGNcJBwp9t8kfiSMG5AVL99SJ5/tERFU9y
vIZWM5knPcpqAIiDtmgQRwHarEp+g1/Pc6Y4rOgVxvzvcKsh3MdCHa6OtDEvh0MK
XYnH44tE7eSgHvP3fTmOrKghvl4GmJ+HQg2HiBnryhUpraLj2Yi+wdXVZ38j/kgQ
54VEvXEUHoCsFp+TZ3/n24noFKvPJrt6bjeT2BDxFtYQ5eqXTgYZP2DUkdN8QGr0
qfD55vRp/eZ6LXo4x/Wy2MmlwupMgq4rbYFUOly14Hpo2ul0iUsNypIWeIlpKeHR
dY/7Rs/iueMfCHjohABVn/lA+X27DCcoawX0Q/+7Qt0sTSQmR+BOWuktQGC2svZt
N60fUhVsY0GhIUhU9NeWCfVC0IOpilnbor3bNKYopze1y7xpwvZ5nf1M3p1ShQdX
aL6f68rr0ELbVmVKSPt1wC7PmNSenBrtmZTy40I8BtFoMDSJy17rdjii/dPMXZIL
uaTAnRYljegrLe+65Qn5Hce1G9vikfGrv40EwZIWXR1rq67LcMUWIUsGTgbmcNY+
KMzBPWvas6bxY0GQclw8Fl2m5ocRM17q5qXrAzh5ZzFZQ2bXX4uHrwyhuQlj7CKQ
QBzGJWV+5UtJ+EQwdMIVJGwwbApsjsOolD1XD1G5lD+FBP6QNVQKcZEa5cbZfftN
roqXla4XHwSBCDFFe+kdSHmh8IE+I53s8sgUzPYRJZsu2xZlV+CrOp4rNXzMLcEk
tdDQoPl18bIydATDOI9IUaCuWCC87rhk0UpjhKrCONq0SvoQJ5rBn8wC1Pb4K0ou
bNXiDFHr2ur4Q3zy92Slc04kfbALWcWggUzUi6KTEV1pDtOb6wGEPT6l4jdcbbZv
HXQcj8v83507/gYCs9i0o8ID5i5KHzssa/k6bVNvMd93KkgEEvqPB5TM+EsvMQDT
yxxn5KdgEgaOTaQTcG/8JtL3j5dXK66DOjXq6wwGM30uR//C/uNQjkEMX6xYsQT2
yeJfV3DqXl8oV3tV9l0n76FP6TvZOa50oEvoFNZl0BNA2LZ+9+EiuDT/7BfxE9SW
q5BWLJEq+BLmhaKo5PdxscPd1A68i4F0tLmijEaUGPg5BxLvoS/Q1EeJ+rZvRFGN
hKHVgFV8FWh0yvHsZhKlQMdoxBoAdxvjpXWAqfBd8x1BmC3Jem6fJOtVRvg9Z72F
PZGw1vVpbe4iSpHySKehLnH4esV/dU3QAnD7G5r1B57y7aDU02WGZJI4Yo048G8l
B1Ji9u/hqPoWcrDyXRVbOxqLeLbuOi+DMo1h7vUrL1J0DC1ipLky6YIrcs5oUq0h
M5jJbHOavWWbcZ6vZyas1gbrVllwPxMRmahdkw3ev7HrPdOyuYfZ+M+JoYK2Nbr2
wknaQF1dOLDGMMO0E4bEsoZ4vS++w9cAtbapoTJbCeykOlviHS1Xz+m9TLQUd2/o
Lqg1kSl2zCagtoK+jxdx481K4KXfscZs6CEKWR6K55g4Cg9z9wVzUteazgFdO2Bh
K5mv/T40YhD0DvBpzYP3fN9x9kWnLcyVEkQQ105MVxM0ZyORP/PwtxzV97NdrkoJ
TeGjso5XupgVbLlhoUS2IQU3EFBbQ0vZRUY4TZFlRQxgRVgT/axNwq1+m6yDNuwL
tenk3rv05c5osJdU93O3sYP5844E4iabkglir4KgwR7qqQAu7iB5lGSVABiWQ3+/
dir3QZhSk0hLwdaA1PleWRQl+y7MCOlvDJtMH9HvVYQOjmnKE+kzYhPbsCO2T5Ck
2ztFKmXvgCQJVxomcaY1S4zEOYvBi48KV0aZrfP0q9ivlo/77euM2nPnOTFvfILq
20EqySDuoI4KyPAK64PkgNVN+z9vJWlUCqRB1aTzGxEAx/GgnbkHmfUwBY2mdF2p
+Hbn7IJCJBWVeppYZkGKlVsTHc8+kKaFEi7DTNiVA8cvaraLm3RSCzdNQLYFcs9e
f4jFYmPBbca/9b6y4lkrv3nygR17TDElz9RCbtXG44DyyoEFU4M/dL3DhBFECPOH
5H8MsKWA0sOlqHwiNEFNsqUalHyn4w7IhBKd11FhYaQar+mh5Kq2FJlYkSRyrezV
UoscpJmSwFPrpjTBuG6vClrYShzgUlo2lo8QV0gjOcn+3oQKBp6G6TZU1glkoCZu
efdfk4gcIoEelitvYA74uk7H61sQa68otRPceOaOKQTnOo4Fbxu7jJNXb1brv2Fr
dfk8iOm3OGEg/NhnZEV101HGIJf46drf9bgmUaUZghCkohcMNE4Kmlds2WVFDYQg
/L1aACMWBU5xFm5H2msGgrAxRkDO8dwWS0xyxxatoFpMxgG4il5YprPlsuWN7/ei
/nXkS3tORB5hoV7rpd7VGPkhrilt3h2EHE1V3YBTPqsKAwEAn+QcRiTcop5nIFRK
Xmv7//cjfo7e5SPMGINbFWtS8caiNnMujVhmQJhYfRLDuMyr/yRTiJcSZ+FPxcOl
SyB5vndPvXGqJGvDMtqg4o2VM1VVqaj8FK97aDwIlHh3W5g30PW9QTRIlLrHpAUs
nNWizQNOHVAMrS9be2LYW9lUudun6D1unpFOBnvJ20Y5dc9ySonkBT3H9wRLXGsG
twDicwelG31g3l6tzZC91M5WYj+JE+QzP/Cmq+WxdWDTtYXPT58r1C8FxjcPVLgg
iQIFi1UclK/Ex39RUa3i7uI+vDAdTfLoOf/z5wJGAxwZGMToAKTDL9uGeHwu/drQ
L3K6cTP0FSc9iNycCWBnnycCSRt/zewhx6UIVVQgnbmDhaqFGziiqwCqXtZP9Q7W
i22OhGQPVbtlhLjRH8hVM+DZFGOPzRSyEzolcTUm1aR6M3id5QEJ6D8N37l8AxOy
QO04BDd4nu6rXPV7ScNR7MlWnsT4KGxjSBKViduHp9j0mB1Kt+XzsPRizAjb9s0/
JojSSYmJvENHHX3q3ev9lGrWko39RXtjWx5uXv3EpdrRDX63g2BxtfbEcSma9wZD
FnaO16COdsNTwKuCIj14gKM6fJapfgQJw5v/sXg9BSkuxidiO89KCN8l5AQGKAg0
PEWbDU6MCguxkRI39TCYMGMinOUPhwE9JCuq4WVmY0Jlgg/WiUforh7FmUYcASBE
G1zNEp5QQGTSRVBh45GM2zya6eDcesie/059ZdoXXrZ48QHchfEU7XeOUKi84pPd
lsfo3s85p+GBp4lbxxVWx5j1xjsAsSHww5RVvb6if/qwBr9qqqdaBVeOZWy41aL0
LIYbU5gPdqvlg45A+t/F6kuI2ITZroazG+6lkDHaUWAxS8g5pd9gnEAU8pP/V5Hf
0FeSuJyGKg4+5kcTCkTfBGFAMJba+58kJ7UPdkPS79/vqBrHXvlKE3Q+30ljOd/r
3J6VRxmpcqCUDVSRA+O0qVISdCyY/74CaqHRny7fw9pOkg0iDFWCV3ge2eLhOD2X
MwNHmOtHm/J7H54Ob/iGS9ajy1CehZiTqprb2HeEW1oZsxM3mHZpIXg2kTgeGecC
gfAe5uWhfIPlEl6MLzRQ9vYt1TSoAxsTsgXakgK5cnCnBo+g3i5oBxA16AuXL1l6
eLQE0iJl0A+/K/7oPSSIhCakZ0uOxAuUZi9zkTQ8qkujMre7Vd9qQ4hwWrmvdCHK
VHXlrNpDJ4J633f/fI5pRQPouXhvt7PGDjLClPIfI7FJbIL72XBLhiovwrv0cwQZ
TtKlWOyLObNF1tYsLU8pvLegHPbaPEAwz+Dhyms6WLjK3iHqnQkoR6hWw0bUCV0c
+rt4Mgki5KEXE7H3fqTXrk07Tzr9UAlYUjKTqhzbMbMr7mlIHwn0gTmM4+Ox4xWu
97pKpPIyl5IG8zK7j5WCVGVDBJbnpb1qmEXVD2EO3+894i4Qi6p4flr7gAPjRQQx
rzYTvbANqPQzBSrI/6lhdLO0EtAzmDTO7bsG93ND9HaRkB5ZTDXeZmjanfPE2U/S
qMmnSuJiy5rlY7hgd6wKoy8aaukeBUtSBya6OTIytvgcshbdrF1o4d1L0Y1AnxrM
0gbq3gphYeUHdqzedNoemxGGM6WGtUg6N7fQ4dzb2tKbyNnOwyOfrgjSAUsWUd6W
A9TRBDiti17d76Qkn+XsrhAUi8oRnIUA9oVmLafUkGoG/rd+pKU2Cngk+Nf2bmAI
pn+byY0vXjgzHNnSbgQy8rBtRj8k7Air6GqhgKhBCwYV0Jc6ue+8wD6UE+vbi3NV
F1PbBGmQ5ULE5VDBMnaBcX0Kjk332aK2fXCwQaI58/Rgr+bnKySWrNcD0IDPpfUB
KO1iUPBDvS9Kph+vbl5tJ4HpwTvHmwO0c0stQZXoJ/rUeUu+gcwzQwoN2GsvU58t
Qfid8/Hp5JyqwMrwzHAGAsXxoiT7T776vxemhxs+FccPaGEcZ769LbGKFIyn6tAH
g7eenBnuvTQY3ZiermbiKoerr3ZCVeQ/zYWnEsneycAyLxXG4AJ3OnY3r3Kl+ixW
uaiIxmJV7yV3sDUTNL+41G/HiIiSTA844B9Fs4n3cqWpzatSULrr/xZT5ldDpoO2
ymy/+VKH647RvoxlS2QXSjnPrG7lEvZ7RxLLfi3KHanxLuT0j4cvNw51q9rT6Ajf
g8MakdBxzkUr0IYGy6SfD8IFt41uLGp/IUlXZtmozLmIIOsC/TcKjLSP4m9CJCND
wO+zaQ9v5eqnCPuncSrIkhrRigIIg2DCRAyoYFvAhwpPbFYeFU5hodxakoTqu8dY
ck1YjGA0XzfI0bTVSMDzH3SEyZW3WAkVHlX8sNKcXjq/PO0likH/JxVm6AjQ5Euk
686vFxy/pG1hghqD7B6AJurXuwqRkvw58GSN6YvWHAH+sKyhyF5oWu1X/ui2sl55
Gxq5jtSOG/Bs7PQKMUQkAmQVfS+3zukM6AZuIp+CoTkCvdlt3/6/fG6xe8Ny68nm
9xjp66/8OMnQnV/Q4RQFUen6Y4FRIPcMRuOqDLVzgw/ZEJWQqUWN1mMLV2CiFzwX
YE0VmZCN8yJBPVtn2Snvz7ta60Dh9yaAbIt7XqsirVbXuhNmf9s73/3mxVTmNgo6
DFYssjXuGQ9QU4VCUU6/JGCB8rWmaZ+SeOptiXH2AE31WDwdeXzPkP5rk6q9OUBJ
/6v9iZHiW9NpgcW2XhW3TS+AwcxRtgN5yqKc1cWy634GHmi44ffKisHyuojH48nk
YgpOv7xrfG7javb7WLAuwJNLnCuApHX1/TDWdvMGsxF+Rndyz/5gTST1vWHAlpOI
qRTpYf5olfJdBDULxinQU+20h7qkuBcaO4lmW7eBjMAzlLqJ5Nv4P0JE92hy+S3h
AwnP1KtS9/yp0k9fc+VXSRE2NzER9fYPBLp9ChALb641emZdKs0KEJLBXWpT73AU
8NqTfLSXKtwwzH2vS2NP8QIqK3Ih3rFjeg+EZC4u61IHkkXfwyE39nKPQ29Honhd
vaQAiNWSAqMayppM8DQT9YTmvBtFVLCZJ+XqJz7ejX+Fx24I+z7X6ikvaLoCJEBw
KmpfyOuLXGfg2mXGoY5BV9dkWS9ffDAdzz4/k3E/HhvqxTZiIdQW8qLBOvJ1gW3h
nl7BecUZLUbA5QeTw2vBkVS30FUcGmP1LApxJML0zGQR9bV34n8+rVbMt4Gp+e3d
YL0Nx/AlM4qR4doVQcQzQeXGKT/Xn+VEksJbtLm6p6GXOc86Yn8FnEtUczeWtNCP
YN2+vx/9eyjfdlO27ppB4iZ8UoU0dI0b10Cwqvrr113YBxADXFzztPiJFqAS+4CM
2Bq0qE0LnVKSNRiDwltX+IMlbnd2Nun40ZBAe01AOSgj3lEi/jHGPwndodGwDK3T
4BdzdGDTeLU9dQlKGD2K/Wx1/5wbvGK5fGOw9Db1fbu6twT39NHt+hQNO780bsW5
zs8DVyyMF+G2jES0ax3ahO18swyah5yqIY3tcL9kve9UFBcR21ky3lNjrHOz98ql
IhJO/fkSMJjN82dyU4fRBkJrrFeVIfYVmPzNKP8BsVhAzUXv0thY3VejBvaiY0/B
sE6Gon5b+zyRD26uQRmDUgEYHEhJky/9QuelHJ3La4NFpOmSykUvr19fItraYYGE
RmZLUJsyUXwBs11H9pSKsiINgsMK46gjh40/fDvG9PRZhkH5gbvMP2pBcUlQ5zCx
nqPa7w1ZsLpFvvqU4BHlIGwf+FzVjE/XR0DjCyowAQUT18lXZQQxddgcMeWCFDGp
jznIBVUia3UVqqTQyXkt9dF4oxxhfqWf/MaX+ngdrGBHRHJu9dnYagr8T+gy5LTU
liG5zMf0q0pBVcg5KfJ096VRjeCLok1JrTkPJoAUc78zi1lO3ieAB9hbqoFB3Mwz
3MdhlIW4FZ6/Ytq4p77wt2WtODp9NKReq0GkZunW3BKsH0HAAgGkmcziWzfg7KcA
M5Ys0IYYQr87Mk4XabsD0Clt8VJCiZtxvi8Ys5uR1yJ6ULHnofb/lbbrY7o1Qnc3
G0kLokC1ca0pyJf5EjcBNfjv76h7ROm3vh3HJyDsuCwl03Oqy3XTMR3snJophWET
/4yCUhplQU4GJXloIISF3Htu6AuMclarINd4E15rDFyKvWF+iBenLiTBTTd3TTNW
CirSM2YzB015FDUxXA/o0kClLbdSf1IGK36nnDSgKHEDfvcLCBh0pUCHucrDaCyy
X6UhPa72OXhcLP1HAddRlWV6pVvKlk2a5NN631DdmHgLR4PLhOnfLAK/4GktQxxq
oDaafSwp0C93dvs9t605w7FvfEm+QiLPY7qxUDTg/OKLR3iM2YGGaQiLw4KckxRO
0WV0x/pH0zXMV+iso4X1xIpTE4zOO//DOu9JfiLFslpx7WCnpMOdUdo0/dx9+zjF
mJjlTZZEzcdXrQD3PAmgzffaEE5/uBTAJrr7OkmXUbnXp6PSbjeNBc1xP5GwyyMY
fNtGTzH1mcVu5tcTS9KbdIcuh/UMIerGJcQIXiKYZ0gQNwROv1WjPS4/J8hLL8GA
lMP4i6lsEuZ5pz/Ubp8L8P1anAW/NEJFirvuGsAyTvRC+EdKRtkR9spcJ7hfLcIa
PrBXC+Amly6C43qC9upIKVYhrGMJT0W3BFZevZsaBF0s3WN9S28wsUOQsgXcLY1e
hzicHJDt82oObADVPRj8r3DURJXPSopXAi4FKXTmyOiFxzaUNzXjMf0cnooolZCn
pB+wSCxY+MwxE+E68vkK2M5Zwdsfay/vORDE4jTWDooFL757Tq9sN4DOnavZTT4I
i6MwVpmrMbtHvRMuNu8NKmGTFG0yjHhNhOfY1goseJIQbzDBXIzDQcOoMFTvYjDV
anzUjBfUcZGD/T/LFLI/3kC/wD7p8xQvhv7/IBBXEWvj1n4ILkW2Lp18q7NCtey4
GGLwIKKMtZknaiZ2K1hYUTX3yOYCGVjhVUMTLzsIEXjatFA7v+69xHPTjmX+PtM8
FmjBmcWYptg/SxoVh+X/bseDUQWLgEcRO3I9ZRvrpCYAUJC+zmqSl6fDnSHXjoMu
F3uT+ByOUgeR7iT46RpkANHYYiXd39mQZqu9jwdo0v39WoXP1Sx3fZ/lETnvv7V3
NAMDIWw4j3jP72T198y7Hae4UuzMPaXted/nOhxx2lv8AvMt/5v4yWaH4mQiqDiV
w+UH+lvtB+knJlQnLOvKE8i1jmmtD9m7Ovdfaenxdg4nxFAFEDUP1rnkUxIYt5yD
+7xK7fvNvv3sw4U0Ew4/8lU0SotcnZrgZfUM+5RRf8E3DbT5oDDARocLwERzNJwr
JFuClbNyaY/0RYXh/KFKxgc+kNHxdcnnK/xPZ1Yb3EXqicx0GNOZG0DktDStgTaQ
P4/DtuwNClu4AqvU4JsFlzL8i9X7pIqCJZ7qOt2aSsRPb4mvAZiMeLKh/+F+l0hY
9cTwwICTi6gpvTktpEm0GgdxeH2es8bqRArlQrKsRDdN10sn1s81E3WnmDfL5eHX
BeTMUQ9k/Wr/cVPW6l7pUfgt0M1xPvQ1QWKW0wMc8xNfNZvw53Q6kpcnEWD1N1y4
EvTMeIhHd6qaMVGlJ/KIi3PVg+dEss++owcUVk7O1V8KjX39c+Uw574HzXSbO52m
s0NkhEeFRQKGeMT2aQ3A01NG4snqtlNZiSEqLbFPu3xvL2mekPZYxOyc4UoJKQ/f
J5uHlZKG1vOzpKqlQjJ0++63Y/f0fN9iNMFvNQUnP56pUjiCeHr26e03f+ffisel
9PHKa7iso+vDnBEho3bovCz5FM7iCok7qzARr9NA8D1tMdAz+HkDHcoz4SaZQC5/
fgSpTVjzPgwC3M4S3LMDd7dM0ZzcvkMCVHhkkmqIb4XkaQuzzzr9P32uyRwDiPz3
4FIuIL8u7Zjr9kI42MZJY/wXgUNm1ZyI3dpuM8TG56bRaTItQDL8ILLhu8suB7cc
TyNPapugaI+iZtgmL2CvrWmEiyLlynuMCPsxPEuw+WYmZS4JEErWXrSVG8ybCVSP
TLGW8fgZOVDp8IPwafYfwtgxD85a3QKVnVOJYBLhNAW51KkTi8juBRL+YD8oFKjV
lfRtTAwncxHLx05LPwdlH+BhHlD+Oob4M4f/ORVddNtNc7+UKCR69A7Gt1JtoOOq
BAbnnVIywGHwgCToiq4nTVc4WfvQHnNVfm23f+4Wl0zxYwza5TUpByCkAJXSnbPB
1heYhEI9Q+sVGfVXBYdsiskYiV4WwMHd4TsnavOs5qGxZXKXJZCfTN0NTN40uO9t
rmYe7YLsUgjWa1isEnJ5LWHCQEXHxSMMADdLA4GubgD/av34GH/nfQDAJDVhsKlC
ytI7jNDEJ7PZftBlofoC6uV5wHBxeqbVnZeRy77o3/O381u4CrfdCQMvg2LVmM8g
Vdp41p2l0sz5fzDMZOXKZsZcSGB+Bi9L/Tkm1YxHZ8n9KlsOmZe2r5Buu0ItBXJc
ltdAYOeRm6/sZTb7MCJ4HIU0opw82sxFMdQprxGzoHYMqQwAJ1ChWqvGkQ1Iko50
pD2n8V7ozZb2TBE6X6Zl08HrYPKDhZBMhhMDAjJsw126PFSsl9E0X0VsAmy3Sv3p
wZDJzsgLTmJe960bmJP7v1ruJNcRhSHjHqITJd2h7Ejw5UXuwlHQ1RLQK1BFbnUs
RU6Ys24e2JrQRLVo3CNDiNuItbFRO9pwDM3YuibU+jqYJCPS7YuRtYMfBbQ3OPSb
RY7O+f4bx8JkGPXr9uC0fau40meB5aiYiZTzuJs/HzF9qXXzoiptrSUnsx2Pp28i
0dqFoWFhQF2Hc/CxfDjX5AkRjXO+zrM7toi7UkWuTrz5JG8DrEeWNhNe/08ylCUG
PBOjiFPx8z0Tla3U4fthOqWuaCG/5cdGjhMCUTbsM5HWd+K+yVwlggXLN7wZZBqH
PfmJobbtdna/7d/a6QTEioMZSXod8J5oGDKA7qoHpi8L8BhUDz8I+mXI0G8g3Sut
GmALh0Ja09G8QrEkWl+xtFzxmuoL8zaVJF5m+z9SEu+aS3mV45Xihmf83hACgbJY
+X7J1B7eoNFo1xK3x3QVRELrUMXI1RGzfTHbAxNqlRTpAlB+PDkmKMAjV+vgLEfK
IQhI1ZOWSprHAwypLDgtBOMD691TQviQUl/k46cmUYne5F6SofgUxLCaxwJfQx6V
fj1+ONnwcdA2s4zR05RY3D7Q3UMufEpPBWanBrqcfycrv7h5KX+ld2TIitKJ+fl4
zU2MppuCLp1BTGTeCTTKXpngZS3uvfcotPK/fC7Myd0g0KIuGY82ObePedLeGrej
80hK4wA9esfobZwHjRRY8kMZwVqbHtSb0JDYOih05CzZCgd87aqESKr9PL+O5c8E
ifAHRInw6UuF2m3L7lTgF+Y/2SHqtTWENcTX/WwdoNxJykDkTwzwEhL8KyFALJa1
gF4xObLV4PU4p2Rn1p4HjP2qihZ4xpmpqvVH4ImlqJ4UWW42ZJiBZN9y3+lU00je
k4fauwQpVCb94FOn6M0PeE1LUnX2Lg7VOlxZ4Bt7iaYITimQA2Yn5LTfhW2GqVzt
TfykAp+TDWBJOBGp7O6SPLiNbeFR9wuenT8aQuy0m3MzQM4GIZ/nJWB9NVBSOTeD
epkMWbVvI0WeUCY/Rh7Z7oXDPI/0gqF2kU4+Y4s6i5Hgu8QLRfgQY1TsoPONbHd7
CC6ydIqLdRfdjekKg2SvdXAdfZBb5F5QpZoBEe/pJwEM3c6qPfFhisAoruIAdxda
V/0x/yD83V/fjzTCF4PnHBj25I6RITa7931OKPujeYjEdrreu3Sv6Vy+IDt8MIEE
OdVnViXksKxFTdL5J291zpUFN/JuUM4INXz6F/xVwFajhCjI7zGAoIm9hmH87Kdp
QeaC/W/o980kGz6nhBDyyZBR2OOIU0HF+DEc1GCzGqCNgAauZe7B5tRsOv/+/j53
RnZWWE8sKx89rm8BbU2ywsHlKIY7OsdGizcFh673Mn2vDxsFjdcniTpdGAPWVsaY
o5LRmzDiLLWKnd226PbwCorujDCAvjZb56y5Ui9S003PiXMjbdPuzSGxbg2WdpR+
IgaD3aRFj5V6EZlh6uvVnX0CcupWMcWK+w+qCvFAEoXWSEFZH+/cnqnblfWyG/lc
dbt4XTlrI4fNhrbgEGFe0JjGduPjH/Cr+zPMWAtIHhb6IKCxfWXQOzE6wAYq/59q
br4cM+0JQu1j+fDmZzJ7zikNgKd09jqRI0Ij/JMGanaAno5JJrZOzoAZZslgJcWo
MXVQhXiIc2xnB7CIdi8luHIIFeaZxlQsDKDC/u3wO6ajd1g1iJGR/BwbBYLWd999
P2m2loDdtSY6H6QO4/AwlayxV/aRDKm10J/Swp+JmhjeK85pW4P3GnTjHVNhUVbZ
Wb+LGigknuc9c29L2E6Jt9AXMXlh60EEErUvEkk5XpBWYtYRbLHL9zpnXFiXvp31
eSzMs7LUaQ+QTJ7nXH3meK18SJ3/puC2zHtnnUkofwlanU48wSryDt+cffhPo82p
hPmid6LW8KCXrwS5wHyObUX0oEdWBTeGwMbLr1ZeoigLdm8AaEIeTGzkqP//B7rT
PD0TVdtSSTj51hbp5ZpcW3gf3B1qiBOwUay1MYhGMDCjGKUMeC13LqAbC8EKM06Q
4H4XSI2B2aKf4XHfC+v8IzXpV5VUHLhJHGhkuu8wfJZ6c8SGtkGSVd0BENdRWirM
45WW6GKtq7XMJJX3RiJEto0wGf+528h9F8HSkqMXfFwP0zmCqwM1EGzdZ1GrJTkD
tbmWSX/21hL9KzBWKi5ILamrJ8kZSjEFqkzmJeUX4L9mcjoOIgTU4a2Tb1t8cK+P
1buc33i0UpZ2sDxBSi7xNc3WF0ZPsk8acjBLCRKmY3+O8YUQNygHlsKCylgAFGvG
861I9vZH3xh9XSzZ9Z56OsEPJTI/swapZiD+vBzOaiXtQiMB3W9b6k4U3/vsT25i
aAMcQ9vNDHT0VuObyo9E5ZpZgOf77KroS+6bGOfvwypRulTwtD2hCDbc/fPgKkA5
ZhsnCrRvvoCnfnLyqJsc+Gz7dv079pdwlA4C9tK5cQ5V0qRL0oqAmuIz4P4WFLL9
wYdCAqrSv9Xw2ormu0oaW8WFk5PqiJ1h29Zpo+xruRZzwaS2bZCrnLhXaKmVsrRM
QCBfoDX247z0YaRw4J5ZtnDF+Zm2x+QtIQYb0mmV0Fa/HOKbMVnBOr6pEkVE/Cbo
TEViZwr/VYMEnkW4BA9vG+IqgRsGZqdWDXgWVvODrYV3UYoGuvPj0stHbMWb+W4t
2oCQXJXSXBocXXlny8sVNc0Ry0YfgWJhdKhOTfI9SGGV1lOiC5jlhy6q6VV2amah
dPu1GDcrUJc/HShwmwlzWg6BcRuAssMJa9sZVeeZlYjbK9YgxiDtKLhD8Rb8k96o
3j3mL9EsT7lG9yQA5fvPGtWDOdlX2hJYPwWLRik0R2Oj73uea30lLLBYev+U+St0
DGYRG4UKCPsnUO8a2wX9CGoCS/39gA4SsiBixHxBWG9akNukPHz3rOMK0LhTGPQQ
amMzokuHY6dLIhwhRjzCEWw9CR4Z0G9kMe+HMk8q3VZvXLH6G5hn8IHF2+YVGnxh
4UHrRKDzeRZFwTrCiIvIiGh5HyhkURbUKukzbTGU5xUo/xqwHmfFDZBaSMoDpBsC
B+ebAP0LiSIQKXnzQNFAUO3Y68juKZk5DIOuaAgfKqoH59vr/cUKkf9k/bmfx4H+
fJVdLDO46AqJGIMWXLrnWj8GuObA3D8bi5hfA4NTnHSE9XxoxL/5qs+bXr3eq0RJ
qE5/55mwE8qLh9YfdLATcjm4yOR8u4MrDpdOnQSwwt2EKrZ89niHNX5/UAtEEcXA
esQqPDMRKWutqxYvDRJhAvlGjQNSdG2nufCXhHFmlf7LJobr0/+j7bc08zxh8Kdk
I4QtLjNfflECyi710YILtmUhjyIujqAbnnwzeE61l6aE9YeI6OKP8aFgkElMF6aj
6TOIZH8Qppg2azpmHuV1co4StDVSLYv8ntFiUh7Nuci14c34xeDNyNOW5dvyiynr
f72K4rHYXSG8F2cOFJ7mU90zuOzrRcdS5U8Q0DkQp6zT97w+cPEbC8oiJRA5FvdT
d4iVz79rvQkJW7zeOa+yOw33Hm055G3vpc4dYus2OlVoQ+6tYecg7tV2nK86UkVv
Zgrpozn6KwvinvjMoqxQpjOqioOTxx7gMfaMokDgGNOWGdaOKWo98Ug3Zak3ghBO
FcqT+OTnNdoyTGcoEouiCLJIu5Ed5SMCA0omc9te46a6u6KQlFLJ4yhbeN0cbHtT
yqOmLxE4H7HKMIQrc5WpF64Ad0ev0w2OMDxZxZtWubRyNCqNcLMI05/6Cl5ijvfj
U5UTm9v98uR/ec6b1bvXpZG2CAbNuJ9ciu0SuzKGMpAidqkWJJxqeCeCdRbTd5Mk
EFRYLCCkQjvKIpvqTx1b5jUSWeVSjXzOp32WAux1aKge2oMOF9pegLQSygrwKpT7
D5LNDnV45ZeL8LAPixYtponej5PyfCAjJqNEvBpyoAxQvhcz5Sa6HauwaDBPgjGH
Kyju5ZBHDzV8/F/3Rn+denO6IDTq3dS1ekF/OxFtsj+Xnl3Idr6h+dH9QqFNcS0m
LdDufsxf64NoI6aWBESbZ6GNN554PtzS2xnQl6zhze6UxA5jklheC48uS3oKhxDa
rILdVN+AsIEoNFpYQ5JBYlwwblTwpe74qaQdSEHgDabnE69xv+h/JKbwqLYFBwrF
Hbl+L4E6O+WvTGQ8pw7H/A2dXXUhvhQzrQW3GrjtaSv46C1RfsburbpLvNK0uZl6
UDxwD0jtu4izaMJh8imhYkySSubeiIQ7Lm033u5V71YDlImkLsTqVs/EcSemGIB4
e2+4QyipCbqwrRnYgbp0uhSekgFZwy6xlnMjE0ugMZKuoEO8diL+9AShOfnIjSTB
UQPmlhOMPoBNn5wB23F4SzEY2EPCDXZ8ZtV2H/nkRx5VmbREjSuknk/thfXxs1NT
j0NosTnBbzPAaZm1Ljzv0f0C5ZykPVTbIvHbnC+vxzAGZ6hY9TYjYHsPB70o/2EX
SO+t1Wa897MSmp+l09I5q2vvs3M3dl0gnyaVYCMcRSWcjhX5diGbxhaln9xEyUQd
/gIbNkKysFyQbk/X7rTdDuWU+j6Fl7CpfI2I7Pvwxj8wVQHKOKvuDahPhMaGHw3k
FM6/vvgqdduSpDkTLzIIjaVcPW8fos/x/2oRzml5kSZpvZL5olkOnizHCdtwvuoc
Fbm1L1eOKn1aS/cwMkRurZwCxwztoHSUzfiBoSApLZjuAt9iOzKS/dl2cXsFmKcT
oXHjKGGeNnUaBpK5nOFAGEuaoqis8XsKuNLbQeZjMUkXCbhTYpcObGNq1xbs8loC
zCuwWXSWwTtbu+70nCWBdB/bMHzzuGvABoTL19N/9LPOa3LvLLkDqyLh/6GR84N1
m153GXFyRcV6zaaPphEVGmM1VjAqMhZE52BoEpQcRA6/7qpx5x3jSq27LYgTgqCs
AF1lblmXIqWJbv2KkwDV6SSbcyTfiyT1XPAy5wKQ1viBq29AiSlkW015BtR3rw44
h8GfTqteR3yHdKrvQZPBUbbyC+cSFzKxbvvDUluzHyJfornrgMp38nSB+MkCxtGe
6/DrqJm4M77dKaskB8IkR7ecmqNXzJrw3P9uY/4L4tUtIOetmJtFSdIv+LVcIOcG
1gcdZSUouO5hzBADFxsdzFJLPiPXtars7QcWItwfpiKXeJPHuKdCRJyCGOhop4Yb
Wlch2VKw02OyLVa2QytTxnds1kRuBuvBPxkbMGY96pyli/NY107KH8JoSaX0mki+
EOtCBCcw0zvmFFCA3xlE4jZcQk1Je2Tw5tfQnEi1jNQIZ1EbmF33xmYfHHLFKGR3
/aGcg/7r67XdzjAX1qe8tNyPem+YeA+hBIGbatmR89I1Z5EYlGStiVyrzQZ1oOzP
NDkdFzWtil1cyc63JEdfc11FPBjM00+fsQCy2KdF9EfdVTC5HeVt2GjDPe+NruDF
9ZkFFohvoN8L/WCsxdznDrOlHOcNKvuznAmRapbx6MNk/DjzdSkpBJe4Pduww/hY
LjwgawmY7abZ0yT+iUTavn9o8n+yxlPBZJmYydr0nlcbz7+og5wi7JTLjVcm5aHs
ZbO4L0eiQ5MqCtQlfGQaP3EoQ+FMBGamEDYHL8lP+rguW7Ppx+bpXLo4pRJzusW+
IJ9NETK4lEHUznrwKGzwJGtIjJYP7DvVfS2sDK/4ZzoI40JBN8fn0QN+fgD66dcB
nvetb35D0ORzJmio+18aiup8aEzOzVx6faiqGghGry4EXgB4tbakQSSsV+XWoyKM
+JGjeKxZOiqb/6PDYtfEl+EOpm8RN/MMus+mdwavbJuI4au6h5ildm2AtJjbQN6i
mdXYU7xqwXPXrbZFQAYfSIwIWLnosDErN8VgUkR54aXwZyrTn1r3ocqeemM7TzB/
b4anPiQLhvePO6dcsvj0TY+46fUHg4mYhKDAn5owt07vJZsEGOt8Nzv/eFYWnnUR
CgB3O5T/eScdZm55ANAicbGXOH2wlVVcCwhWiep9kdusgjFMs9+RvvE+vD+HGY3v
ygmD9ydwiLWBLcUnNLjyJt5I193XYMfkhlIqUJXgVqXe6oKmlY5w1Czk1SyLEMkC
HXcNddRJECIOAQeK0L5b8abQNX6qFcubRn4CQ7fLEkNL0PyFfBn9vlG0z7Len225
joe5E77HmZg5TQChboMgzA017DC1wqDcxSmMrdGU5pH2JvWy0oTqkTTF4JhqEfxx
/d1LtdKKrjnWHry7KtvlbLLHv93qKKge+davqrSwZCzCAW35lpV5/cpN3NiLsWgs
AcIWPAHsHHL7FW+680aDjxz71KtgVH4aK+U1SC1aTYgRFBUv66splv9wQ9hB8OmF
hF6sfNRY8sevW3mr4EfETbGu2XUo233Qwp/y8MM7rHLI2bbzZdslLg02q/2+p7Lg
io6F1CxTyBkkxFZKzx1eNtRRH7zUeTL319OAHfS57CJTKRy/3ZMcfaFdKOYkh1aV
80KdPmSv6PVzcLV/9A2U5W/RSiKS++9TfKVQYc1jechJnHoF1ncQyo8xZHNl+der
OO1QUHQzAy2+/rviPCdTve1ghP2yjms8ZZrW6BphyOvkirKiQv7YEZjwbnpmR8Ou
ZVgloHBDFue1vIwuDznAg0k5TcOR1e+FhSfGtIMYejphLctevhRKw9L0L52kionR
Y8pD6UllAT0OAeNmnNO93KzAYKz8U6gCTTsFEdie6w9iXHb5GgrmJ/RJ5+cNvgOf
NwGSE/yjGONrPkgAQiaxmRvXNmw80OuZDe6Qjw7uw/aV1zr8fA+Os/Ov/iUPSOML
6dVXe8I/yj75Xxos1ct82EotbYclDFZCfvI1gxx5h9F5DuH7lBWaT37TpHmWgje4
1EquSnuOfOff8F6jAjhoVjQ+q9fz6oZAYABYqj5ZOehT2XvUi38W58+1UalY8sRG
E3Xfcf0xwrYlOpfYFM/wEUhUmgogKLPMCJNCaMT01kbfT3plY5vAuP2IG+WEeQwz
mEXjH0fJZlg0l1TCS1PuKSzhHGrSuyk9+PPg9AHpOdXVBiq46OE1Uyg+oMkeCzVK
V9nZ7++Q2OMV7PmNW36nkbmnAl5Eq2x/oGqg2Kr7how9R6TU2IBD/kBJngU29OL+
DQAWxqCEMxyoYhBuU567btjH2YG0kpi7AyM8wQd4iZ2bDYcXmyHIEP6/hTiBT9aH
9h52FIRXbbLlOMMwXcWg8kP8zPaxUh1O/kOBDl9OWEeXVDArO6tFiD2V9NRdFL6t
YV6DJLBdo2JGKPZhgrUC2S6KYUtBtlaGEURB8DnXj3joRrgszn/rVgjuKM4QZ4Zk
CdzAgRcNtIpKFmobchPG7KG/HffWmuqUxbzq07kvVZnsiEac9DXUeg1UdWyjH3KT
m3GsAu8uEyYkAXfqMarqk7wOzPGx0qEkZkCWzjashWld8gMMLdQZzJFfNUBBk/8h
WjShlk05ZIu+IUmMADnKw3ugrIPhTN5e7OqiMUQu3eCosgwQKmTV1r/9iUxghoSt
KQDXfN3IUhv5sFhPXgnFcJSkidCw2Hv2q1dsERlsmFwBmTwtKTB3jUjQFIfUxMcO
0gnGK7sojof/8XqlmFQREA74wks/MjaaJVKrnmdwsUIRRQA3RIAHJlHd699nyMoH
ouTCg60YqcCLY70nTijqIoZk7Osm7yEUKLkdOMwINL+XDQs899fJlsH6uZDdVAC1
Klrrv9kInqFJ08FaadwFgNDsmW0TU+/TB5H04qOWyV5pFjezadeyLPPfhHJ+X23/
SHsMly7m6bm/zbiBzZcyMeZk+nstXa/vIVIJ2b+CC1Lh+6KgMkUZMHZC4chUbPiy
j7oZQ/1fhcJ/qhIfI5hBIjTn9NyVgeTLQ/gp8dryCGR5RPNSUS4/t5aulzS3vwg5
UQQmKmwgxV3W3GjfMncTQZsdhUisDS87SgsB+1ZNZ0jLVYxDZvFpMPEGOoiJSZfL
FpbD1IDJ5f6IyduZiEAz7LDHYIVcvjsafnGnRH3jpZVMq5QjzHCn6otIDKlS2XLw
psa0rYnuZ3hgstX5Ven2yV7Gk7rZmGG5juGchUfrXSILUhx/WA799tfGGG8/AVHK
sRfUGq0IiIftqJZ8WPak46p6xoVPgWKrVCRPpYvFk+Ps3hqzq1aCMC2l6xZb69de
3CfTnX74QdJxjJrI1nCQ89pnTQAnOq1QpFGjuXfJeMxU26G4R2ii7iMNDXyBEGfX
+a/ZS89520Wr4blndkt/wBjTI6/gt5XlKaqHjep1haSUtxMtQJm2+Ql7otFiuNeM
F/g27oFuiSGZTxh8NUJmz9qcb8vEdctTCBWnliy3VsT26XmpABDluSU2PdBxqYAv
Kcbq47QA//Ek6UQxqSK7oMxMH9BCahQZqGLcPQSmHHVzJSQp2ZbeAqbjNdsjV/9i
DjKKBdU/VW99Aw8XLjz2RJkkPLpxsclj5IR1Z2/rtDlfztW59QJ1SXQxVOFPPmHf
srlbCeztJ7nsL+8mlQFGkWKowzobvqu3B2J6I2QiX7uMXU6/HYcN4n4cEn0DaLsE
YMVc/JTKnEN5wgFZpq0v9+PlVVbEWA26zRB9OTJv9SCkR/zjEnHQtY7HLfnvTCdy
Bc8FlPf01Ahb+4STKBY6h+2G0vIX5Di1qgM7KtXZhKFo4Yd9nVpu7o6IJE+sFRyf
AtNNXk4X7VwDsYYSusDGCkr/m17NEQ45D2mTge8IfLuIcOp3iO4EC/mrjKjJr/NO
poDHxbdgv8RblGq0ve/VSqFlArn8lgguZaimFDHwBCzoqwxKZrXaK503Q/AaZGp6
euw1CQs0hK66ODn3P7l2o11+IISOMijlwkfC2Bc39TmTqVBQ0AW8eT64fLiFop27
1cOfpe45Oms3w/7mhctUeuHq7llyk7d9REHHtfdWcJi5HESja+ZM5hDkm6Bih09t
8uTBWZ3CDqcjrY4hIPMzAgZjJDd27eiEH4UNmzvs8QpqbXIzISqpGnD8TO37HEWg
X/FFiNh2glMkIRMlXZll5fdi7ovV+4rs6qU8CgT0svsqzjoLyYSTDeQ4kJy7UeyP
RSCfFj7tIv60sh8ASfAMVfyvX5GmoBAR/wb2RukZS6ldj+ND67DEYjXYrncibgHg
SOBm+kR3l9erSo4twRmSrYG4f33S9FYjH3gxe2pK9909ud0rF63W1Sn7IRqSbIWh
SRw+LbmVj4GGKp1mTrrB+m+d9QNJBKvD+ObYZEp0VfYguZfFcsy8QxFajzDyjoHk
yEUn3od7FwmarkV9v0J6ctdN4yNaEBHl5KJNZ983oDrmgAag+bNPQsfY2tFTROOx
65X+uGvqA5PMzrZYr1IKrgsI89h+cme0VKuS8ph9nsDof5cgCj+JHP3qVFQFWRuP
MAUvYWLDsn83v0f+XZOlG88s+5kUUGbGS/RHL6S1IVKkQJ3Swl0zdNOyTRStMc2Y
mBQmPoM+mKCp4qWzY7xpshETWST0VJctAiAEefoIFNSkogNRfWdvs8Tx0z1FO1Kw
NQauIH/bzfjW2qcX/cap2fjsgk8xxOr5cqY7Dz0eGQrRJmXJEjrNiRRfkDGj30ll
7GCrp6wuvh7mGsynP5whwYKKjQRExeKxrSl7xLHVokOSlm8WIw2oYrapLJiyi6tD
ThM7weCPtg8JNmaNc/ypAwwuTywLvtqwRIkajDFLmSE+ozxqLSKVTR7uilCoFfrA
UBtL2dbQiiQG9dTzTA/ZFyZb1XsUNXM4bF97qQFtTSgrE443pxMwHfmrR9qwAofo
Yfe2ARR/W6JaV2rcj/XF0nyljD3R77jwldsR8SyFydtlsR5wmiXDmGLEEfNeDLqg
NZL0bDSbrBqH7QKPGCKCl9kBNyG99jdkQyqZf6qceMcGnFFU2F84/eqon+Q8YI4+
GPxBEgi4fmtR3ZPsrRU+xBUHZXiI9ULKmosnnvn8nihPTMZBSBUOjxeZg89QYy4D
vOzwxGTjRZ7aqATM1dJSdO1bAZEtamdI4her8CVlBkVa+u76Y6StjD5yRRiVKx78
8PSCboIThBfin7N3UxueX8YqaYBHQ+5/vYRl1fstwIGUCwiVF5PzMXAPTh0KI4Rg
lSX+FVWq181nm0thGtNxo5KNOW0Pp6zohs8Rrs+xeNLA+tDR3QGKtooW+k/IiUSE
r1JCo6CPVNkrWdLjn6kaGryZE6mhd254fknf8HOF3X+U2WqstCh1JGWxs6+bmece
N3JBdQihYUCCXZOGAjkDNlsQkj+gEAFJEevMua/+xYUEh5MMOk7pKe6N2PtBaTDN
827l/3pk+kzLh8qQxFRSFLrSIL03SCA1nj7Klb97uJ6awy8Y17rltenUpQBrCw/z
Z87W8U/imAfYMiCPHfuUq+7RaKDsjYXxhJqnKAYahkpzs3DTwX2+m5g5aNmMaxqy
Z5f33vA6+7rjd7WNk7UkdRc1+X7QfMhZX97kwdfLrOoNHvfVdP/+PIxXEqYvFaos
ZB6SkITGLuxmmUOI+O0HiLoz+QARu23ql+3BnKnqxGCzrSjmc3sSsgbip2omELeA
Ul0cx/fbj+pxWNVWK0PyoAXl3Ch78QSvZG5YxKnVcbm7A2R2NLQHaswSi6h1VrLl
WrBV+IGpYXGQ6/XKkV1lbrMjOjDph1Bpci4crkVvAyd49q6C2bTtLHbkNR/kVpiq
65RcqDWoo8+QNSZ4Plb+zD6eRWrFg6Uwvevfuzg/uRZqMMGO2tYDl00cBGXya7w4
GxR07h95bMEyRXbQdxO7Rt6DEdTZCj+r2I6nmohG02XN6NV8IcmEfd4x1Qz4prnw
WfT0NHbK6a1ESTcmDreoMl59GvFWMM2cQV+8WsVBnD3UzNHPENmX7/FA8A23oViQ
pLNKXVmvuwjUP70ym/TZfFBiBcA3Vxii376nLhk0fEEDL+KkfCXQ4KI4rEDu5KeH
YWegICOGyUrQxFvuyRQh3lbWZSrQk8BqPodYO8V987Zb/LTdZrVwKjvSbLHTHyJy
s856rpRz2DNX4f47n3EcIVj4jEs68lBHKDZHRpxKoqVexg6QFJJBPRA0ikuBEdVP
2S4BAJv9UAbL008frjM9Qi6O/cJVqFX9/f84PbkyDJCVUxjOkqGF6yiFUbJj+Cvl
5YNDs6QqcTlgPU/uzaHPlAOp3EqxCKELqBNSlOjasvNiI1LXgJDoDlwYxzbvU1J4
mnLA4QP3jwKLMPRnTAIsbKsEqjxKxsGHbvL8NAXg4ry0Oc60JFpWcQxxD3HK4L9u
1yhnll8UBEDj/2NI501gkkRqmY6w4Rj8H3ximgWBbT71MrIZuF0dTYInC6s1uJX1
6DP5TO1HixUxs62CsSc3BUGh4/zLJBw38dEBP42UYwC1jdPVoKApkeE3oRiFasAm
zYGd26FmJbTNMAXNLpx1Y1LmghotTbU3HIj3PGPxnBcUtj5T9CuSMBAWJU1Akef3
TYKAdOFj651igUYjksKxOtvU8JLqllJH80SxS8UtYYe6BmZ+qFGMg1YaogNP5oNq
VZuBHPsEwjpzXLz6mFjpVVK6o3YS9hVAdz273Ar+ntrwXRRsf3JfQM8m3xRQzJqH
m7Bop6n+1iGa7G40tZEe2dVzxWsymlmGAee37RP/qxZKC2DNlXNEbSdg3MUbPWm7
ee0rwQbqXZoYZLsyYVuP+W7LRpC0eTAYJjbu6BJpZDcebJp4ce3mCpwDp7VvkF/1
KkGy5krN4wAURGZ/RNjFom6/cbU/sK0UlI9xmWHP2kYwrD4uCuAy8tnDEcOsXhnR
Eg4yIXAPMYPUlMmhDl+DKDYtdmR6TBEVVQ0IIHQF+leVKUoYu6CqcGnY16692eG4
trTkVODuEad36vuEiI5tRtRWSd0sieZf9UK/F3e917EsJzXyodyoko8LeIUKuSvG
in9R8RKDM44jzQhf9B08j9QQKbMBSjoHtJa/4HLnbsLzf0qnWfWmknm+mBlW4JWl
QfWN974lUfVSNVf/A/RXR6M9JAFwYbxCf6RWGYazUlZ0guPsqmWyfbpxoVtEktsh
BpO12LyVy16OVXwlxDbMLeJp13DCGBDUH/HwHDRhiyFl7YzvCEWW4KZEMipmoJdC
InlqlFYGGM0EpgaRg3y+8dxOZzzPNwCcOtl7ba3f8F6b9WY9YaHz+jNvgWbpln9D
kwku9IX0LztOqTlXEougtPjtUS+2BK/b8U33iY9nIIyVt7XSa4fykKIB/iCj5dEt
WsJfnr0dol6y49BZr1oskxCJo/HXVCgXCriPwP2lR3IHY9us+i0tIormbfxh1484
hIz8gDq59bbPnC5rtgeZz/pXSg0A76zsXL5ok4F8t/K8NvQv9EXZKw7uKLaNJYct
JijoIrvai0mOtpmljtgiDiY2TfkKZPB45yRjUwXjVg8q6UJeGJTdXFIwHd2f1A7N
`pragma protect end_protected
