// Copyright (C) 2017 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1.2
// ALTERA_TIMESTAMP:Thu Jan 19 05:43:28 PST 2017
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
nDFgI7vC5fuKp3n6ve2/1Kdg05//Z0EtGi5klMIu0xGCqWuBj2QRCdsjeFyO9AB+
EJ8ZCCkGykcGARga5iYezmMDtGHiQ4DoVy0SvUV4HbPcfexU40DJ1ugo+46o49PY
KKyts0j4zH/yw9TtnIIeKtdYKFQ0UOTZ4+QKDxkoanI=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 37216)
8/8aonjHsSNlxICiMbhu1NjXNm5H/8oj2yO5R0t1DMRP9H91sz1rRwOmhTqNh6qh
kFHZHF2/UDbe0k6USFEf7UXTLfSY7URrOBCMd9Ci7TN7LB2z2m4FW1xoHwG1SHp/
N/nN1whVXWtvEcINUTCtsTuxfJPEAlhV/pDtcv89PFsg4LxcHeXF/pyr9CDDU6gI
vXyZCDXS87lJ/CI894bisUe16Csh6+zWlJRyVwQUeH74/JjobxVlcamNl2R/UfW2
KgYsNvWbXt048k7Cvrml7FIbz16V6XGWwQn9O/yQbV/7jzvaDg+z2DXjMPSJusge
HPtYYFYF1OmZ1We6Vpmv4C7MT/C9BeAtLsqeRz2qmHVHKlRg+v8NHxgdGN7UC+EZ
a26UG9mLbFZrTjhaig4fXYX+m3Sumju1M4DfcKG0ltrMMlcKeVfuTNEhNk2Kmoij
buxCEmtnGYneOJHzLTqx+1+eI7dOtBGSzixdGZDfz+zp25gV0HUIykV7h96A1swz
TUXqHORHgj2luYAuhCVqqrtiCD0WqevYXkzlfHJKVd4TBWUVbFlkuEyLCXeHIKWW
FoD/XBK+eG2cunnd2X2igjQy3RNXlPN2lBVKB0kIEsD35JpxUNUa89BMtcbZgUVB
HL2hsliIvpzlMLgt5O4W9JNmPBbAjscJSEiT+nSanlyWPq6b6hh4R9JEEywtwr3u
Cfq25j2A24z2MGM9BVxOXYS2uPjOd2laLS+pfrePEfzfXci/zRZPxwyW2aU7gQj0
nLM4PXYC+X0Z0MjipxVsOmcuLrr20ZwjAeiQ7/0NukPCUqNtBn+ohqjRq2XvXFjV
A8tb7rD9ChufA/iGIqT7wYliBlwu3z1bGl2MpVxnmtSbX3Mz4Wu8pr/8uScWBqgn
j2W1OhVGBw5LmM8TWuilRW2Lx54gklX823xLK4fJ16uNDI7MXEM7IXFbWitWbgJu
XZH4C262NFY9NW30yAwtNswHlNK1FQ+3ihFqsmKoYgx9S4l0+soyIIVRBvBg+heV
InZtPb+3tgWYx7h3dYDfe5PClK3dCfQxUnP28TT0gWw/HSRYinW0iKTERFhN5jR4
9g9SsL+HUSYLb6qLqmLYQI20Lj0HqtXN8RN5ahJU6wBHsnNNYPncuoXKy/OQ9ymu
SyQYShMQb9ALPiP2bpN3Vsq0P0l1GCBnUWD9mwlGvvKDERobHhkA8jAr6ikQm9td
5yuPFugOxdba4POFrEaw0I5qoLcNY4xcmS84yOVEaLeIbRJaqgZt4NGecIo94dTd
lAhQJPtdJ+hnkPIokWBuIie2V+ZInWcwXn24UfRLIq7zLB7EHQmvxnB1ouEBhNf0
FuYpgTUMsv+JhQA6PiXT1BWwxsLjXYXiM/gBctbf5ouTXbXVvc112/b3LXLxHVue
gzvPLJx90wnUxH79zjG1EJ0FfqMS1S91vp+PWueNwX7J+kEXnkN+lL6uSpiCM2Be
syBdt2vz2RqqUHFSYttlw8DAQZ8SZSp1cwL+2Zh9duYrkXlvm97q0pYPjyuItwkH
MLMS9k+7Alk3ZRQrb8sClFEx01rtueDYCZJJaN7NkZhD1pIui6jtB0o/VYAv/FoE
i6y4aPMJTuR47Y+veJyo1Fqqyt9ECJSVLyNsAsrSjjTkIuKFnxQiZ8W0veUN4+oL
N96XNWnPddRCFDyAxbq4YJ8X/uIbTJRtb7vIkgkKXPZcz2DNvwWvtBrxN1ti+Rp9
xq3PP2dZ1TqqyUPHrWSczRWO8AY/cAGbbHcL7kqaIfFitIkVyb/WG+01qIg0OzQJ
irXbuxNb51VteKlnZ2ygsTsRqZeNC/rtsmkEg/71p5//vPhhchrXbN1a69YPAbwT
OWum5WWjJBYNEwB+W/uJNxnjSBn33gWi80mJ16oCc+QAt4mQwTFJHijHbh1FmEX2
tOAuO9BOPCZAgeanhsQftEwik7sXeL5UXP09kUV32sHwRNkGGWpwCBSGoY0TJfE/
KFcUFALNtSzypSHWGq0Z/uGZxlaUzWvynn0c4mpG86EBfkHyIoTYfUgwEdvlFwYV
AoOxfMsZxpvP9zQ83seepYfKXpJs54b73uCKmi/3N2GybPfPtsru0VGHfXoSDRLK
6pi8M71xuwgH8eHOPtgjAeVskgjAIwY9CSDUDMMs7bOfTtPje8b77FERDvu91pyC
sk/AjdpPuv3v/nGSDswzE3x/lcMe3ZmtSwxD80Lw3hcQriDWTg69R7zmc8qfSEEF
clzP/+CfFF0dIsyYzLaXnR0idlGHhIXWx7tJj7jZF689WUYpl+dkvZ4tK+7mkQ2c
cKsJ/bHoDYKzf6h7plrPYkv5JADaKPxruQEGt8MF0oVXXqvAvkmzkkAeVpw4NNIB
lp6t+XjyyK0jtdHNYrwHZqfMf3maYStURGnjHss1ktLSgm4ByhlhovU1lCE/7o66
4kjlsr0m2mZicP1CyKwq13OHmgiN0od0yhWEkq7Nr4UchTepDZdVUR+aQayTez49
8A5ZAbsap7uC1vR50jEpjKE/mIWsshLttC+kPA5PXeg+viOZAy/DUNnNozOEF5CF
IrVd+awGo5UmFoczJYJoAPGDwvnFuPJOMZb4IMttXVJAdwYQhGWpjltN2WnhqvAC
9rUZRp7nq1qj1VhuYsU427yMm6l8xiOptomUjIFBFR7QdTk/eDc45RPxWPj5BQ3M
pEnCIZt1nJ9cF/kG5f/QlLY4HsXe6M6MhUe0V4oMSjOm7tEksO9tQ7BUP/PdcMkS
Zt4GLJjiL5PN0xu+4n/GMKtRtgSoAOO4roNSHlZ1Pg2KFjhHFUG256hd104KlN8g
QJJvg52gdBWOD3AFi8g35XYERx690h5TJr7T5IVuXFnj0uDJVnrNGJx5J/PJTOH9
7HasW3gmz94t82AqbSajQbTblOX3mraldLT0iIUBc2pP9o/GaGLZAIrPCDtLqQ3+
b+i4/w30I7LwMhoVnphj50FT4rO6ZgltMJZ0GVE2VJurdIfnunMzPK75IIwWkKLl
a7zo6xMBgvcWb0LjdYcYe/pdvyXq/kcSqbFb0gpVdHE9Rkap0LYWhsG3daifyCH7
PVw4G1v1H+/kErhXJOFmAoKo88e+VI82zO+eZ50MhxRypzx9ksAzCfAxiirqPO+Z
dzueYRBANSrEEtRWC/ZsMXxenrjZnIBZZMg5jHY0U56aMWeuXgSQRj2YdnetfloB
kQmPle1yJEMYAeTNsamZqFtnxSmFzgeL0dDPvpOvLkRvAHBfxaNoEoiS4skE0yLP
JBP+mzRmNqd2fCsenjzXnvoYC+Aep6S2JEdzC0nDTCYtT7XUcVYlmpmExoZRayVh
ci12P98DKx3EqWwDlvgppbRf+uNfqV9w+17kpXUY6rIlrX5sbX2PDLSXOOIx9AHZ
uKLj1t+0JEvy/FUtasdC3HJSX3oXvymSDjaALEUfr8xJr/MLyd3WjfTjS2PGxzDL
6+DBl4aWggMkkFRDkfvErnuTkzw80Ku+3gJ3V2ZxkI4tQcJPXtWhqtR4j0o2y3+S
oDivcSkrfOQq7XTKbRATrIGqOMsrK7ziFZK73CEcOgrF4AfTRo/aKVF5QKbnoQPY
4MQRfRN6RGZEOLYpbKhlehbtK6Xroux8w3Qrk4FwKTLFuJxu6OE5eAi73kHwxnmF
JJTQ6+6n0Da3EsY5vz5CIvFb7T/yD5qv8tWG1Zuj20DR1Z7MTeEboUw3DThdOulC
lWZrSNb4IJ3L3mlHpEzDsOGavZBobCF1GkqapQYLzPeaGZFXMSW/ffC29Bz3kmG1
ejRBRr7MHLB0k8+SqH+N5lLcY900ZdqLAZmtSflFGRNTxCVryDHw3LJiQCPnANpf
hTArnDJK5wAoXNJ3kSYv6avTFg1peoVa090k7iiaxHOA1/qTKa7+OgqfypUeTwOy
+8tGjLKPg0B9BMSFtzafklETWqiFHeJpfaxruJcCGZoxUP8FbK743Ps3B3JI0tlD
Ro5b1V8f18Ul1LGKJeot1Q2fE6McBthbjdyWyyqC+Nlg9R9rYzh9XNoNztjJZSh5
mJKuTu9/txU3JravXRg5cwGzFKLatCUZhF9i4ulz+G5AsvPEO0efHC5788Aj0OhK
WrHNs99iIrRbCpgRKKQXzlcU0q0Gh/Fu8PmRSALcuc9Voo3Bf/UHbTEd1hu4Bx8e
E0tKivpI8cVPZtuEmIhos9MrLDjANr2kPceVUMmVKvdq6lO+GIGfYUefkEtjxgLK
mqI4++nQKCko33Pw9DNmA+3be4xHuYcLtLjQDTZOFh3+6OrceN6fvRLYetZaDOuY
2zByCXuvMjNu7gEnugedRC0Pq30pJ5uQmqY17p/DInyLxpXPoSLaWGxG6JQxsjD8
nxqJb5TUoMQPLGNBBFAJbUTIKaA7l5WMW6S+mb4R7GVU2NSvxU3+93q2oY+Q4sIO
pekkiwlDctcDOE3J4N8D6IJR3g3nxwDVEpNWX/FFyiMeNPK5OrLl5971q8SGm1+Y
xkTXamc74XGm3Og4Qt9FOcCRWWyJkmBn7gj/iMxmow+OI4tnHfFdeu64z6e6hb0x
dsxYjV5FnRRbYXjowHMuxdnRxLfq5tupc1XofcWjIjOo/aahRcqORBN4NwfcGGrh
GnESObqrt9Rkx36SCIezVHwqD7wRHE42et4UnWlkZTwKfSfBcvyrfJvIAUiLPWG4
r8V+FlMP/O1a+/aiE+pBUGv+8E62zMAQz/uZkK/NwcEysJsRYe2hrj80U7kucXpi
69ZrRhe3Pn/98X/SIjDWk8cxzh6vuS9WUGOOoURmmf2mV1uUg5fnWepVlEgO9Jc7
YdktmOrtwdfzUa22P8jK+gdCcfY0Tm2rDKoIxpYOBT6UrHjOb3E7vwPuN8nY9P+9
pWS3XgbhiH6U2pZ2D46wRtdnAqDrM3t603C3WdOC43rT1Rb79U+Vj22aLda3Q7iy
L1rAiaB5W7OsQmRRjzoEbNNiW0ESU0878srG6I60H70Heane5cHYbE5opnSyuWI9
XI3wftrAPAlR/g0PEnfyZSckWkXGv4ifUkW2FmNFNhn6T4tf5a2/BBTSiMck2CnQ
9/9xsIkXD7YOSzsQ4x3fH8RK1z4am2t2JcEGabxjFYnX87aWygMQ0Rn6pgQhDcG4
tbwhLFKaDFlOmdrvctD3CVkm60qErtbUjQv4Jf4HNShBUedGyhkUz2ZPtwZXkIm9
MKqACpy81EpMSTHuIse20feDajlH6kI9+8FEAQziK+cCfaK9LqYJ+PECNWoN4yPW
RY60L1JVdqPyR2MAtYmCPGk0Iiu3K5rg/SQQ6ZTQkJH4tj6VVTnKNVJWKoKXhMKo
6Lcgw6HgBoosMrFLaaHYGv+QRhntb1oANMLMauM1XIw2xDMFTCfLEthZYSvzWj4t
XrvF7R/lG2E7XXSpUPDbpL/YAi8H0vpeRUIPXh1YUgT3cyIQ1qLYWA1xKzHBfXLZ
S+aqrtem3UVN8LTe9UywcBMFZdM3YEAzcjqqfDAUqP7M81Lg3ACMvZQ+DlUNXDZc
XZL2kWGuwLi5+NeQc8G9liGzTBkBle9sUfK+Jf8FAtSxl9enYy1TeVHOGrDRkkGk
ZC2fTK0pueRClvgAAhSHbMDKZedWvRjw8pXA7Q3hhPiyqoiGGWQuunBJf6wpIYNQ
hlFgobrQ2vX2D3H1hGI3CKtlnihmy2nQ6atDd5b0nvtMeorMa0SB+5uqsTT5ciAH
Pv4HpqFoV25nFbyI9mhlCrse4hYgMjeEVtZ2YlGw6lWK4ahbN8r16zC0NK4FPiHl
jZSUPbifCUjKJFncNW2gfnwJNWBztNIgudSg4koNGwNq4R25ncP12jCH6rqy8Vn9
3z7hzlVaBZ55bda14yZK/GZZJzKa/6F0sMzV746ciA/HaT4/uj4HxZIfh0oFsyfT
3xK4swDYtylEq5Sbw79L27Mo3orBaLjej7wqpQRUduHk6wuYVdp6GmaqKvMeC3be
KmN8qKlv/l5bTqCTGRLBxn/6unDEvNI1RMs68Gk5Z0z6FuN0tVh/aPVObEvPQ8vO
ewT65xMP/Myid2dfRSAGjVIgmsYXyOaHpNkemvSV/cHR1L5twC2tWnqWdY/IMcDi
uuijSaqKcn2bFpTceKVehKvJkJiS4Od9VW9VFILlZvew9X7SmBjpnaCP/9s3MAMR
aLINuaqdQ/7rishr57WXWpXwdKj0OtQij/7yk+OEOFZS3hhKoqFR/WC+o5wz4i/t
vtCRWI60UvJcIEpHXBdzjVIvyqQ9uUWm3vmzIlWrDML1D1q/L812C/yFiKfQFWpO
Twd26Ll86cPoN8GMJkK/wVt4aLSXpT7Rl+HeC9HzeQMFcmphFqNqkGlZ/xpQJCj0
bI9aHiKY5KZf3zoVz+Bl8hFyBjRG6qpXZsLIAzOO2v7rcfBPRczF53MUW/lUPuZ9
m4xCkt0xW4JZwm9xIP+LDyeGXYU9VuB7TL/OqNvn6/n5/6LXF5cNtIrzR4+ga+SS
U5vxNxD9PF1hLxCihUQdg69M74lp9oxWOVTe0br+0zEp06vjwz05pPxZI1bRc2vH
vmyKEpHKtvSSNkgEo03LEggMhnFfbEE2aEb0a+QaW5hyeoFKbPM/xyVFe31f+vOn
7Jt+DDlcFGotfuLXAHT4uWAQ/ibUCdnNqwohjZ9wQEnfxowe6qSBm8P92uMQr/TS
s3ZMTI63RxQfvuWt5QM/25lKr/lVhuf+1IW8dfmXXCIvX01UN+gaDet4c4MRGvpd
P/9ok30IEPhiHMO1Yyh5hJP3hMfgHDk21GvAmDnBn6v3Ejmq1jh7WGm3jm9F6PaR
FTiQct4apo12QVqSxa1S27KHjlauRnDSl7IjZ2xRqJu/w//n/r7bPrwsRnwBwdFN
0s5ntXbz8u5sKI1krjqd/0iQQL/brNiBfgsJ1YfsJsS96YrfiH2QSObn3NzX6XWK
hcv2Qty7+hwxfGUb/qT7pM4ZzfAfVM/Ss+1UWG3+EYJsmLqM+9rM1mxmII1G1IZD
IOJxSBOFM9lS3ZqeeO0ffyrN5rA5P3rsg5SzbgrYVvJ/84vidR53WG/nCb9R/PBL
kyrFvR0l/bm2JOQVxjK/w0usnECiOXHKLFgK7fj+84jKq4ck2d76Z5SqYFD9S5LX
aEhg6IS/22ZTkwXUgiLXOgvC8pm3QAg0/F2qI1DCPqPHQ+jBeHvzf0v8E1gr8RLY
5RseM8EPdcfWCXEyns4jy1NaXSSSoqfJBhO/Yx6MEM6mXZpH96UBNmt/PlhmDfvt
2hB2drFZVcn+/A5ubeV95l49QKChT2n2qVklk0OvPPCsz3KvrRlqWOzIfST1bivb
KVGpNoNPSwd3kuK06EqTm1Yrt4lBQhtBxytfP085bSn+c1Gqbvbix+dMEuiY1pD1
yZJqhWrWgaBAP0a3sVzuiBQZZ2oFWUoWovhr2jyjo8U5b9ku8SG6BsARFYh1ocSd
aaD7IEcQdOt79Qt4T4cYIZCqqHf4eWENn6biQgroR+d2CLCaauyK2uoQSXfLu+pd
sm51q3tXjjSg7agwLmQIv1Gmw+1RQi5wHiNU6YSwC2uMoDBsUIN5htJf4yu/NurQ
qu2FbuGuKQ4eafOdbnxHiJ4STt14pmt4l4b4iStNocykoHT0vLOF1J6LIhpY30Fl
GnqbqBYWCiTD/x+mh7/7D9vRICpOgR/Lk9lpoj6tNpWhPvpgWUNsntDkRwbZdLJb
Le8eVCcAPhVU35mgaYSE+u14G2jdTHDgGbHX5Dvc0bcJe0owUHbmiZY3mvPd7FgB
l6cvqLAiNpZgdea51f3BHtyqdAlUt1labsB8yswj9CFXYmyq0+j7qaZ2pOxbnwBb
0dbcX86jIB3uhPrTRyTFpTqFk+2iFQv6O9ThgahddiaEV1d3coP1w0WgVtiTrxUE
kUbGS+CNz1HXa+rbtDoRIAiAFjTg9MJ1xUWrg0NkEJeM2pnsxe3slRa7HSyjK/vl
7XSXM8+2uMA1DWRHFw/FSiijBm1KudX/EydfXAHJwiwvKlhTzZkHx7+yOxn0gF0U
zOMsCXQkkXsrnPoXkO8CUwbS9MseAlFc02TsO2R5m2BGIw9y6ZvNig18h8Uz9lmv
9tgCsmI7vS9lS3XeWh5Gg2LGqbimblj6znHIlUid8TVRkdh2SB4Tasnn+R6T6uwB
uG/F+ZmZEKALQt1ilb0b3aKZUi761SiN1xEh7pEhaMRTzPPdhDNL935YdBj7oDpI
cehSzHD5jo9BlbZIDACApZpnm7WPsZNMHwxKFfaM6bUhgAoW9uN/dwYZOOFlrJ+V
IgYWBWGw+sGwghNhTQOi4Aw8IhGAVcbfN3nuu5Ac+wgnSSpp0/0wqS29LP45smKX
rtyQO7272bdv/3fdjHgS7Wnt/89lCNAr9LGkSRqGH8BdHuBmdm6wxST8Ueb6mofc
WRyggf9+h+6vkqkNzlvbpyQNHc57pMZU3EL5ZYM1F2WnosMHuuBzdU8Xe+F39tUC
FWCm4xSpUE89Qbz/yhEpeUGuV0XWIwdLXRzXGLbbwmdTyLJa39p92mB6zznYCBxn
/6psYHrGSfPiTThs+BDVnAPAPfnNkYZpE9GQoNME0TSQWNuUGPAJH3lxW/ZPDpyS
uF06WTwnhwXWsynvou59NfBO60SC4NGtBOcQF81irkikt9qBjsRuSykq+aKcXFho
fAq5wnM5M5jBYa6mf1I3e5eEIqg11G44RVV69p9hFjHNLdBjCTsj15oPWz/cdydq
3qk9W/MaRjPXDeK6GPk400R1IoHjKP2+OaLiK2/2KGQMo3gbvTJthbwSa6KwCTOQ
duDAf6RgP+EwvxSfFYSTG1gj0+LgnN7fxmlhBSzzZbSEKY2eVTBg9hiHOMdP3Wrs
sc9KBL+yhVmG5dG77E6dfE1ZMZPkfk4rq9DgNkEK3wO4VGmWdpr578Od7P0X1Dd/
UfHR4rUj3briKQ4TgkycRNPuncTxw6cb3d6amE511G13r/qdUhLVNQ6D4DbSSJoE
SjnpVKX02jpNzXlgremy1rgMJl89Bx976F3SdU1pKQiTH5B3ggL8Oe6LKVA6SW7q
lg8p2u31ZAWGFV8Bqt4t2LrsO/l2rohOpv3g6xPt7NurJPHlZQTpoPkBLW9uyEE4
aZmQwMHUagBSRayHk++eoJQrn55wm7f4ugbZACR6aw+O2W8AbslhrDRj4jaxfCLM
Ryd2o0e3E2/4MAEP0vU7fBANNQOyYAs0dX14RqRDxNNj8G6MCQgEvMidyiL3H9dn
v371tbrTXt7D5jeguzBjHcH4MKA0ugOarTgckZa5GsK1ZBveH+d9qT8V96ZPxxtK
gwWzuuv52LOKKKBIVjqLNXppbuVI8zvzRVoj3R/SDjEdFiueyVusiDjaSkAwNt1K
Gb81eP4ezUTAVfoIx+D2KipKZHIj0nchado0CERL7yczKjdmAGXHsjK05PfWitFR
yuKPLg+f8uIX1yMeT4SybMMQz803Q2omXuoXWbjm9Z+ZttE3WdYJtd9f1nSyRAy3
J5Y6yeKN5AmAkuj8MfI0bgvqHsWKmL8NmL3ZbZgupY/2pJdIaJn3ePvCk2rpbWie
hESRbV0BevnNMPT6T5rkpfvdoYiEJ4zQ44Q3ZMieCObUHICbP2Zx2Uq3gq3nTk9R
kFHJrVIqp9FvQDWd5oKPc/BV7iWebXqNUWiWJVJL8ZoZ+053G4PVGLtij6Sh0PHz
UzbBWVkseD4mxK+R7Ok/3kEGg/HgHJzC2Vkpy+QvKCOSRumGJw/gIF6dl7zev7dN
xg9obn9aU3EAM40+QkccRb01BlzSU4Un49m4IJYsyLPu4gC6n3YWxJcYupxwnnwX
S9Iyg2OzaofpXT5UG78f0/jNZl1asSF8gKlHKey2/QiJRiRDpo7fmws426z1lm2v
WouHrZ8ZS2a4VAYDVkAxL0plDoEGXcNFHUCWOU/AatkTTOjpEu52MjZ3ve1Raodp
C1W+rGD0HB1jq7zFehZp2pAters6VWiqKVpWg11JO9wrQAFX+dAdo2rr3Cgtx0ZS
Rlz2dnjKPw7CrTdft3glX1Fj3H/UdtWfWiEH3m7HdxWOtbU17G3/v/8xPnU40ALf
Qj7NyLYk62PYxcU6a1dcFZueMeUeu7hmIYmXDU7/v5tGhy7JvMe9jPtYQxXViL00
x5UZhTdo0mf53bNcHkRWq651FI461XbuZmkI+JVP1NWZmhSWOXoWiLc+/qcuAuvs
jhnQUsH2oIZQq8hoysfMKNJCMngQMjTH6IFmdGPlkkSH3Oy7T0w5Umljz0wi8Uvr
SsNIkv+dX8oLos3oxl/ASm9dqQ8giE5SC/vCan7ZtnNEt105HyOr1ejOm48ty2HG
e1dAFcRtO2ZRqVwDDEytAm+DGleFqnzTTQEMHD6aHHOTMQj8FC+14luzfxGfSVg5
wGyY+vDVpQQ6bm+wmAnw/t4zE5+ejpnz1aUnZ6Ct24klMWWJvlzU/G/MLA2KfFn5
f6ssCPmA/Puoe4S3RsWafJOn2+U/cMygr6x+FejmMP1+Httpg7GAwWuFewI6G3bO
h1Ve0sOcusDMr2CKJljCMo2AeugoD8WsLYSzVun2igD7zyfCN1kRzDOar3n1UnaY
yydCVk7TGXu0kCNA4uiSKa0iQ/U1dsJrGnFffA1AdYqNz2MVTtON8KY0TDAs82Qf
sgOnQn183WGwQ3oE0fMj3+X4c1efuParapWr2Wxsz7Wc3JNyZUIH5phkrvl3389b
55Xnk5tRUPzaEWSy/bMMHDkXt7NgTsoVfmLwcSN+BcJTyKUmuE42BCSSYLhe67Hy
O2Qpxz/h8VUimgjiGfsND188olyMz2X17MFyg1U8orkjt7d9EMPilnsFUbQ87dd6
HkhldgPczI8+SRhW2+IHEZ8Ys1dnH5f8cdsAEyPl05Un6+JDzT2g0QU2I/6hQBla
xbZen72Tb6s3iVfHziwjLXi4gl8bv8bc+IC8eLoks/Wmd96HOInE8Hvzl1ArFjv1
stZt4SibVpLVE8GKV/EuWTLptHr0YJYsOVJHcm3fTvl0vNQp/st9rNp3766qcB+X
VuDBiY3EoqqUaQigHo3xzQNNVwoA/rc+Gy4IcifBCDCjh69lI9vpAgWra5vpVUnT
zUTwrr68Kkq7ifFEOXMMbBIHaYw2x4CadbEh7YP367J+TYc8RUGAeZDd+1uKZMIz
k2rdn2pcmdpFnpXwlpY4a0tZX6aKIYpOXTBGvyuFrkUtIiBN+PW9hlV6YaoE7nRy
9l7ZPfHLkpViD+FVEzu5U6ftVi194mXcMLwDLPOPZO5YP88o/QFsNWjNBpYYwwfY
4TMn3ByKZEodXhjDIBQntqLrRSsoFoc/7oQU29h/Gw9pOF7W0NSBQQP4pGd00x+S
HgczmEeZO7pwa8K2a1Z51QJNngXLSoyKh8EDczxxwHjD2c7aePkiGDnUplRoHwWG
KxlXdZn70ENgAkbMjcjJEwwZs9p6beVWMnndsQFLq7+2FOnGm0JAK34J67ORpLER
Nm68grn51ah9mU9gtgRXcKC1v0OzWVLKMVVDgTC2aF+gQ26l0JEpHJuPbxS1DvbO
3CJMW/cY6BFON4mv2zAob7g1MiApiQECNPRqWJiqdiH39LIFmp2XEMaLY2gKZ4Zx
koIQUIGPULAkGEu1EGcVtdsMbEriJp7Znc1O7MZ8dG6CYJGLWaGH/R1LoXHNAelf
Viy9/0WCgFlFeDsOt51Qg/GY9i507k3hfz75pPYLJlcY0yhCQfmGAG7JEVWWjAM7
NV/JKBRYTh+w+LPkfhcndjIipuAzwK4bWCj431cy18rFy0iou44hNMLuWBHjzSO3
+/7/LzG1KHsREkoiOEtONwa8NykLM06kZYsm41tS7bX6cz9qw2NTvFfTYp8rJw3y
UeHYIU2mQI22MjF/I3sd8gWdpF2b7/O+RVyW28BcBvxVBp5834aJK55kQw3FrA6H
9pBij4gY3PvC0OXu63sYvIWjp0qmjExBM7N2YDldUkFZktWDGL7S+ZGen1xZQ+KY
tGbgqK7PdtyyqmDU6kfI73fHb5odBwWQx1m2hIBNnDdrLfLaAtx71zAQWTAMavNw
wIOelglsgOLRMj6iZSEF5xlyYDqtPfeoS/IPmMYbtABBCsOuXNtgMCJ5y1cKaJfH
kdlTK7+b7Qqez3Pz2DPk/07HdRsYXhO4zLk+MNnqqq4O0XxqNV4ZQE7dSAWSSuz5
wX9dljPKWd18/Wr+7heLA+0tTrq0c42ZERsn3yFNRt9Qaq+UW05hzYdoLY+FGZ0J
IuIBHUVLtAwJCZr5HjjcfwuywuOBlmAo7LyfO7kK9Rc0/pupvY1288cKB3dFOsLj
VvXJiB89n5Qr4nke3wlMis7SAwJOPUm47fRzjXtQJzHl8vyD+Tj7LuvhVUSQ/UgA
AbfH/oekz9o6uQQUbvrhjYLOy+zsvxTCg55XiMtg9DmCVrpr2maUxNB6WFp5pWwG
Oq00W0ch+pU/HXhSrLmI4X2XP013Ts+DRbU+jKq9N+lsoaeU9vb9w3A9p0t+Z8xl
zCPFInLsBYk6TEVJ7009ZUytx/EhCIxwXeaPzt4xXHfc4m2Q2rN1QhLsHGQ/DkTb
g/16+dxbpCbDkLFmD1XTYiPV+5rtE0RxtJ+vXdcuSG+nD5xsW+uJAN80x+QpYj2F
kh801VptGVL9qG5kwbZtNSk3VQkMKy/dUFpNV0Pov34AnmmTZJFJLEfY/GZ1W87R
vgh6z1uenl2IJFY1oX7H66MopsH+48BIoT8RKM7aZ2ShgLYuDjgEHelltA/rLkLH
UIAL68AruPuMSbcQJ6XfXH/tfKH9uasNWu9OWPsYXZaFf8e17zceV9IXD5pzjbiA
tii5t3ZOhpGG8cD7YdWn0qyJ6xtFc3WUpfE4nKSbaU+pbJijJPchXjgj9tpJCIKm
8We3t0duQ1rp6ciju8f/DDfqTKcJ05NhjoEqSnkB/5l78M09RU9cILF7bs7dDWXO
TPQRkN9+MMa4ONfZRYrUgA8+I0L4EuK7+KEM+NyMLTrrgSWmE4TDEfr5SXBQ6GVp
AeofhYQynR6X5uY9MOCgTJ1W3gTw6JDabjw+YiVzo5nMSK3Y703viSgIx6i1L7iS
SXjv/BKmkWm0TNDu2StG/+QXxuKNTh387mO2aD+HdkMHpjd/M3/5VCS0+64LONuZ
HpOn/Jg2YYwLneBs/IOMrOCOPaxFqfM1TtbyPz8dYmaIzrDXiZ9SgQiupXSC34XL
qko5eTo0amMD32xPs06Sf8ZPsLBI/d94mis93IM57McHvAqQiuQ5CFv9b4HFckvh
2G5fJij2qHSfO6z9nmwT3EZCDGFICDpURGI3vl17xRJqKUsp1ZqeF2jn0LpOZD9w
04nnVLr6+0dPI5r47Pyk158zyBKA9gxpvyZ0dlXtQtw+QxNEywHexQD5kbcMVtTl
XMCtYCX1VVa5cPTlVmzX01tOaChoI5MP7rStbvgh3kcgc2VC95zMas7NahmnGYqs
5a/VfLREM5NhYsh2YCXu9/4Y8bytpvwRQe0hiGvfNmK607vGdNx13v+/zeKweYOE
eLURgJYIeotHenZ/447UlQ/WKAZ35hFVDRUDFpM7xhE958GNP7hxZQ/DF0OuKJ6c
c9Ys95LN512eW+DTLO/aHhSiiUs2cETtnm4RgLDTvsdQvQrL+uQ668uUmJQ5IxfX
ghc5e+3bVaw92LXj8jOGjdgKNjvWfQd98natrDkL0OLd4cvYC8iI/mpPriGjVPRs
qAGrQ6EdSEnc9HDKHFi23SlAogdalhuerm7c9PMbW9Q4164JZALYNiy6ScAtCadx
GotjzUNcdsTuXC4s3cRtsnzKI7MVPt/hQ7cgVP9cTu+Vbi+maQ13ft2udexYODe/
QV3OxrSOi4IoKmvwe+DktatiCGBAch0XZU8aahMr3t6Zd2aed22Dyl35lk5WK/0f
/nJ3xrXepwEMAq0vDG4aQgQ3U5iih0/4q8Ap7yBgDRgfpu2jPlFNamUCmBgcYJOG
Syi9xtXHEz8mJUEtqdqvC2XHzrgDLVt3QyE1hLlZmCKGYbP3b+ZYRx1M5oDkNNXV
A5mbVht6DeEcplMpil2k3w1JZs5x7aiTem4GSldFG3IIt0B7/HxqyMTZ0SX48LSn
ilBjx4vw+Z65PTU152Wl0JzhUctkZTU8OPc4ktInbqAdQ3cfWTpkSQORxNTEFiZM
0yL9YJbOPfn37J1MoZ8sMI19vWd5gn6JORWKvXKp/m6RrwiZiLAhqWiZM4aMqwTz
WOCUF5TD8iVTDXR8sxyYWwSRLIWE1cc4UvMLmFFfYFqzwNq2ij/2NNGGr+e+kL1Z
tnir59lCcanFXnFHRuKPsuBDO7CVbKbovBObI7eBiajsuK8K0z0ZY6tibvbaAC1Q
Ug9VX4pHpjEeGESgv7QO7dsL0ApoUbbueKIdtBd9bvt8LhLoE4zK6FLgFKqVjp9G
ZIzRfhslRYqiPiZjNHuo+jb2ATgedAUTGgPatC4XfoobBL56LuZdbctsmzcmFstp
m32rJgiVLzakD+QlAH2surC1VCVHM+4FW8W/1YZ1OJIf7grF4Yu2uD3121gwkBsF
TxbJzCRFNT8fM7RehZt88ljZTPAIkPBFVuPu7h/jh9ZS/Ih+opLk4W0WKo/tmKRF
c+HM6/lzuDWA+y+gZWaa/Qj+RtkS4b4mrYTARkR7fTimBomJS17tB3JRkHrYSUTh
+jGVDNdlnUTeLsMa03IlzyGzv9HVn8MtIL3xFwjXHlRnByJN7ogeBh4vJELGvrg/
G3tcOvb1P0e4EFjAvts+8g/XYls+s5P5wvJUDBMfGkbKDfSfjvqdijs0gJOJjLr1
R7WH3Uzrw1YDh5kSnjPPgykPnExvcZwdyXeKfoQI32NCjFhn0mU/WzXASLqvZyB3
sqx7Vv2V28n5QtO/sc9BMhaPMhNzFzuPRJQG5xZ+tp3p0ST5egjQjDVdSlt4DtsP
LxmyxQqroaDj8F9LeFtLA5/jjXpqVbHM+hVaRbBaxLjxL5ikCVpYCxra/RFTdMGE
2T3zpMPGzj8PeZAwJh53mmToaCSgtLKHKE0PtjHp4QBvlKYCBTVQJBEdMzDYCsAe
4x75glYobLdIw1gH9NGnZXgCVXOERdnf45RBKe9cEkPb3I+ScZD6k7Qiy5cDJ1sz
pI+y54v9G97h8jasljZzaxWC/r2VikKUbh0bSU3mYMrE1xZUT3rzyv8em4SSP3MB
aaVCcB0BlBK0uWs1oTKDnrsRSqqfgpDSs3F3esV7ZucLN8KMplLPIfKX5z4EqV3M
q3BRypPGU8TUTonrcsSjY67m7eqiUBCKXdf3XhljY+Xhi96U2MtmnFBF1YuNJg48
3IzTKvo1fiB8BS/WFVDL/yZg8lLXYncQ2NC5asYwL5fZ6Ia+P6qJcjCu3dMrtKhj
wy2Jq0FBE5vrjhWNoztrSOgDw46YwDkymWre/JuLNF47S+VKyw5O6XJ9Km6q3AT6
29/e+2L+EMBZpMN5/bovIst9dzz+jobIj+uJ5nxh0t15FEziOlf3KIh+JxG5BHsj
4ABL01B2gOAjvDFwNUNgG6qR1kvvo+2l5tISKKvqRK/n65VO725PxblMyBtGJVfZ
gY/ktE+gFHVMUaJ7JdV0BFq59BuPPy3FfsOE39+chnvo7UGPogmzjoPnhMdNZ0+/
47mLXwgAiVsVxR1CmPPLMHsiX6iNch2aCE9qLBz0X/5prNf5IKZGwyafcbGWWbS1
M6E5plTrxNTJcmkyt+2xkWC086ZXWzUqYRQ6BRnBdA/VnzoSyt3LfqmjhTjeuEbH
xV0wUzidZEV+6Iu1lGGxOHSvIotNrR0ZR2uZb8gjAuu+zKjBg7itrzsTKwCiwGWp
GnLMKWsCk7846QA4ZfUdTRIv3QIm5qolNK4b3nNltg0DB0dRiwkhnDDZCc0LWdCm
lgy3UkirOZT8JsPs9hBvJiq2Hxid5mTq5KRLSC6dAOzArYmgqAIEGKGm2tqy3oLs
yu6zlSUx6fST/2Pw+4O2I1w1fwP4RJrDN1gJKJAbgAqwk/3HHXaSujsdlSK1KjRV
yq9T5WQqA5yV4srR9X2pd0qGLNcatESI9Eh2accHq+qRDWo4+kHzcmHsobP2SefT
S4eXW00LclsvLXJ/mgpik1ehDOd7VA7V5aXXenJ/iuAyw455EPQDjddwPwQu1qtc
ng6BSlr5fUU9MjuW4uHNUgDHsJdJHrOwORmNNg1tYo7X9o2JyffvCVmLgsgCeb1a
r3F0oVykgFL9jYspikcWHtrgTTZdm2FfVT39B/bKgVfNLig/MIF/NmQ/V7ROBv1q
f/CPaKeHiwrLxsjFgvkRrU+e+zaElm7Lb/bkb1UvhBs5Uq7KB+MreCuPgcM92xkX
wg4KluLzqK+/uiOtpyaWHkXiWg0QNeRZmTFY6/4F4MsZZ4xAl683tpuAoti7I0qt
PARdOV+IQ19EhooTHCqPFk1IO5yGsYPFf1MNt/kBxh4FBlDKqfPZGm+d6M3BLqUB
I+o7vnw0lXS9L1IcxnUoZ0vMXpYJU7HZ0M6MtgZCnApdsQ9otcgsE+Y9iiPmY4wv
Ly2HrNHY0WcN79XlgXsK5an+xkaHyAFL8i1NsmwhwFiX64e4TAUMh9pgL8qU/BqF
q4BPzEmR2WJwBozxLD+j04w7Bx4KDQuZiDrmBqMVTme/m56+T9GcvcPtazDLKdMc
btsL98/QKNt80FsR+CA5ngWbhb+TlyqqzNAOunredzc1KbUkXfJJoC4TwWofBy3q
XDjj8zrJK3vUY8Ti7E2J9Wj0GdHmlHciEMgN1ouJURkejdr7q+SH3LUgvAKkRLrN
OEd2yCU4PMVP3pmSwFiMVM/Z8QpowzfW0fxNjgRcgBjXHI7xZpTvB+VTp6qA5XOQ
7zNS4G067l+4NH86qUjKyhA/a7qShgSzc6VT4M8PItpQfa86ylmLQXv0pwC4WjaE
Ose0nes/p2Xk4Qm9O1qXm7i0eROgYB9ITGIu1rkf+I2wWkuh1y2JRcUVgFH36jEX
gbJss2cAO05R5cnJNRvgktuW0WQR6AHqA+wcJdHsTp7+CuFLKBj62SiWl5oeH1L5
51eSE6QX0ehzNMhUGcpn5gI9HDLIG1igzDK8B/R9MJstUS5pPqDJvgAySQIy+zyW
cxlJx20w4suGVTc9e8Zj2SJZtlttrgfSxuLeASOnGdsoSFIjg+Iawm8vRruBBxfL
oiBsf0n3poDMHr6eC8Gzo9yR39s5P994GH7/VqP86rg5wDsrycdyW3fp/353a5UM
C1ERaleSgc/UZHn9HCAZ0QRUDd8QCUd5/1+Gu4UXbS/aaewDWJeGHZFqs2CAhoiZ
QZew2mb+pcLIDqQDDEmcOA096K3NAK7P2FC15bYPZ1ajGf2aophRTrWFl9+iElMT
Leo0Pw0K8LUZfDX2ysUfil+cSOel6H12HJ1ZXgbjqDkTBj+FOLJRXlXL5kWzIw2Z
HPec1Jv8Djb9Cxh4Xiv3Edw8fr6oxuHZggqykd8v84ZN5NQPVd5QDgPHEKSa+ZS+
HJ5B8zi8qIC5RrsWK2zxjvZiEO57Hczs4Ep4sbddqCCy3bjwLNveqeo2fePbKrTh
lWjbNYHlf/VxFCA6RSS9nTGe/rmTOZ6DLb1FqeRwv/SfHHJvjy7hnMRXKAzTsNwb
SFewJ3eZEfX7YFs9UHhQxBEvJx9wYM910uUWH/SbmVh7BDxahgp1opuwX6AjMivk
15RFWxfGXVvNLIzQnuHW/sThtRMuP+WWC4GOWIeEdkUqUQk0dKb6iup9PXhA+Fxt
DSRGa8xAb0rtek4JwAB+9kaFJa+E8fDukJ60Nb3130KudDMn+xRMJQz3bdZnTDyS
eaupVwkb9kkMZZMHOf+Pqm32bpkUzCSA2/Gz4xFg+wTvD6i5U1Ka3MFeidNhfuZC
slHbMwRMofenDZ0eLwFM8Z0bvE7mzAnZnyBd8y987uapVGncVYUKxkbaIfFHpwOv
amki71jKmhDCiJ53Ql6ofrXsEZlDGykvm7YS3FN0AbeeRc3gXcmTUHfhD21CiXcG
RQGham+oUPrDOiFB52dcMzUtqW98MSpF3+xNpIiIvLp0hSLkZCCSrg4YpqStnvFH
XvXOxZwilxVoKm5+A+91WnGewW7l1waeh5cRI/GPktuzb4GoXAQQTYyX7mMKRI/x
fjjUO7/YAjjI6FwfzYtbEYGneqqx8xnSyMGCFetMOrr5hIFR3J/SSMZgRz6dPRS4
NX2Ysm00uiv8J8y7D42wWh5A9rG5pIdMJpdVulxAnlykPENggwFn9XvMsWtMdLIF
vpEdruQC710IMpOC+VZvAgqmoeOzCtBXCezeCeTlsDQioNQvssdiQOaQLKF+z5Ol
A9zrB8OvWnVwP399XFKeEVJYjBVAu3wqj+PZFoOAJ4G2UIvlxDLXJTqkpIUGokoP
Uobw1kkMFAuf67Ppb+3Aj7jUo4EX25pS8nNoSrT6TvqO5IghcX1iewvHzIMZtZCk
XD4m6hWCAEZPY0pKWChOD8AA0bmKLMAeOdUDRvVKE8D3chh5e+uoUgXN4bvuGrzH
NXPbwliDwslpMCu+DeteZ8sG50/QCUIL/PpiWSxHKLhs7Xmknaa+XML8dQVr1wme
pgEzADMev1mMgq1kbpKijdixtcKfjvxDeibqsWqqn1hu9THVGXIyfc/JXNQjW0aJ
739Phpo4EP4sX3MHp5rzjmTyrMfqKETgGrwdNGAL4jy8B88GmBTsR1VWReLosA4J
IDy1ZJFm/SA53ogXENoMDiyQbU4wHHERx2D7E3ZhZvtXTuHxbY/gD5k8Y/thxsJh
jbkWPW/JdDLqrr27dAahILNCNaGy5TFnGQSFgRZlzL0KWhHV0NO63YjRJLYmE/xG
LGb7tVNWqX6lJMJiuA+TnwXjZs3yQhrVuf0FWAzB+0VG6xyNkURT3qhzGzg9ihgd
CcqSbjlwgLzz/6gTmAh4U3KWnn4c3lOiJeKPunSn1BNtDY2qGYY5yTLpp/qJCDgI
TydoLZwOyuQcWvRRZ8z0icCLW+1CSaPdPTuVvmeLGMdp0bgrYQE/hEQx0HchIuJm
5JjAo/pDQWeQlAEEoX2Vc1ID1IBoTWJVonGdMODV/GB1jRmI/YUUyaZ2beguCPEY
X1tsYyvFs9+0hZUTP2DOPqPDzS2Yytf17J7I6bLX5VbUaWonxqgOkqoLAeUlGw7T
2spTmKGCsB/3K+BR/rDy3/A68BqiEvEUPy0feQ7ScGcjPn5BGtJFcN/f+fHi5bji
aDprSMq5IWjDNJgeZZOwcKt8rV7rx0pD6WMLR5UE0vjSiVR4Ngjb7xdpw4o16oLt
bKZ2FSzSCfAo6y7yVz+eJb2wrk8lfM6QhH8/kw7Q/UolTQQpoMId6wLQ1qOxfkAN
IC5NBkN17bwOiHr/rqlTLGq5Q41IH7o5PXSS2bCmyP9+yhM/ReGds/iwMBNeNQ9q
/tO4qyAxJ9DKWzlo/DYFYDh9upv7sh9G1AmG5oB7Ta6MHIAqupoQ1qnF6ASp5d5J
U9IO/Fvc5zDtEwxcALwpE9f6WSxokNUqTuwpnXkEgiKChB9YroV7BOJwZZZVDnWA
qf3z4GYnGOWPK+bmr03qRyNiMTuO4sq5xpIyOutGWQljZ8Yd15uPIu6ZuB18yXU7
ETvn4UMy90S9ltMDmME/dXHKMqXyJcNlJLloAUypHVhVup1O9FlsijikQY1GmSCB
iRfq2KQBNW1b/ZgA7bwv7Shxn+vRhlxTCNEDP8zSf0BN1BzWxkMeD7aifAMcFxfn
ICNt1XqDgUTeA/1yFtWBrfen6vr/r+raQWQdFwOHv9ghtwYNl6czoQ8Bkf3pcxiw
O+D+5mE4kTC1UatoqXtSowJ8fC3fcVGKvHQ86+/3VG54PfPqzxRKIaZwoV8h01Ah
lVy4PT5QYflungx1cBDySP8wIFU/7wUoX1NmHUyABJ5pIXx4N+prHeb9BSw8UKkl
FrUys28FjGOVCI4lg5qculUZ4hlJcYpywbIa/hlUUvJNEUDtfEDpB73UpM/VEbMg
tKVjG79uisXOEfhwhVCr+8TE8HlyzZvl3M2ygl4KVqMRHUNSyoE+i9LaE7ElbU0Y
ImI3O9F990eR/ZXqRU7s9ph+tLcDTLOMZGVmqd4cWrDzKF4ReT1HcRJdobGpGSAK
vZNJdA+icTBEJ5BFwCykMUBn8Sw64a6PxJPsHzWyB53zOl6LvKj0Hiu0vdGfTc3t
pZcusOf6NBkNgtWY7vzPjmjFDPcdK5CJ9PJL9qJSUzrDZKjRYjrgMUA9YKQrJUV8
mi7g1txMtU4pnWtu5I950LXp9QXsbwjoqp/2wfeIV5Uv8+n1jKzAaK0CDMR6c7ho
7yS1pGPwH2C3gmjksSh60iMqOV55cM66dlUGVttWNRt/xqGkAOhiO2gJmTbF3RGF
bAcUXPBfYEGeGHgH1QhevS9juEp0q2wXlQSeBbrprhj/+aCS0YFRbZ70ajhZqtF1
T7KRGL+24daUTZja8jB3juTTuhG0jL8z8GgMV+fVO31OAJH5yesjz/YdY5b4WGeP
ugyVnBnAiv1PuAG22pqFlCZTE1O0z+lUZz83TMbN6pF0AD6LwOa0FS/4ZOksNen7
GE9ibBw3cF4YYf3LrX48oCI+pSjyvm0yKI/zrK8F0XVX5G2tzIAptCkFktCNcN2T
bm1HhKZgPAPq4gVXZfVbBIslQ1hIwwUQFynjOp/M+88Xdp5Z2eB5mZdVAO7yvUQq
QwiWJdPryY79K+6jAQ80AfE0ga3hkQZhfQpMblNGfcdAuIu5P6d62eK3+gwhBW3r
qKcfScuK7takp07t+knzZC7vE1tWkm7f9m6liY0QAD1IQ9r7RoDJPfNIt3MkO7MP
b34+cYrUM5U6aFQFQR1Tl4aJUw9IfJgLMNdczyt83+3SXq34LwNQ4Fu0egNQd3C0
z3fwqXbEmIEDmtd01DpQIBbZeMsiCnYSdQd9Tc3BE+f6nNs11vGFYV50o4Wl7283
jhvZrsIfda73TiKAFixjP1fXw2V0kmcwNWZWm/SWRnJBtpN/mrDbHOIZCAD4rrZg
T060JHT/zp/Hw8gGeyCrFLpBVb6JuYjHJZgBKQbArwt9b/sPNZUQnXsw4YYhseYS
fcEff1k8WeuIMFr3aa4NcyF9ZlzcH1nEdZEU2Z+CvtYg3oi6//pV/hmEPy2mcq6I
Ucjf3ZKIyNNmGsllrVYdl3sVAR9u1zQDj6RKlYcoZ1pcjkZlB5mSjmnWStps1mJh
s7wLvqTZ7eSFCMzJmcub/OBuLbkMsPvfEETSll5C48vHh9k55NJeP9VxzmmDWyl7
E62DrjYmn5eGqjZx8kPycgKZqi1qIwFg1fcgB8H3l9t6GUQFg1clb2jjF1VIuzUU
SWo8zuGhZKgQ9H+UMQ4/auvIirepFFB4exhHLKIrXdrLfFM3xBxMntj68xXPhym+
qCWZdi35mTa1Fui/bt5ONCpwHZpIKvF0cuLiQsYn90a3IduPYGwrO1QGdtAcR+cG
vmxcZqVw/5Hc+B9MYMyuwmndzK/7d2UP5g9AWULf0RRTT2eoi8GwSww+p0bpDelu
DqzGE1yuBf8txKw49i8Bfh4LonxqtCAyeGaAT/K2M9YQnyh4o5Q/LAfaJ1WN7RZN
zU+U0pkm3zzUwjFqxSjAKNiovhxJvpLhd5XqkFmxaidu87Fwvch4SREJ0unyI6zJ
uisrLlBwpv+j69v3jpiRykXxNCE0qOlO8RLo5ttODG/tmGbJxXN6AzQsP7Lc6zqp
TdBZ1ZnBBd+qt7Ck+xfCohrznrc5lCFrjqXpMUOCC/7gQELvxd2Bu3zzrOKjG+1a
XegMGr6pU7O/24umVEx5p+7fmNt2qbxQ0pXXLT8bcRR73FS77WGQ3QVdQ6xYulX7
y24iMksDb2oKi6O0EjKI6Q7LTndlhkwynfeadN9NWykakNE7oyKstFSinb4jxLAS
kzMgtwrbhGpcUNMavrkgfBBEnCVAvh4kZXnApA+PUVuxy0BHXD+iZSlDOrQeDrl+
j5XxfRHQpb0rVIaDLZ9fMDI388YopZcroCmiVjsInpINF4fG7VmghoCl3iJ2+g8E
i6RNRekWe/vKZGoWQE9xdODc6vd/QbcNWX4BF3JQ1suw4B7fBBqutX5CpMmnuRmB
3DQd80P+cOPkwgZRWpnqBlpWJ/XNuhiZ6++LSSFBh6fmqT6gofbUgxK2VZkW/NY3
0fx52sGR421Uza2VHQVurPL8kYb+3AzeISfIa6Abajam9EIK0jqMCWJ7vI2Sec9n
Ib3BSVuxfyzH517ia7jL98ysm0hAJt4kVUNzwD/S0RTP5+7QZQQo2Xr0Jy9qfi3I
a623Gc5O3h9ckB2sW2Ei+nWkBT58P+JlRyIghs4mzxbc4OKzHav+0CrMHFNSsoBl
tp6ecq0VZ+O8jBwHOi9KkaaqsTt9jD21e0+VlqnoZ9oMWqXd0oU+Nou4CqLhzcMZ
FyTxY9QaA5vMeX58xlSA12XMSfgXKizY44zuvV5cMdF0MlX6Ze07fqJrj8+gSpAC
/1UmZHbYXns8Sagm/JH8va9JJIbXTUZ8WHFsPsGHJYZPYOmWcJr7CYk+4jekgCwF
/wE1SO+AlPSCLiqpIAO+QUWoBjt8DRUAQ+Ew1RPG12kOKC7HQrYvRfqiUoy2FNDU
Za5XyMSm8kSIonzgrEM1FyzzruVayL6x7l3O1tuA/R1HXUPgo6qq6ffNJmBGZgzP
7CBuAu64dhIsgutDaNAKNtHzubpOxoQKDnE74OAe0d5Gs+S+Sgegu/mAdBBFZkDH
R02rgm7h7ZmiZdvKtQUCC7wuC+kIDDJKeBjWosqooyX2HOk39Ynd85pr3Rv+tCHy
O0UiQ04QI3+hZeQBaV9stPwxdMHI2rh69LKwSLQwyInxXPh48I5LpmEwqlnybiL6
aht7fmhqdyioabhhL+BK/jBExPbApBRrJnl3Z18DcrTnTl7UMI7pAy2kL029yZk1
Bxv0pX2cgdFJXU099fVkgOXb9/Gd7xlZalydt2JofTOidz+Iq4Twd/QYLWv8RlNX
3arn2aJlV+ZapJy9BERLOW3SXrQh9ik/7zhvjytC+SaLVJjduEBiBrVoYIE6oiwZ
0edd/YcaWob8LgBQrJ62+pKkhsSz8qR3i9AeQcqTqLTmUKv1RjyAGnYPeKnQQjZW
3okmzBIGPLDPExQ+EGo6h5w/L5+ZV/UH7ZBB2A10Wcv7i25hMPP/ymEfqXAP69dL
48f6xhhr8m4diTI1Tw26hg0VHvwomF/FmNMPJhXhWPJboIN3AkFzSWxzplo7axnI
3+34X6nq0oKSxM7HoPW6Wv4O3NMMyD8jdUyw3I2h8/LDGTt0qL+ZBw08hPgkiZLe
SQtO2WN/W62eoFNKxBMPMoipY/0BBJP0rf1rNIB+JZsg3lN+GZhy6ab/fl5D8fLv
h8b34YySTyy4ZDkiD6RQ72I0XQB8rOc3LHfuW+g4koj41FO02KZFxu5Hd+300Jz9
ZLEIA7j1GG8bd1Dn+ziHCN6BLmaBktQivgfDB/ZP2bIjrARbVMYhdMqDYbC+SiQr
FbDq30/nRdrq3flEEVU9Qj11adqvecS+hfSIrKIPbYPw4FJHDgZnxpHd7x/x7NmX
iJJ/ATKjhaP/p9Y3ONEPC86tJ4/1HjFqi1XHGmJSEQn1WmUnR+1Atu7+8KWl0Zyf
8WsyuZX0kcqrDkCPLjAgj6m0ajZYP6al09zewdxT5n/L5U592SeQQSUH3jeQUBxC
8rnmXAiAZJu1UiCA/CZ+XuagD8FteiGWI31imVyYOZkmZZcTxRFU5hXdH0CBHpjO
t8i3kK7q1TZHNtmT5rtsYyFjRKmjTG/ZsrclQp8mi+EFUfBRmWe6xzf56MrkqZfL
GKeVl8vhv1/0T8lq6eqNGxeerORhCQr5eQHXzac8PpppISu04D784KqHqBcitz3C
RRJM2r60tyOhfq6wRpZFf/E8CR7AXToEpep+CIXxROUSK0YEYvHB6/7qppC0+ri8
mQRIoYLWLTwjsqOMCkPDKmv/F54S6ext4EW7ujlavu84lTCnkgpMAqbW36qIys2M
sZ3UYSxvnUEt5HZyJHT1TbQ5XK7f7Tlz1s1ao+sA6wbOoe8hv4CLuuMhjI8BbBZW
szMtA8XXaS2Y4ZcEK6l28YSin0Y87feyHvsIKykezWWfEyFsB6vRCxwXcp6Qrjgt
ivCuvLnp0GkUbzKn0PDaLUH/hJiTovtOT7l1qUBcm4/XPHvy0m3dA9tTKMunxpUV
WlNla+qVBrMUBvcUu6l70cRmju5v8m5WtZRvBQit3DkaNb5Ds4eYapRuZAzvSfnt
+zaVKL2/XBZ57BL7uKzdB/yk0pjruxBuGLC7xyhIWDT4QDbwtkgrV/PJUTxdKHVw
6pjcbbDv7FN2m1NRCG6sjkfeF+lMKYwDcCsRQXUtTGYrMGrKJbGlPrHEVrQSic37
FmclW5g6mWFZm2ianqp08ni79Si5cncBTPCVi6xDbWwXzlOYmYaSFlAxeQmRHV2Y
R7np9/nWgTu+3n2xQE361+v1wuRtgiXdlc9dBs68nGp9rt0LAT0mmisrJ9B9JCMl
ZcM95l7RQca2V8QCRnKVTGCGh64BnWOGSNqDivrbbTYbgIr9BneFnE+lQKfd4L9L
3EQ+4w9iNvDKoErf+wMjVnwMdUDSQZUBoSsrBtZ8X7iRnEbaNKa4Q9zXQIvgl0Yg
jgf1rnEUP7eLZM/cHfCCc3f8lP1ZaCK7v1ZlFcFU+24EyG5KhNb3eLTRdbmwgyr0
dwr8j/JIHPYRdU98Eue3jVIAGqkluR/HSpKjAw8rtOS0ALeiDh4lwfsjcX/BabLa
XAi2+4nQW+w0JuhxxGJbMZ5lfGMg1dXfKOxEYd97wuebCHNv8n/zOA2ZWNrokFK/
36iHj6KFr1lY6yOXBD4MFCSacT7lM/lGZqBDfn9m0rRkGLRlHilzoY1bNW2EpD5i
UuYCSJHHlh6S9hnGNJ7l6GOeLdt/eCRh71Tas/xOb3/Oep7CKkby2261EFJfXiOy
ILkyJd9ZolQOGJog3OgY+oy3d7rr5cfpKjTu/uJ2UtPqjDf07Bk9otE1dfe24vjb
jaFjrB142L9ePgq6RvCxZQssibhvn3OhYAfwASmfVQdfGsi7yFqcLvJKk75h4tp/
k2aca4+HYL7WE2oqF3SrduT1OfJ23q1wG1hEYQz2Gg85+KUKPoGj4G0Kr3ecRdaJ
Z5z8oAn6OxCWu6B+CzqpL6jkPWS1CFMM/WF/D4D1aRro1xx26fOzZiNlA6Po9Vqr
47dmk2kl+V4BW6QxPKfyVhjR4WEFH+Pfs6rC9zxOHBEO0wNyUOA/OBnvK5HX36+j
hm5I+krxRsMrNp0ZY3zNbpwYSvUO98SGQFjoqim48vs1EyMxqG8Rf4GT49YZ8Dw7
AY8mgnf6Lpj1HITn16tBaAJ3tk7IZypM/NJNtgzdl0pSGt3VlUcm+yvkPKr9Nl4c
OP557y5gNFl3UlViVHglZj249mDedlyrRltGRhHz0Ezbo5h7qUyM74I6NuzcOJ7/
HRJ7lP+5S3btPe5SwMjsPBxZ9n3+KZ5D+vuP+XGvZBafDjiBOOOpwGfrjpdil8SZ
W5WFND220CWtmi8lYkYR24hlbKPooqSezDWSozoU58XnJzaDF6pKOt7X0ZyZuu/k
AE1FiNQTs1YS11tToJtoLAJnNen4cUVP7G6zrQVN+vRhpXO6gvd4aPqvyfA5ozw9
GeOw/b6eFjzPgSyP8O64JLw5zCW3zS7DIXZ8MmmfNeIuMhZ1WI5e8vLsBcWCq3yQ
PSI4QxFqqxjPkwyn0gpO30IBfz81ye+5pOftnBLpRbcDGwnR54zivgNxFVWl4Lej
B7epKMi0hLntEC2jG262vdgoAgA8Q5AWSJmOq9IhF1N1i2Ak1IR2EMDUCmFRP40a
pIi9+zhwqsl/XCPCx3uNmyTknelEszTLaXXLcgPfUgjlIRcT+W+IusW7AY3WvCD3
carzg47L/+CcAAgrEOK6fGrbWOcAqzag7sFUPRHXyuG9Y82a85GFSugTosHS+hNL
jLAl/DZqLhxS0aZ/4WBgfXO/u4vyOTfbGKiWKrs9XV/Gs+dMSxLj1XbUPWBhnybE
ZtAAzHVgauA8wuTrLXpKMi2JTjVi5LtNnnMeNoLzgY2T8CHa7EyqODY5uJQBfw1f
rW6M0y/rFlw3yk4egTI9EeddAqzACtEi7vQ3vwbZsDwgvQ4vRUjh0iw+C+gLrs6j
Ljf/8e/H9VAcpQV8lVyBvZzv5/Jefh92KzawFPjYKd87unTVSBCP6mICLNeAHCGX
eaqPYGI6ExW3Y2tU6yHCL1TgZTgv/lhb0u+uY5O5G5GBzjrt4zDmBqRUm3XjWi0d
5gTtJggHXc3Cff6JeiMGJl9/qBJ3CNpeG4t8NFqgTa7sJSq6gdFElUCE6bZHvLN9
oMIKBGHmNJDoCEh3DPPObqeNVlGk+D849oBSz9UWN5DFTZeRSgGc+ZOkXGs2j8N9
fkFj+tmCdM3XeddfAIh6TviH24u9nI3Z54SSuBR9As2HTlBXPvWdGuG8N5uY1xtt
xTW0/CklKqAZs7iN0I83wudBAxOffr/QphhkEcK9cNqd99QOlWqgAk1OYEnScJXi
49+UP7s2h459tPH5U8yImbkosOqZ8XEIw3Gj4OkRGY6MyAXApsJxL3rMAgkuDvL9
LxWDZ2ZzVzEh2LcOgOURvBZsrM3J5omBu71xUUmaC5OAjW7GrG4HJz7GHZieQLD8
Ts60rW+dEYHw1P0yEYfbXIvJVXJYShyAatIG43GYC0sVSGIkw5tRSOmavUgJRbKj
0DjQGxgeXgB83zcV8pUnnWLBnRxprEKAHPcSbiEordKDnwY4l+O7SDUySW3N1wqB
4SXDCfuw5ZI8xIGWt2Of15Z8WRtzdsBrweyYO2ShWJAqqY8z/wkRYvI/dGsOCdgY
8y3/5c/mhXs8io3WHuuudZYX0KQPpIZC8kHajqmbUx+88CBvxGqpJuxuC+v37MX/
K4MBAt2tAHdsGRHPT98IGLgeaGmiCHbcoH3sjj6DNWcd9K60f4LsiQz6ihBriTql
VHIPBtGYQGMP0qwWl6wUHNDOff2Icd1RgZ7k+mpHsFEIshglo20xtdvvFXnmrWP1
tbz0cP0KHuaOD/eXuJ04YnPZ5smAirRoznVcoV7Ekb1CAsRK10dH+IP6k8pX7sd4
7gCGpx44nlz9FpccwcBlu1vvQKCLnSv+EkX7Sr9zxpCDQLDm+IC6oRO76SScIfIy
o7ivoWk2W2gr7HaiGPxXDZhNrlhL0Kal6GX6qNaKLvrcRtprXhHjJph6IP+eyH3K
knn218ZOS5jYCB7Bko2FYIuQ0RN88H+xh2eo2lBM37cVvFT38W+SljH9bOpo77g2
KR7PKkZLSMBKP6OPYc2WfdtBEXNhESPyefpQb6px4fCxcKPoUYhtWexFBtSQzDs1
N5hstDjGpcoxvmQ41TOTBKR10LNVbU1cK9dk1MQ1lVXOlUnfqN/n4duMbY82A7Zq
CzLLR1gemTKLBOlF4sJd0nuyoaXv6ksfwhnU0u3D2wZt/crHb6uLk8+KCH0f4z1X
C9Ir1uef2J92LW+IZ4hEMfzplvu9Z/bVhBoyg6OZ/gFGfjtlRrqDZNzNnniHUSrZ
RlA5fXmnM2LlDaQYXPjgLNHYXP2qeBO45tymO0cRmZWU6VLElF3bevyyfl4JBEox
k/yHMBnNx7zLhPkblHSgwMVzNZ2kxv3mD9n7FVIifIbWDYnijF975uaGhqAY44u8
c/c62MA0VzUO3kFJ6eiK2BblrqaPLXAk0SWfyekDxQox8ikbnXKvwQx4s5gNmW2j
07NKfloplrqHhNmq5K8XZo0h/1wF1q7qDtawWSiw1HF2pZ5i5bu9HEulyXu6U5eF
nY6hpuWs0TDx4X3HXU9aRB2pBeKU5j93vTOfX3H65Op+T5ESuYJM7V8KlBh9gHXn
6TjLp6FAhWy02/1sV16TdJ9mznfMnswHSHIEhRrjd9t5EUG4oArEl/kX0cYqWVMG
AuCI5FlxWjoPLABpXs1XQ7x7HvzKqoYC6ZDknJKZXZRiRlMYIxNZJvmDxMle0+Hs
RodOh9i+VuF0XwsGbFQV3goptXRWD0v6vbQ4nkgapz0N35/A2teZXf1uzsOKAw8w
JQzGSlbRrHOGWdo9jAJ56zEC0T78PAWFlm8F1IqKJWAJ6BzGVYy/jtBl5llJINfK
Chr2HBIb+NvAouvdN0FLU6fVxSaGPbEvq78/BHxD/iSxjfDUCCK7CKjS5E5/a1mi
fhgb1M7IZxIKLHtK1Ah6XAOOfb9NeDwcD0k87siq2M5/q5/EsIJgyP6LbSs5nMhX
TQM+koL/AxlOCtOPepPwWIhHI4dt3XFT8Gf5JrYlCZkcQa+NexJfVj00GRkHYkYG
agkLgqc9xWOPGrpbAZ9K8RZGwNHAHnva5GsN+N/PxVryzKqImZRiz9Q4kQUiluJz
yCrPuomJoy2LsQoHzGg0QvzxJDEXMV9xh6E/i9yiW9fYkd+ZTjpn0lNrGyxP/3vW
Z9FZHEaSQOyrTgjyGSWExqGNVbfiZcYt8vhviiHftVVnBrw4FtFZLnKhLcZmZ+Du
KaGsNs1MWGOtxwmMzOZPsowkMnOruzdTccegz+zsrZ0VvV8esHli1qCRlvd/sdXY
/X+tToFRJh0Hv6Qvr6e4TH0OT33jx5FLhsxbFp7m7CsQOKX++fYl0APWdLyXRpjc
fKmIPSSJzg1rulkD1sG7Lg3oXfOdyySF4I+ii1Porw9qFvLmPtafo4bRYhC038de
SOEULDuUkwZHx8pp41wBVG7j4EE5AAHUvozNBk/tGCbYyzOlwbhpDA7Z0207E5ox
bRjleoXsCRKqoAjJRHaPpStasT6GPKDlBa014aCWrEXHtf12FGc5LnZx609b2SO8
empM5wM5kNerryeU2icX/YwAHH3XLcF6Sx/l143H4VDZsIE0TozMo/En8LYXDGQN
eAKUjISlOwP3QKZk2xXTZkpTZy/LUFpPU5Muu0yWSCTYOLjPFrS3P8V6PK8XhXDu
dkRwUZIKuZx3vZw3ruiUvOfFZlwXbgVdI3pzHOQ63/IHX9aTliIg7MTmf8dInW7o
t2N4eCByzo2nAaQqRglflkIAg/VFbf5NMw3SXahJwG9szoGcHXkYswMqZZYNWGmG
zb8GinZh4CJRq/5iSZikIL2+fZa6gN/zgWx1NmoSkQBi2FOl4CnJYFNFKzuqxRuQ
WHnGq4s/zrYpzchEYxCBlWYOh5MAVoxeyakDJFhGJx7JdKMfh9prqa3canWeSk4q
hQHzBzfLCVdINBity7dQgLFhECoCq6V8hhGWDzwLvqD+Gz/AkYsyyqfmFqG59WUd
XZNFoNCb9cNMRhZeMD1yQHVsQVMm88yuH0xB2t+rqmIhNTnJ0Z7Cc8Y1kbX7XgAP
acvqST/t4zP1O2HzPSiOH1DX77h9nxnZCo+/Rzk5vnrDgE9hjukgU65cuUT4lnXA
FfhFr/HKHyMBgwr+hyBmQ3BFZCvCVmcgLZMwZpR78LuM2eFeMLyUSHwWbCH0Nelb
zGlU18PDXUdlW9cizZ5yTk8wfjQXDmWstbN/NobOB61OF9BIT5iVhbPTATbZsc6A
dma8zbU8KD+WlyXYnoDMcgUYhRjSvmclIVkpweRX4EJe2fyGAK2XMLQNtZkUf5Be
J56WN4+AUah42sgOropEPfXXmjYTUaK3vc4ssTz2z9Rpyt8X2LrmMK9AyT3SaNdz
DMYovhhfbqoiQAE14mwssXNtnH4DAWg69MXeocwu0Ib2PbwYhmsucJeez2w7qbNu
+zv0NdUNgTDSzGc1uQjsytAkkZDzvofFOwTZeO9pI0qiyPLDTDdAeWuUlo0zcfg3
PYWx3490s6Q7W3ruBkvBwOobvcxPpwzgBMuos8g/BEyr4gR5lVI82XzIG0sRuX+n
qd/2ij73+ri6C572OJmf8og97o/eft/RpGyjKMmw+K9fMoYzPGi+DGz+H1qXy8RQ
mNho8grsOT+mGX0OfT3Ulhwp+oAQY2OxncYV0+KvllF6ZShJAMU+gEwRTIRtR5kA
/H0nvoclR2aKVRjSEyE7tPGDeaw5SiY1tlZ3neMO9Xt82uFVqpQmXjs/+VS89+ix
vmjEZBZzgAXU11MNbR/AbS22l2yGA1En9keYwGpnjZfJ9g/fGtT2ypSeMql2zLTF
Ep7URQGM6ExJ+p6/3igplnLn8iGG/YwRx1E8JAVLCo+0kF0nR3iEyhNUNPPhsykp
aRjJXnUU9GEkaSrbYnjcc54MrKIwd/Yz4nZUE6UsdNzZ2KRJtdXpcx1+jQqOzAvG
iB8tNvFAhrsDc8QBR1YHSOz4edgb6a6fYOzVRYAhHMgPlqs1EdNPXvRRwfbI3fEk
7dxI4BrX8BVUNx219QCZYgGllwE2BjEIo/1aVYvp6nnNaBX6N0TfhyL6UH8w2maQ
XSRKCh1I4obz4q31+XhVktri5YhJT0miVJJhVUYCV+K7Q4cSZZ/wG7m+1yvrHMQJ
yEkUZ+I2jL0vy+DhT/dx/06IyeD4FQ36/bUtq4xAp5FdmBoK3E5+zxaRZiV15xpd
gawDE1nrA2aTQHRgTYNuwPZhbNCCsX6KSZ47XR/72CxgybUE/9kAi8yTyH7vozzE
pjIIAjmZafDC7k6WFIpr5Qc91jQ6H5XsAwhOkBq+AOpyt9ONpKZ53OzW30V95LG6
/f3iK3QcV1zIutnOgwW0hTWCwx34ojqMndsunAyBrRDKA+zyGurKwvLC0l8SKW4V
MxCXUEycnlNT16jtCNZx8kn5vnY0UYbC2kSzj9r7Q8a6Dy/T1iFA9jWDrS5Spl76
7XHVJxVgpihcwPv1uvip3g5op710KlZ0TJ0ovSLUH3a9gK4PafNaXep6AgFMgWpN
QMkQbqWnUTeHGhpDle+umRH6aZO+qAScWqTY35Bk/SmumA8YsXBQd1ETpcYw7mQp
4nmV4MsdMsdy92weCFF+jNZSo2oxlrFPN9pYeJEd6NBafcMNKX0ojQJKDFxae3yW
Ym11VgVb5VN2bpYHoqLcVqDdE+tJQV26J8VJH8lcWWrERQR6l/Qhw4XV2muwDZ++
VvTtv3+QpNF7XWIA9dvHEpG/sPUEP+/rUayn3DUzPrSwQDciZLP/rw7DdH+Gmipd
mYtu6XlDna01rwE44gVHNEQ3E+uMANqXDh3ICx5661e5croH/tL/Hr1U6kLLtIZk
+E3RSWpr4P0U71Yy/ctFwlg0nd9TDRpq4xJtP6qpO+9FWdYB/p/+dP38hfIIynNM
Rio7Uwf9rpsbCPVe809ifdgpIomAVEc2+6G5jm8r4IfyuM82Yo8otXy5tbuwi41e
H1KKyqKgD+RpiQPb0lXgP9iPGuhhL03gidnJqJjs4VIYYoDgjF1fiiORWGyDwwa4
nnlYnEZqCHzHdIAQeZxVRMFkL3irFDh5gdvdwyAQVvNQZHdNP7j5AYxxAMZc0SOu
LIQc2w0tsomPhmTCOwJeCoi9Y+SjP3WmTB8LVleWcwuAWZdNp6yuVXEvWkvjA5Rv
Xbw8JcWCvKh4MI1NL6+w/xYLUgduKMEUxvhmuqkQi6GUz+ueiJzQw0D08GcZjIPA
tr3s3PC+fPFwTu3V1rAoIlerbi7fzK+fMLmW1kSXYb/aIDVuh1GdzjVgunC+SOY1
Ts0BLekPiJmLpgVJBxtfpy6JZQwwzwMc5zvRiBO0XbPW1X5XAs4s+SQiT1O122tP
6s42U9f56kpNripUXJHZizORMWyHBIunRBoee14ZzjPcXmR0pwTPLBZobCYGpOth
jft0FqoNwoi+cAHxGx557NEgkWCvRA6EzRt0nZVlW1ERi07nf+RRDWzP7OwFyiCY
esGUIgBl68coHNsG12YeQtCxoLKQ1JRSTM1M6ZY7LtKa8G1yMp3Rb4YPMxZSXlSX
Y/tGhMMHbF1JHey2n0Ct6Rwoi+m7sKDRfMr+C41KR3TxuvQaJZWr2qq35gTgrorJ
Um16soitvBKVT24UEKtOB/ywc9TsbjmAZ9jkdQgczr3FNyMA1X5UztQ+OPKQKytc
fJ8mGV6pnf/QjAA/9XOvcFAa20jiryHNB0VsbC3EMWFTRdTtOXqZBnbVhBuFvgFm
izrzha0Xxds1FGhIIZT0h+ECEsb5V4gV+sqtrLd+r/ifrXPy2ccSGZg1T80PsdsI
sVmUta3PimEoy8pwalsu5AsYdQhYOO4p0pGdJ7LEDwgkctWsaYR1UVEd9HU6w3sL
oF3yhqctSIlKDrTRHsntY5BBpkly4shBRrd0xNLed4qzkdpCCK49IiOlp1VISLaM
Paplf6uWIB7GFl1JannX9bBmjTNOw887407PODjCnRf5PRwFUTshj+nOGI8Gw9V0
nqcVn3asGVeVfPrH91p1Q/dG9b8c/GHocIeSUn16gBlZjvKmUOnyvb9oHADNcwBE
UTZAg0iiko47BWZVhIp+WJo9iLUeGF7h2DvuDc55Ac9nad1FcLTL6jinxDrtpiaD
utRA2/sbaqrSXnMtZJhA5sLGtbxtsEt1mO350fOACXqOa/ylvJzeuMDeXxOkZncZ
0JRtgGrAyUGKVC/A/p9AGcjA37gDeOwbMA3eCOcLWUAju6OfWxOJHCboeALFmIuC
HC1JttmYDecTx3XOzDxmnwNn7N8i6Pq8sTbqKQ03I/LKIgTghN06jkMT54e8xjPE
77px+Z7v7aTKFlA0ZWQQRs8Tvew8bGiE+FgnB1haSbposo+KNuF+EpTBdA9h6RY3
d8dwT2XXyx1kHjyu7YiadhcO7yNc7iwmRCyaMyQIvQn0jiN1DQiiTq0CtJdYbHz8
OHV+XbOHWL64pEeFZcTK3fNx0lpuGuHXy5uvGPwm5a2dBSTUb9i4NSRdvkhhGh7Z
+vl6vQxrzEt/dVgVW2mPLGXSUnBew+vQTJSb0YK7skPXDtGFksZXgX8pLIE93d+C
Kljr8wah0ABMSs5XeH3benI1bUKTL5FC7YiUzzl+SGtNMWr9s0TnufZ3MIX1FoML
OqVIwyB4Iqx+O8oQuA9hmqxZphnnRN2M26bmuJdgr1Wis7AeyC2gx4IIxzN443zi
mqDr3GkkZyU8K+ZfEtyepQnfy3nSKhHH+tGnkLb7++XliIpvW2JIbpKFj4Kj/jvN
JaoUIpvo69YeDCosXKRALsoIbw1FcwxAxYEV3L7Fg/cxzXP5jEh5VuyVsTZ+Mu+t
Hg4l6mfbv2/TABFmaxuu1lv4ptEDmYKxy336u7avz3Uw1wDGHdNrOd2LRvLPFnT1
qdSQ+wgxDHWuGrX18REnRXM+5pv9WYXmYKf0iAbdc0Fb+5tjdswSD6IocyfhR2fP
48Y+fggW8pAdFwb0rR+3p97imhp+xoAYflqqPS5LGt0dmqRcFo/qpaQF3fHGyJlD
+sktR6FjKxOatyey7KR0Ch4ijMXluJyU5vBGuv8eVpRBDfCj6MVVqrrx/7O3oKDf
tSth66gtcQQo95DDshlO+cOjpiJScBZcy337+abkHnDgd/MVaIy6dT/QTx+2b6tA
R0UmuX64ptmOZiKrOOYWj1hfqRCVUDcb4qIt7vhVjkEju2+6nJGu+2oeoe14DSVz
wth+Y7FE4s0lRGwPYn8Tm1cZBrfGmc7qabExjKIZNHe0wP7Vck10mIPpFZ5++8hj
6JInXqEBdCZ/wQ+pzIctmBjrcvIOm0jWIR6tAB7MOKX9zFM86KaDkROphe4KX/Rq
LZo9wUWO6IcuSipDGTxb4sxgXr9FSa7LrbpNv9+/hQfmcaYG2Tyvyp+eX+S7eSlv
2pbs2Bc5veId4jQtg6zd5GA+qLnxaVzGKlfqepbyIYDCWiFN8Es+PbRlJAbJrkwm
gRUV3ySMQhFr3VDN5H2G2HWqefG3G5wL7NSv77JPnSqfcset+vXg4vBiFz+msUPQ
NPSiuAzOkUm/6JCNf/sUdB7wI0c5N5Ct8EZFW5jj7+RTs5fRQD+hK2bUFTtC+cvz
pddqBU1aJAQKiWfGpRx3V9nnR1LokRQBjG2Hom7bDtdfsgehubc6GSli2zadcidR
/gwIieZC03iTg0ioEpAWEZbnDBRGg0FxT+ljhwoPqep4woXsdT03/q4ytV8SVXyn
5uUY7mMAhzqqRtxDw6ucwiQ+zyEUFYLTojj2gb8Y1lIgenGhh1yDE+SL8K/Gi8Tu
FlV4J4Av07qBkoGjv/mfbHwS800OQ2XY+Ngb1ZHwkt4BCC9VpXnpDZ475PP91pt+
zFESSxu6vt7ZKhOwCh1eoUHcHchqOZjedpG15yQ6ZDgBj9bO8gmx/sabzhvmM/EF
Z0go2ZdePV3RCiVDJHWHAOfbkh44sO7H88lnKVCE0mUFk9h6OBWdpQPGMVTuZGKT
BVNzHaBRnkC8mG6SVyKB8GSvDVmfPzLPgKwktC3RLSmJPMVw6uvNn7pdv790kyxW
CCYkay+LNCt/KT6l7F2xLzlij3SRjLMib2kYcx6LfOmqHBRTlKVem42BRi8VnCBH
Ft2h3eyBq36QrDVWYlob/W6SaX49oo0a+yGoEnMz7+LgSU+bV32QuWkiSiPSdIMs
gJM3m6PjhcxB/b4pn8w11umishIpeX+95qIhMIdcLTf/4UkOEUmjivDrc9la9LlV
4/4U15/lTMluAQbHz/onbK4D4TZRpk+I7VYdBmgfypdQKQLmGkbUcpyW7Q2HhAxl
XEcX1bCBJFWzDh22VQLojpZk4Ooaf579xJdlvvOhI/5hA1ADEXKyiakEgqmHuVLE
WxhIwwJ1QHuXrGTzU1PSLJQV4r5YrVJ7sfQQDjONB/mP4Ky1PrJWbjZyvgeghwBU
qOOAFLWfvhmLMpxWWyUoiDZNfkkRUSC5msEPI2hqvrHvSrsYpMX9FKmUMRkB3Gp/
FaT7aL+y3wSO68Ii1OfrfZigX68xJVgviKJ6ElS/6pCPoDNv+8olfyK37Abpnu1M
4SH0g2oztxFCOAC01WGzH7gkwkNLh+jTlw59DCAFT9QiRBT25vxH3uL8vcLi543b
0GHL3ZKE8l74QDCrgimmUxk2xndlmplafuLYn14T6Vy4Zq83vzJe+b5TWhK7Rg5k
GLAX1GIO9Z8hlRMI3MP1udoKpFgBHZv76qTWDioYNB0pPWZBxp6vBz0l3JHSHv8P
HR5M/Cyurb5riQulXL0W0iyvZe3U2ZfKdCzdt4EF+2RReaKsqny3HOyFWbEs/VlG
Mj+Lq4Z8UnKGDWLFGRd7f4sGURsAHd7MVVvwXLD592Zqd8UEVs1qPur0hi606cCD
cstiNossy0v9rIoGgLHDj6a6MPex5o3gbOyL5D1h3azaUDCETmlShhVyB06f1jIa
HtVD+wPFlaTfieUok+pGmVQXY9g94uejIqTVjQ96nZISbX4RlRPPDNOvdDLCtYVC
5ZOnB7I422pAJyGo+8G6WTuVk0QOY12S8gcSE5CVyKNmzB5iOt++p5iCbUafTtPD
TacYgdncbD7dMg5PNRwj1jDemMZId6w6aCIvwNZo2sS1jajAd8xl/j17yguANOQk
Zwe0+oFdVznzmWkvykbJcPNQXIF5WnY2cuf4sjtAq+zH4wDRtdfAXoHuUxipKkQ/
grE/WImdgo1TEi3UXOsRXDssZGKSsZTw3HMPD2Lcbs3Lt681QeXMlXIw2R2CvKu1
GP6GuuW2D+UkOQHwhe9b18HMkquOTxMFG1ZUqKvQJy2ypqUzvyjYWahTB9wJfxL3
1aTtBX9vr9n8yXJTBiR+sQlsNynR4wOzU3baaiNea7zvIg4I97qBbASF9Up6xpea
mVn7S69ggT78ZkXP+dWvqK96D7W5rdKabnn2ndYxdqiRspXqqMdkLPmhpJ0iegjk
DHmHMlKxjEQzPV6r7OHn64f3nXqQA8BW3CbL5TfPyIeDsLVMB88ZNVkSQgqhlVCZ
wNuLKhGfaCMM/Nv9VeFl7PN0iM5KB4kJQMw4Kw8Qxfn3xTh6dwT9Una8MSTzJST4
CpNRHqkGF/NaY4L5HKy5Z/+N5a36AN+Jw8WhpOK9kgIJJsDwMzFdgLjlvAebiId2
Yhj85pb/519csWvVCjJJpESi8uHs9J7d0nNuKurKoWqvNgYfHu8QS3cggVAyr3a7
Sfqx1tkv9X3ExyDpj6W1QL9yxohX4dZeKYf2mdvKVFGLL02DD/DjMUGTFH0DLEuY
aItC5SktJ66UcqLHuoppfjknB3pa1nrb7s1aJo43VwDe5oDvPLS/OqXoFB7wxafT
xm/H9w6lyF0qfw3ggqCdUC+UlWulWGzBe8AtI17ZPmuuhwc2AzW/ptntYkMd7rTb
pGs+92ElfZiCkgW6IgnPNbxYpVvG3OLEfhY+egeu+5Oc8LdiI+lJl7obWk5GgTP2
dqdNI8WMrnityw8zXX4K1xoQefUHpgFKT/UqhBvb6yrWmECS2Kuifc39P7iNJ/YD
1C/Dmra7k6Zu+ZEJ/PHVOQntfQPIAtIEeECrdiXBPWNkqdDRgGH/YxNfmt/a20oX
Z2ED2Bdqn8ssJuc7G9Z2ogl+osIGCbPpDR45l3K/qLvxEcTU/DNHFz/inhDlNnBM
cV62cRb3waJsnr6SZBC335JT1AI3OmATrcmWMUH1Av0UMLbAg1D8vIoV8No7GJlf
7cZSdaEwdccJE122iPSroSjSp5+i93nIfIUUhntguGBmLi9GJKs0fRonzdnAWtHc
cpmDcfLUWzCoarWRNt+wygTP01tJ+nCbWBeQtx9huRwAqgjVZG0OucU2Rr5VoDP8
VknJ4PHJFbjALevx7QEJddFufgFZHSQOxcfFovdeWFSzTnPvN4OmuqLlsZmmbOGL
MLaEKNxqHY7zcTPZxNFaZ3+cqNAKptdd0VshgcjMjNCVtiNjvqSvkjnbuD1F7HbT
H4a61BIU7z7w20bNZmznh/kc210+ZjT6woNxyPARV+q98QfPKaeczwstOCskv1Vb
Sb5JOydCscw7Rzi7kKqgLu+WNLZkW3xpcUnnz/0lT3IBhUAR2M+2lI9XFjvjx+gT
VjX+4HT0C0fKfPsYTVXrvtZWMBOwWqyHmzaGPqSi/ao2hUhBHAyun1qM9064LEwE
yA1GRWwS8cYgYmPziL4sSMwCl0J6JkfjfnUBcAL3IZX4xalATrzUdA0VRMw4hTnG
853FNHSnjrSQQ/iwuTSdpEZiL3OBjdmX9u9aLykBXGSVWX7YoEPyYZ+F1tERWpxN
1mrUCfMCAz4riVf/zqGCsXVmDY2ENeFC8NTddzYTp6+mGpJZMPBDjW9BiZ/Mp4fM
p8me6KHUs6maC6KncG7ut3aJVVzTa8QbZskAiMP8/QQjryf4mikWVp8OFR7RmGmp
JrI35PPf2uCDe4cg8hhrRoYjP23H0VbqgpBYciELOt3DA2ypvGBVQFX38g73AUiM
gDoJENxsd7HTDttMDCuycHnI40KD/gnQPJ/iHkh/AOI9XesQ8JaYH0GvlUR80jBb
qlSbyD0bz1HF1iRHJHnkyRYE1rqwboZBgW//LptwiL/pFu7X/0tDQxYhG2TY/FeF
jDRDz/kZ6U7/qrZBcWpD55aZBd2faUW9SgFTJ4W4MKKI8kdqAiqDaeh/Qi62hqEy
rTWZrwmQAmDWquHNEgrcboIkr0EJ8tirKZdSPt9RCsgaaD449PpV9g9WtdbTYKgL
BJ26K7JnNqBTJDy22CV5v3fQwpo1r424dWHaRze0sJjDDCIF/gLgFdezyzGoemv2
brCLanojFEWaqyxXb8pR1z+aWaj1ejjkrZCbIFAoN5hMbBkwOVM6l2ooKPulE4Do
piWWDNDVr+Eu7UYSozDRWbq1aKuq/EaVewSHgqQBSE3l3DaVotuJv67Ey8nr6E1P
88WeHn9bZTGP2AzpbPIivTnMB6VjK4Vx6EPV4faBTSGpb7XTmI6tQgZriZ31HRYO
+SdsmSA6/o120J3wW8ycHLTv+4BE4HtqCODKAdfZid6E8b4F3l2Pl1bbX/gIqx5N
1ylE2PQY2G2ZDiXFIcrZHOKmIlARQX1F52uAMnZFAwSrykkddunnCTKFoe0Y8COC
dx+b52HjmPhYgTUprEdnjyNJhnX6nQp0MEZ7AjCitaiz93DOOvTyoXW0xA7ckoG7
Z3ftrRHvVadu+CLrMY7paK/pART9aILzsqGXraozH8knpga+8xt/qPgWNsNR5to0
KEnzHwjntT9GbMJqe3KBMQZQ+2oNWOGM6cbdEZohGkeQRx8RSJVSF+UyluBP1jWa
uh0F5ugBkICsxmkrX+t0D/Ntu+MxB3iGI2r4Fi/xHZMZlBaOBWVhZJwwBcPYfxTI
ma/cy7xP3+9HQSUDHuodOdpo9cPfoU9vfzwvjvga8+CH/KDQjt9uR0WrVRcdTyAx
pUBUD0gSycQ8lc/1fDnFivVi7ffBSftfWGkFd5PhHzTp4Bknqz01kJGOuvU4+k40
7zqHLPM3BOvbJUjOAwpFCdCfwZVOF/lTByWIb0kIlmcFpACTA6IdGm6PZm/Pczqb
Teo9hg4pFBj3rFxP6yXt6H4VvLbORm3RCBPV0cwQZihMIGhJN+Z3ZpbyMqER+NQ7
vVvGTx4X2UyskFwTf4CC3Kktnxv52wahx1+8xq75BzYfrXu1xWDFPYhsKjDmh0Nf
8Nkyl3S3EESP1I6S5qX2hohItGSCpwRiWaM7BOlqmD8FcM1wLPzvF8XXlJjohgGS
XAKzlEn4QHr9Zx7tnQoyvyG2p0+NwcDP0C1B0hMoSDkRHf+G3N9qjUFya5p9q1xN
FOP54xRZUkVsTAAd06bHmLkp4aMQZx2ODY7jGySTe3nPk5HvoPtsRuPa9uIo94df
Kx9BhkMb0DsUYNjvMsdoC7nc6WVyXZsVhbyVuRKXa3pCbqux6+trNP5+5jy5O7bh
jpui2PGUfK63uAnAxdM4OZA82iTEIB9dLVw6RfCU7kxhR3WxTKsbQ960cG2Z2u3r
zV4jsFCN35ZHk/MJGUdWZFUMs6OkT+vIS/W4KISlYMW4L6ovvq83YqD3xCPizv4k
MbGOJqgDUC4Zwq1OyTKol4sVaLh86fXcdMu/jDoVu7he4gpzC+2vD6GuxFE/3BMt
NGl04Z6NLOocYyPItGQihKAWA04C8dYwu7gQlQ0Z/ZgDzdvERpCHjQpxwmbbzfW+
BpWeCiP4Te4rSGLpfblR90ysBvRuhN0V24WuGUuKiCkeY2Lrg4vleaQnvjyjwvBe
iYzyd9F+G4cjXqvMgR7cDYHoFz+wA4m0WMoFSfYc1oqtMNKQ8kERyiDYAAZMwx6v
jTY1Xp2iduWvbnH7PyH4UeubNeAZAVC7gwimA5sAXFpaCYQTZE0LqRQ9O3nKlwef
AmKcYJx9H7hGIaR7GvZQKWv+FCui/a0oBKHnp+MIuid9JdwS1Yy0kQXpu2DD6OIc
Noev2wXiSgSsvuAQKAwbFZlRLHkub6sgpYaGeGbhcf/r8o1Nb86ko6Ptw2Y4x0Ku
/MG6AvxHrWPQt6AIiSYYp3gTPAr4kyei5k+LPT6poj/Fdi8DisMTYwWkxgfx7PDD
2SyiAMJZ6k0WG8RduE6IeMJKmEA4DTfl8l557lMpHQkQeAJsx1OiPia/SPWlJt2r
LaMEpSrIFrLwGBiqBVPqD3+pJ8jz1WAfVvNQ3isKXmjXp51/ISsO3GRcwa/XQadu
GTyAo5Nliv1P47KrjNOJfo2eFMcsrJFzuWvjZ8+LiYTsYDPT+dwMrt4UXM8J/Jva
n4fYvMrcirIWgog/+CjNnkKh+dLj1pTNm+jR4FvtgmYArJBJtIgUN3efQjczaF5h
ln74C49LqjJkdCLnO3tcNNdyHmMzDxba1NJrhxd+iKyqUV3Lj6rq+GcrmG4k0JHi
ccvejQzy5Rd3zYt6k7PQhxn09m0b+IBhHVbz7zlMllRp8IGYKr44HlnuiUsIOOP7
zypWdlMOBqPN3ovt1f+EnEOG1qlkZI9kc097d4ICBbJ82Tmfje8FqwQd33lVAx2W
YPHZnquJoUWx7iYnrvbwuDEYLyiRWmUtnwJECBfkdS9jgymDKYzV0fLkvP4A6UJi
sHS38pCZwkvrLPsWLw4/4IdaTLwEBnUWbJDF4e6E0HHdfZixSVoc7xt6dWyseGVr
Ep0fV1ZxYK60lUVDmKgz65G8C6rza2FMnDacxpvNm/4yQhmOpdgK5nXgYB+ZZwig
34xMue79WCOOz3zyYbO5WMz7g8DjdSbYPq+PbLSZtoo93vqFmhw6xO/1Yo6W1+Z+
5eQPLB7k1BJQD2/1IoKcLSb9iMMnxLaef3rJarfd6MMOSWBSSgZzf7BUYvKZvt9c
fmecmbAL/Gge6EBAMeAWvQ/T2xj9zL1vj2ttSILP4RU0La/ZeA9itJlJd4xg3RGJ
1rwQeX4YhjPh2p7C4934cRBzg+XgM6XwpnfAtCI/gIXOADWM6WYMknXg5pQkMlIQ
mtiJ3M1LcVrXbWU7dyuQwjT3rHliOcFyCrzFN2dRaMT9WjJWA+sJwuUwxXrc34uO
F49jR3zwEU5Yuadokr0hn7GlDdhZ4Ry43pBix05W5J+/0we8e4+wyXzx0+jGlyLz
T1/PE7dX8YJq0izUOZut9bQhUviR0G7yK5Wyc4/7gfrggqlttFToADQ2H3AVHEQU
O8PJ9rVxOeoQamriMTwdRxaO1TmQMQXCLG4o2OJE+DKb/xspdPBq/MWLYWalwwAP
Jp9CN3IqvzbGOhmC8mXoj0UDYInRqmFtNG051x8qJHmwgSfdk275iuHL+xY7TXrY
HSmOgLEj0IVDy7gChhlpxaQG3aY8PLiFMQEKwSltmOjfF0jPWEtEyDtSU+GHfLp7
iQ2UB0swG5e6Yd7WlYd3ilCbq1jPSkEUJeNfolGe/nJClc27wHZ04iVVx8fK/SAy
8ZXYPPQC+TEXErhI1TOXIF25ZJjJwKCap/JEsVc+ulAli8SGxiGJDoLy0SMlW6rs
mGtDrDz/MI3Jd3jtqjAbsK0dE21eyW+O+WxSR5o5K8Bx7T+Eqpc6FjtdM6yy8Jro
wPoHp6QcctvoWZeTQtwdYPtRpit7VI7feeHc9aJeZT67jAMwjD3eBkGkEc0HAnTO
omg7TizGHsbk5gXYRd8Jcpp85hXl3swdnt13AtgYysrZV4MTt5uvt5Ktf1aD6xtG
qIDjW+ZV813Hi35pCE+jXJlOE9cf8rB8gMVJ+Oi5bnlSnt5qQImRRijyGLuvZh9y
Aqr63Is1rKJADzw7Tvea+pmfA8LnNdGlEllg4EURKg/bzQGP3YTCiajdStq7Bh65
3VW+ql26smHVxLpHYnYkpQQyvdp0L4GxK+87dVLQFYxANCMziyj8Y+F3APh7fWp0
zEBXt5yMAyrgVnh78WIqRiJdQ4/l428UG7NGUdZlz/qNRr+tm5J5seVmOazFO8Wj
zoSURfHXdh10vXKvohLA8fzcfu4NRflmEqJnCaDNOZ2EmEXEF2gryygu0gEFpHne
wY9v5BSwrOng50F1o56HZG6Rv19iOTW0zX5HCdRVYbNs97ERaDAhQPULUoUsdGy/
AJaVcx9ZM42O2cHI/NipOvjDMLvwM+esBoDiEBORt7DIL3w2Drciu/2YnM+FxOxe
qdY8UEHzZQPeLNK5Wh8Axyfd127P60cGFmw4SZp71/tIrYeAF3trK+tnlmP7hTYv
GLubvIkRlZiIi3ks+pcuABoWlkJTBcO2zp7FoVCxyc1acJHK4T2KRO+G/XGsu77K
54b5rH0k1klB5xIkW3V1V/jQ/xzdRJjB1Wb9NtyMCASAG/4qTFKVLwihfLN1cmSM
CIcHkmZTr18/HSsqwHCyTykZ2kTOcGY9IaCY7mMvPh5LKN7TCOw7yqOIKDsldjsd
3ZPA6OrxomwWYDBO67CvDiT2JFg0s+9tJaOU1IGrVbXtP4hi8UbIBVTQCEQCt+Io
F205kMBpIXtMMWE+Ld6NVuJDwpuRfaTDOekMdWcoJUniceqV7YkEojfuLJhFE3/m
d3abRTJv+mQAviy3NO+d8Ya7SLB5yXBgq8jbnQlwQf8nLUgAYlwd03F5vIb07dX9
7sIwpKq/UcR4oLyFNqhJd1GaD6vULPwWyqygr1Ug0qtYDi7pkqUjLwTI6lv9ZyF8
yel4OIGZdr/gr/qiulWm0Bfg5kGY1gVyBmoE9z3z04kwqECS1jqS+sv4vFqoar7u
4gBctUHX0zILPUT7+XSYmBdMa2gX1yxWpObIloREkE75JdSFwUPJgD+LJx7ImWac
/zwwOfHv51XoHUp5Md+bJw/V+RUpQuSpjuQ6fdXii64A8Txt88Dz5IvHmJmDYbOT
5a2S/sN15/HavDban7FaLywk780y63Fo4cF5pwg18BZHCEciTtFgT7EcEoTLl+n/
xsDNgcUaDv9ZyckorGiNYR8IgtDWHMZbXFDZBzjhH5E1aRfANR3/smbIoV5Y6EM/
Sfjay+4QPMcntg1PpS6/D2cdhSx1kyARSIRGbFgohN4VzEMepH+fVfoPUjJWjIYM
4x6cjswY1ah9Q4ZpVqU22Jq7xm0+str4Fms9YNESwkjvDjlQbGc2S1TBRaR9RGm4
1eTSEhE0hWbj+KeoJnwMzzJh99g/kO/c8FbP4MeVO2F1h/aXRlVvA7xmKQaddt9/
O/yPxymxe4P2nz+TPnw23fv4pcGtqu8eTvgm68aQH6SiFoFRFcpMhZMA83v9tn1I
XrUOjuClgIDX00BxrSwNDnhD3aDXgcKRgCeM6eFJgCRvSIrQRzIydvMhFbg4xlCd
Bxq3W/am47/0HP45CA9MHonY/j2dqWWneXGthWdUqn8AgPOsEzbxYcZPFW5+53nO
FagoLGwYLxvIADQTjh4emcmpLO9eQBJsI8IuBK0MVvTkcsO9YWv5C8nAi/ffNHpO
fXxxOp0VjrijguXXYy8ZLq8W1Bbz/7GKv5L/fXKmWMnnG0p68UGIqbDUBx6u1fLa
8Rw4arQXdpa1benCtRyvlVlavtR7OtCC+C8N6ckS4b8tH8le6+Hktc0cG+1qnJ/F
u+XScWqMx1PFuAIMe0PkCctJaqsLj+aP+Iyxz+1Sqpj2r1ukvk6zJBJ6X2Pou1N+
fG+5NG7EDqwWBbWcd5TwLJIWwML1Lnk21ErNtaIg3lSkAWLngTNQiqLPwusRaN6M
UVzRzrWaccDCl6LfWkkmuXc3O3h1yGe8m9z+PhPz/WwsGhNF4BTG+UpMurfztD31
wWg0Ga1y6IIIK5NtnfU+IuupfWRlIwoHOp3w0SsSs+bNoIz/1LLKQfbyPAwrSljb
lBwnxUvOCM29vtyQDgyvwA7rvGX/OnQpS99LXMcRDb0izfPM8WSiHFTOnRRKvtNX
V0dKNqeYtkdNV3rxKM9562wFM9Q8ZeuWSseLEavTuFq4ySCRRI0qncRUyp80e7IB
u22MgavXKe7bTCCzprHyPFo8ecax3IHcc5UYXInVDU1xgOxKYa0L7owT5iabNfRp
C8ZsjdDneRm8hGwzEHDAfkaf3Twb/TeBWaxPnksIqiXoqgeVm6gLuci3fUgRZjFe
wHQ5wAWQrdLmlA9v1esWcfRobhCWpvgRK524qDQMkOlJSJUFhh9EkOAWQY8RYpwF
x2GH1DPiS1kYCTqzhpd7dAvxlBPXrbW9E2fHDaJDdCdlQGAB7IeBDINKkOPkMTz1
t7nV5mcmca2Mw+fCxiiM5fkFbxmhr+vjghwfgCo1r8cSxOwMw5qVTK3imIUSn9Up
c/UoJ8sSIWv/ygbRkFrCo6of+FirWgzzvfp/i3DZYXDZ2Tvm1tMxWWluuGPWlJHJ
idF/FaFWJGhnmRT+RsyR9atgFwoY9lBjVd86xFE8R6keLooZPdA5gBT4Ene7hkF7
qETJBOhEbq4vEdydNpg8Zz2RB594bSo2pEwNUUr3VpQM0tenuiKNN5V1uenDM7NA
K10+35drjcPRmid+FloTpnOwF2AIKgDGbDNXEciU32H545vY1gBLQEACBiVEfYqk
6LbtCjZEet1900z+nBNI4e+GnAhi3SeJZudCAoa4dVtMcZrkaHcZY5OwpoeBH4y9
OZAjb9rTsysByUzaKXTFqKkgMl/lmMnweJKW1Q9i6LsixXXxkX3mLWbfCt5fPoFh
rhSBCG3QZhiYH641zgkfKy4z/vp3on/Gb6JgIG/SyS6NfsRRYFquGgTAYgvpJWag
ryRn4mPhYifuVjqH/o7VegnRVlezl/O42xym+BDNmNltLtaQ7HFxqUuKtAw96hFe
Vb9YwKYpxBeaS5NS+GoaUKIIHde9evG/AlVfI6PY3RNAdRnpilnxkX9FGrtTIeId
Dt4irzY0kLxYdukGPSHN36sYnhtfIHrnRlf0gmWXJxMy0xC6m7/MLavANYpbKgys
IzdFtkQVD9q7vd58H1ggan10vCK82PEEwIDL3p0LJ8qyJwl6gWmb/ACnTjPCmcgT
QyNtx6ksRO/oRWUttDWllRpdHy2tPu/YlRGpopTP08dsNkusBPpYq++l2EzcPk90
3CGFsVWleFjauDbFicg5RxPo24F93YpoHUZHN9C2a2iDwG0RGZyx1huCzO5CKxi/
upXn89ioDLFhJjiS4uRhjA1vsTxJ3mS+pMBEOJEXb2HzO8FM8LcBpHFgl3inBjua
Jgr3h5UfJBe1gbmAWZf4u+QDIkXO33HB7UZpeD+Nuc4YFNHejhWyvROSZ94a/b3b
ZgXyMyImwiEqv4zUJqxOYtBi//Gq4dMPXbF8mVi4sErGjcxvCqB5pfcJYUuSa7sz
1YHQ/nuNNSJRbQTkD4Li5/PSZSnbRKxc6pIV3rQNPTadjd/Z1MZSnLEJT1Jdu0Gp
VI0AvCQQB0Zc+KnYWzOdBnFAHPHCNSAX1iDLmpz1bX2M4U14ZgXh4Xgfm77+15EZ
PkShBGXLjRyFfvEk5NKsVgkbxyP952vh6FZc09mViIlpgvUylLZJhFkshSi+WuPW
W8DfRA81nee43wRZTf38HL4xYFRCSo/+fidrySAKkzovH5vYLf+mnRC3R2zf53eo
/KeSyr/kirxVMgrhGpyjS2lhguc0Or3x91IK6wAuAEpuoIm9PmKluXmmrHJieUBN
3GlrwifXJGkyzcWEbLto/mCsJAC/ztPzbuGt8jG3FEg5m8oObeYRM4FtsfkwWUVt
tlRWt9v6+/7TcIUf/spip+fGI+jobE8Krg8MhtVz+1P8Mv7j3aaf4M3HV8li6MVw
KuNjklNXWE410ODDgwBUhbQ4/C7osiG8Lc3/oCf1QO7Pxyj1w4qT6FsCbEAVORvG
dPGN5wyWmS/lnCj8wPMFiZ7AQJtrKO518J/C1aqBYFmlsWMPlfMu76HxGZfr2VkR
HbwqV91qF/Nf6P2+HV/9ZqiIGgIqiekXGOMYT94xacvQfIuE1UzJRXzuPmOGFdvg
ANfyztQWgoZ7NZBEanDl8eRbZ4f2858n4LbNdGcENtBh9b31NiXW0X7gjXdHSM0E
53pnMl4YqtF27qqgaFAy67rxw70I+yx7Kn4SCJew/GKlOasSoNIbQSyNOlqVwV0u
o38+Y15MM8xvGF4cxrehecRFmhKKHb4EuQJyARiFlOk8zd4zlPDWZoPuys3iVYk0
vapqXCIUM4O5t5vKWzkaxgaf4+uTdHQu4dO7DHWP+am6hqzizZPm/yXcWk+/2v+2
vsCQmdb7avVNveoNmWx/wuOVlWlVy81OvvXdZKufPVPgdynPJTXattTtXNMJAvvt
f7RH7gyzhWCVTmoZuDisNAkbI/BUBwjksS5B6g2xcdlrdW+lZtOr802mwdmMc/xU
M/bYgoJHjT0BbPMUZsqQIuc7G0qQHV/JW1L9l8TUu7yZM2/MyQsFQd3A7DcNRAAG
6GtUu5wz5VQJVf9yYuSL/hZqxbP9l9D9jMeuBff/OIZ7bsYxw0GcK55G2smk09m+
t2bkoWs39KuUPaahgV/t564zmPxHNmM7k8yxCGJqaeH4m0ajIbgfaHF/S6xkZIIb
JYgwgnpaNGVK10Ibi3bnhFdQoAC1p9P7pseiWSLq8kBzFFukQ4sG/AsZOY4i4zZp
RbILUuonWR7HzrHTbJEbxKG/ni5mODAc9bzXL2kstPXsVsdYauE6Vcpe5fpeBN7U
YLMuAhvv+zplhZ/WLmp+DV5CzJzZb0g+jEnmyXMbwn+X1hcuNxfOsHIFFO+X/z5N
ooU5mJvlUlYb4Y83F9rI5nhWdGFXnBNeUGqDnWzzk+NkTdkurolg249ceGDIQeEb
UuM+85XoN3YlBlD2VQChwG2EfZqEajfEu7GCn5A5byxClmbKnft/A30y3t9kmz2R
uclLZZNUMoB27xURVjq5Fy3owT3rpcnVSbcyzSLgGf6Im5u7NN1A7+x5tnx93CcY
M4E2vquP+ZA6EJk4EvJS7xghL3NGhoUJMBPYIY23SQVjxTqo9LOJxnculfYXXYRC
oqp8xxL82vkh7CVIGiZO3eJA1y03yRUablOBk3446sPCoNsmvoUF19w07qj1AOki
CyvBs84giVsqcKo66BsHm80p5dokBRYbqyF6UXrMxKKZtXQKcJV3i50JYTmmVfQ2
igOOBJTWO9zqDcudpCc78X/x20qPPOiAPsMLxizGsspLQOEmZQYUx36XGVnuO6Wc
G7M7E85soIFu3QD12W++n7zrq3f7j3i1nsgMlVNPWOWEo7GoySRzlUV5+GAPRORd
wW3p1s7iRQh0t0M8rnkHDAYKWDnaPJc9glXKlPwQZFimAacRj4JWWzhoMzTqK7Em
/lVhhyRBnZpNHo1WqNflp0+I9GDb1fAjaIzCFQ5hDVNoPavFBPD5mfNoiFVQ8Yh/
MXcgQnPJuXHa7G32yRHFkFBV+V0FoEfsWwtLqcKRzmHTXzYVEvv2XUDA52IExjeM
7535FAmsF5FYt6+HcUA3+7PVJzOlj34u9eX10aeTpDdiPYjW+qw2CkrC04OVxIIS
mczO1qTuD/uj390OHhh93pTZCvgrTb91fBnaGOgTQuh4au57dWBxpH0Q7PoRWvxs
En1rKHxTszNO4urHn8liwj797Xra2R4gV9WP5OtdNl+LdQ7vkZWmAw8v2cycOFVB
LHvh5DblEGAriNYB94ZmZHAEDylx6XMMTi+N6ydNV4kCnsKo1pMemltHxegoPR5h
gDJs+bqIFucLyJQmGwiL4qWYIS0BI475WpWhNKaLLj6vzEotSGZLDn7vDszZg7Mn
fmg+EhBD3ZLyZ/5Eh+mcw1YWoE1NdWqRHFb1UtvQFlQUyoeBld9ya9zc68a3mXwk
fmT4/73thPQ1fnYHdapsVqft6g+950yBapamkcgL9we/U5I5PiaaILSjyl5k/pd/
wnctUyJmfaVVRb6BdV6v+2LV/L0X7S/kpld2NxcG5HUcwDRc5pRe4nLyy9phsEar
bp6YoYeXiJa5nuqgZPfw73kmMaqmjtJw54usRDyAhG4kgJbBoqO7+kUIl8qEFQWU
zSOgLhpEwwhWy55cL66Nt15Z7e90+416s0SMu2woeuyczPMHvT+lHBdD2ssxetnh
kk0R2yRiqVj8Dhdp7N3PFshoelK7vELdMG/q2wwGY7x9O4yLRa86F0wXK4PVv5Tx
R6PdjMHq8GLjOeIz1WP/LSdVvUrpPSelNJ1wluewyODyTK4jv9uN5A0bDFCINaSv
ml7ORiYWgUlxRdBfZerT6t6ERx5QhRT5K1+GeDwhn5M2eobqQ8w2sgaauAFEDqRS
YbJHgEEC7JSfSfTbJmXtGJfRh7Hya2SoDhU7YNT9P8jb15KJyXwDtlpayrmyXKzk
sTrbSXvfsLxxIZdDdDlYtFYiylzPLn5UJQKDg/avJW9XNeoqpG1taPenmGenRfT5
JoSTaAFY8vi9UeU6zcztqrCIyK6l53gmIxIK+H1/+Nhsi36SABrzzBbrzXxh4mvN
K1ueREgso/327K5Nd5e5io8abwU39JD/idzniM7j8F/d1bcc3piCaRXM3SE0yo0Y
IUekuGJy+q6oCftzvSCbtaZUq9k+N5qtNXMAUulbkJ3UCpvGgDnDAxTsZW+SGe9F
CNiEvunjs0xreu4C2E7kfmZ71gFlnCJ/hTaXoAodboa3AcGSQcjGhd6mhM87jvip
9WT588Y0vQJvwpanAC/qs8F8jCnhKwbgWkeKxcyBv/UcPsi+6I31MdQlNKijmhTV
QUQGeFue7sC5h2GVsZ6NbLnN7uzR7haXNeiq/JdBPfYCWAoO1HGNELJLB7+k9SoC
ZpbXn2PvBf3ZQnEImtnkf1bbKnSKfwESMrdZqgZU85v/hipyqDoF0soiyxVgxGl6
PfS08qhQ4ZaSs8eWdYgbhkxFM3bNiercGwpPiAn3GULbbiC1lWQ/pDPs/wcXZ3Aw
EzNMfv/CaHtMvBiu3sblp1y9RQh2a0fx1bbbKhdQ+nxZMR7asSQgdw9FC9cfLqUj
tquFwOyfeSZdj2ItNOpqg+K+c8FDFKihPpSwXN9Ns//9JkkwRPQeBSaRkvU4zfa9
5VMCjCTbmV/q5ImBsivwUtBPiJ6ySFZADeOXCDm4n1V96pf3ww81JC6f6xdPQxMd
n+4l+4dhGUwtX5M8mkHw3SRaDiPX9lUEEw4vuqzoE6uujc/NZ1VOPLv6uklOTW3w
G01KcEqQ0Qk/p5k1fgzwQcyeInq6SqtPeTyvYAUJrOXuZw5W15lMeAMGAj4rAA6S
CCISgGNAsf9wOqt/kD36cWzogpdF/6tChUhhNiD6rCKtzwQcfvYCs1TCYgxrOLkt
gsGi+gfw6oUCUtkwrw63tija5qctzNfS4PKwdp9pazyfwjr3Y8z9Ue2KXb5lNqJ7
nk+Q+rc6llNE/Qj4jQV2GqfUiusj+NCG7is4OFUZf5NC+2NQnXxaRRFIimA9AR5n
X2byitUJjj7IbYILorzDJA6nM90wm5xYMwvtDlzDGLe62eEfQact5Zk0tFTvJLwq
rC/G80/+dXUPNdpUs3Dor5EK8HeMsUyvIPStyJd37LgZdh5KCwAgcAUbRojpBgp5
FZL0fOJM7hPcFSahYzaQSnIkD8AJqKuIOotSfe0ZljbmrgCl+PPBSBTsqPQTgDVs
3JA7KN/HDSwZKlR6Ntwfnqiaq4doab+FcSZ1KsH8oTe8Ox3xZ78hRvfRWp6lLa11
p1zZYBb9GzzG2fRp3cArABFtbnVuoX+yVs7YrBgGmHL8YHl7JCqr5wIwqg6928Ns
1e9ELTbufUfBAvJ/e8CFhCcmtZfk0iqOT+XdFFILy9921VGSScidjeiDUL/Em1zn
8vPv/qWzWiQpRscFnjIK2+iiuuTC3UY8TD0XdG2+Nb2ZWeeA6kmH38n12FoAlb24
opsS0V7OF2qAL/fEgMwykLzcpXelfBXK/kXn82Y2N7cLMn8xbmHZeV2LNW+2OT38
uUetN7Q+MAiAQrbPrCj995BSqwJcA8LXPvsX96QPsMeLjcQ8L5e2Hd63lXT+f/tK
dkgv97aH1kbh6CzBvr3r0EoGjnNWjaLLdsKKK+I/ODQR7vCokO/1SeZt1v6yRSIG
dBbiclzcmIfnhsYlk1k6U6enYym2cdK3XOCBx2jRzqbdZ9s4Q2F6HOm8nFz0PqNN
Ox2HyUU8U9P7+i5YIvHYRxh4M1CFF2475InI2MFH1CYSJI2hDZR4UuMXboNSvCoZ
/E0WsAYaVbfa2vgwoWpiPLQyIKCSlDrH9I4p0uLTo9C1zjz5xNgA+Z76KoCfgkKZ
yxaJ7pmSuOLD5CWhGki8GI0xYevNME2qF0UKVvC+Ub1PXlCqKdD+7jtwu9ujlise
rEUTu2a3YrUP/M8hQnWYtg==
`pragma protect end_protected
